<svg width="493" height="421" viewBox="0 0 493 421" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<path d="M301.826 318.342H191.176V413.409H301.826V318.342Z" fill="#D2D2D2"/>
<path d="M321.165 405.833H171.847C167.904 405.833 164.708 409.229 164.708 413.417V413.417C164.708 417.605 167.904 421 171.847 421H321.165C325.108 421 328.304 417.605 328.304 413.417V413.417C328.304 409.229 325.108 405.833 321.165 405.833Z" fill="#F4F4F4"/>
<path d="M473.154 2H19.8463C9.99006 2 2 10.4803 2 20.9412V329.059C2 339.52 9.99006 348 19.8463 348H473.154C483.01 348 491 339.52 491 329.059V20.9412C491 10.4803 483.01 2 473.154 2Z" fill="#F4F4F4" stroke="#F4F4F4" stroke-width="2.4048" stroke-linecap="round" stroke-linejoin="round"/>
<path d="M19.8449 2C9.95786 2 2 10.4493 2 20.9473V287H491V20.9473C491 10.4495 483.039 2 473.152 2H19.8505H19.8449Z" fill="#2B2B2B"/>
<rect x="21" y="21" width="457" height="248" fill="url(#pattern0)"/>
<path fill-rule="evenodd" clip-rule="evenodd" d="M478 21L21 270L22.6825 21H478Z" fill="white" fill-opacity="0.07767"/>
<defs>
<pattern id="pattern0" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0" transform="translate(0 -0.0517716) scale(0.000633714 0.00116777)"/>
</pattern>
<image id="image0" width="1578" height="945" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABioAAAOxCAYAAABrP/8FAAAgAElEQVR4Xuy9aZZlSXIe9iIih2oApBZCniOS0hH3IZFL0rRfobsyY9L5JjNzf34jsxqQUD8ygK6MeMO9fs3NbfhsevgP/+v//n779fOLAn9iCrzfBou+4/f32/v72+329nZ7f3u9vb293N5fn29vL99ur8/fbv/pn95vDw94oAf/e7vha0+fnm6vLy+319e326dPn26PT4+315fXGz6qj/O/+t1/P/RfP0Whh8f69nKtt/kMy01ut8fHx9vDw8Pt7fXt9vb+xt8fHx7H/bwu/PPO/6/n8kL198Pj7eXl+fb+9s7ne3p6ur29vtY61mfhVY7PhPvjfysx1o/WtR5AW+3P0+OTFvaOHfOe4b26lPaj7zpX1M+Iz7y9vfGaj3iGt7eiEV7L/XKd5Umy7sOTmSWKdgs9sK7sf11D6318f789YI9E/qYn941cpofym9hD0sALezeN8JFP5kF858unT7dPnx5vnz5/vr2+vt7wNWz748PTDfzy/o69e7i9mhb4DOiBH28r74n7eQu496QPbmoC1Z+PT7xPnhPXBZ/h85OGPGG54ELH3rm63/v77enpE/nu7f3VZ0w89+XLF649n22e0YnjGT79mJbY9/Ai1/j+fvv8+Qv/xXOAx79/f759/fr19vL8LOJlfx4eyIO8h5edM4XXrs81zt7D7eX1lecHZ5N05/XEI/y/ou177c9PCQiyyTjP43Q2d43nuD2IrjgHeO6Xl9vnz5/NA6+3KW/yTFOW7WvC+kE/7oCfKfTEPfI+nnuetXkd3hN89yZ5FbqSNo8P5EH8kM9yLiB//QyQc3iPdPUZ6us3bX7KMBki7O0NvPhIOZp7v79KduiZJ/96jU96j0eYsku8L9r0c+C75Cc/m478kGRmiEVXlawAD71wHfl5fIRc0zkZTCuaX8jlnR5T/h15b57hIRfB/5HV0A9Y88NDyzepksfbO8+uaOENLW7N/aasyOf0nUfyxzy/xRM/eVDqvofP4x44F7qm9Gf4tXg8Ap9yAISV3Gl9pAtr/72bRSfL0bt7R7/xzvcrezhz7VGc8t7WiZFd/uCJj0L8eQfKb14ncvak0/UsshFWHpctJemvvdKaSLBhB0QffP/+nfIWcgj8DBkMWVl0HLZUzswdkWzDtDz2ObNcad7qJ32DnUb54jMUu2ISY9P9x50os8R8HXIN/gHf59nDS4s+9B5FXixHeB7njT8gK6EPnyyPKPseIa9aJ+c+kRW0Jbi/8whGd869Fo8/Qv7ibLxBV36mjIG9q+u19aJ9lp02zw5sYpyT6FvwRWyxT9Dzr89cCGxp2hqwaaAnn56og2OrROznX6wDMq/p2fbWfo70zOK/nbbXOuHE99ZxJh70J2jPNT7cSpdCfuDn5UX31WesA0Aj/P4UhT9WBF3gM1OvDgMR/K3nvd1esQ8vL6Ql7CLRNOcN19cauDbbm5Ew0V1Tr4v2uhnOPp6N+xIal/1tGUetomcITy37TjvQvOaHgb7+9rdvt8+fP5UdlP3L8+4yGnxH+x0+1udPt2fICfg2ZRPoqfp7kOO2A4cNLj/nvXQ3aWc79dPjZ4nyeTD85+OnJzxg6x7o99ecoX5dXx26bZ5brBcW+Pv7DTyPvXt5lg3I64OOGyM+vz7XmcCzxS6irQm/7Psz9x3v0Uejb/PIMxHd9IZzZ/pRBL+9yW54spx9sb1AtpOtRZ6xbLxTRw/wb18oY7CXtF3sW1HGDRuQ/DiuWfu7PWfxoO3xq/MoO1n8jHtRbvM8a79xP/mnb3w+/Fs2mPdGMuhBrsx2I+wFeAtnNfL0+fn59uXrb7fX902emm+mXIc8pP1K2Wv/22dI/Kr9p+95e+De4jzL5p3eUjNOfT72Jvjl0T65+fULfT3ogdfb50+fb9+/f9MF7rCH5s/4HvyXdg/48un27ds3+aWWMVf2UvviY62xbRemsWK+2FTIwPBNnR/sq3lhHCE90uMjzwxsBjxf6Ip9J9++vpZ8gA9Mfnl94dmi34+9KTwFtHy4ffv2nf/iGs/P2n/dzGfCNNrPJ9db9ryNlLL1p69j3TceJlb7bpNd2XRY23fowtdX6mDaSM/PXDPOg57zlb/zvZcX3i37y9cfoVPle8qHls8Kfoo/g23iuTX9YYfpfchX74vl/tmfv/LzcW7tY3/+ZMxJ+oMyc8O4TH67eiRq6Xk8W/a2bYr4F2dGC3/H3w0+Rv10QfQ8X/kbpR9XG2nhUWM0U6blHO5nZu799GmyL9FhtLNAO/s+2dOye6DTjLmU/LUdBvkcuYTPS3a8SHZ7j0H7O190O3ha60bb8WeZvJvCmP5uzvfpHPHs3l7vZLKW0TJEa9VP7JN5y7x76etMu/c//G//x7Xtt0ueX3//osC/KQV0CMjYcMwdqHh/e7m9IVDx/O32+vL77T//UzsBOnDWZQO4gLGAH4Jz45kWd8eg5E8/MkDtC6B8CVRMUHwAehBUONC6xgxUDJ/tIlCRNUpgQ+A9UYkLiJIrKED9wQJmiIeDQ5jrNUi1UmEGKgg40LgLcNSO7gTyJWLXZ4mw9g5ZTzRIBIVLZ7roJGNer8FYl5qsfWsEucH3YQSOGEQ9UAG8QwHruX3Vt1cahgQVbGgU6GhHVZ+0W24DiHtusPb9Bqfj9faI/zPI+fQo4w3g+3TiA5LSWKZhLwaG0oIRQpAf/GEDPDxezuvQ5wLrbwx8YP0JThCAd6ACRnPFk4RgLPqpjZw+HQJFYEjB4QBdXm+v7zC8EAyJk/d0e34ZYDQ9jnGNKLXDAaNDYGcGxlwHJz6TDvgbgBkCFdgbASTehQk2Cl7mHa4CFWQhHxJyFZ4LtAYAA0A94NII4MTJBe+Uo/2TgoL3WAVN845P6sLVDzJgBHYgWAXnDIGLDvQUD+8OzwdrEp/JWKXj9PQJRCowHvSHoQ16Zy/ohNvJncYh6UtnVCBFjDn69HCQ7VxHFotn8Fy5XvauF3xpmCy0Gw+4gJaWKBOYPAHLeN6AOHV829BWUEo3vDL26+j7l9U0xm4LBKIRCkeTgXIFnpYfnjvx3/HZrzyjiz2u9Q5mK6MczzOCwQlKTLmW1yZgfSL95AOum8LEwSGD3Qla/MwR+ShAUXquAHaLWMrZ5t2dNwXIzwDgYSXzUM5g+/JRU+AEVhC/GkjlurnnRx9rauDx2o7g+boLoIU3cc5Wu0EsOYLFY/kEeEaQQ48vYFW/KQgk2gmcfv7+nc41QII4xDNYGbAz4O/JCeHeMHD5qc7V4iQN5s/rCFQE2J8G3X4mw58HV20RLLGT8JSQpzxzdgaZ3DGTNaaIGWeQ9zo4gPn4noah5IN2RikzCSBKdwnUlO3UMsVCqdYQWTT13fTf9V0GKr58puyFbg6YFUVnNU9A9vOnTwJEAKx8+cLvJKFhihzoHOgJfPfp0yfaljMwkaB+gkk58+AzgCilE6yLZd+E0/zI4G8G3UbwkB9xgO0gGcW2K9/P8x/nH0Amnf7bjeA7wCTayNgT2lQP1q9PBssMTBp02A9wy8J1jx6QQ2W7TeCSQIfYhwFB8zdtCQDqtP8B3CqgIz3qmM1w+kvtJ9hkYCgAeRu+XvF2ngJ0lJy1biZghr0FeG5AJYlOORsAnXD+YgPsNME1YM+Cf3I4JC+elYBlYBH8mTP4DhS6fLRObgCvKRDb4A7B0tdOIih9A/AE9idB0GGj0MZE8KnBUaxZgfpOiJrPETriGZbkDQeF92fGGl4cUGCggTaUAhR4RgLyL7qW6MgwiOTZTXY4/n140BrBj7we/Son21Cl4vu6rgWnyFbGuzwh+ce324PB3viUSXJSMlMHY3kJJxRhLxYzajNEEoCYoOMmBofoasBf8sdJQ7YhIf/vkjXCsj4L8Vx3mieZCIBugq4IJn357cvtZfih/WyiN22EAaxzXQ64JpBBQB1nL7YpE2Dg/+mzV4GKkvvDRsb1n18gd7TPkLX4UZLOE/e5vrcwofY1CXIJYPphuZ4CpumjdELgQqvYv3NXd+OylGafw53ePDO02dvnKJsuymSzkRP84vnDc7+/MzBBn8l7hOBdgi/c0xfJCSW6SOe37ejv0RaBzurkn2AbDIQZ2zkSlo7rek5moDz6jjyyaaepz3NO7+lkR5J8Jf0mHutgKQMN9ueTTNpyUbqvfAXjDfE3s/+kma/PpFv7qeLh9mcTXFjWOYz4Sry6U27YCwc+YB9Z/4Jfj/a5cafIpXwmMrTWHXnVUuKOhElCJI2teyXnFOQ5/cSmTMCqMKKyG/KtWBy2s2xnZN13+ISFW3AU6nLwJoOtSYjuZB/iMw5UwLYI/+Iy8Z1j45VfGV+M+KGCE3iPgS3rICW/NiSl9Z590r8rUDFNmPjBlz6QkiN2cZVn1F4kCUCnhjYdP9Df+mOBiv/2f17iARc88evlXxT4t6FAaxFnEKqigtUUrKj4fnt7/v32n/5Jmej9M5w3RO4f4ZAAfFPWGR3xZMqusPflc56iyvhwsh9K8Fln0Bj3tYWB5wC3q9bgnjN2jnaDQIN7oFPXgfFHuCtguTNCJMABk/dPu7oju43G+5rTewpWzEBFCc0KHvABDXiP7HUD9NmZuUO5B7JkZaADiB+KPs5YGeJ63hifda0RqKgnrWDC7vRvgnMDJxKs+IIsqlF1IDk8si4loWtPSBsYEjNQYaHPIJSDUdgL8CH27MuX37R39czyP2CsgXewFoDyMcpvcGp8HuIQsRrnJiV6sx4REPV+e8f6YNzaUMSSO9Ny5lr698FkKxjUQAoM7WTFC6IDY9qQZ8qbjEY4WK2jvFMXAb3sWYI1NNrs8HG9zr6KAxgnI0DAYkTRyXNQK3srglRoazd88HaCOFPxToMjGUE5r8mI2YXFLoHugeMBdUyAagvoyPBsNU2j1QbT3Jv57JcGHQ0c8ZNo3MYOaFsVOTYS4UhMwykG8gTU5u+6/DybHaigUW6Ago5bKh9MuIUlJj02wvI5Y0xtwFWyUmLVxenMXm5YNLP1lkCF178/X55rrXTLuRmCOuw99A+dLlee0MCl8SmHldfNMzhQsWcS73xVnLBG4PePLX+f+DygB8AdZqsuTsE5o3nK1Jzpha8DAhhMCZ9dAVt3Z+YHcmF9qFkNYFrGMbfjFBk+AxV3uiL85z0T0NOO6rpGfVv/3cBRhZUXpdLq6MLMnoGFnTkPOxogKeK5Kypy/dPJ5ynXuiubS1Uv87wGhGKSXnT5DNIZ2JN+BtjnLPBkw6bqKPL1oG7F77I3cB2AkXHAwH/QKcuZ8BeSALL7ajPYdydvD/QToGGgonhV+jsAQUAB/FuOdig4AxVzS5ffQ+vJK3pMgq6u0sPyAvgHPBOYKb3P/XAAZe4fvicHXpw4ZRUzgAmwARxSECRJBTqDomDxpfkioJKccNl/Agc6aMaqCQNrkBnLI48MZAAn+Cm94UCIZIHty5Fl3+sRvaqiQgyrs1aZsqdztCVAjD3CswAcBH0BkjGpAdWYDsCDVgyiIGsawKETARiYMy/KrmpwvED1A38BpOB6EVjwPqeaIAE/Vq0EwIrcdWUfqz4cqEglp3dZ58L7Oe2jgDNYVwDA0zkiXzswN/0dfEfyX/6QQDIH1l+cLPOKyvX4Sw1UrLahbMpkCau6B1XEyhpWko1+og/4HLDTZqXiOIv4HKtIUZ2bDOu3R31nkfW6bu5JmiXpwsAf7+uq9aLpSVw6kYxVzv4u6IZAiAC79Us613qvKgUMTOY8Pj0oyIfnJOB7U7UGvvvyDGAKgRMlzTFQAXCbWfy4r74nn0rJdTxfzj6PL7oAP6y0FkCcahTsrYKQBsdnUot/nwl11DFb1clyFoem222SBEemfKbMYrxOiRuyB5WQdPfj9a9+fH8q2fmoSiBfuHqDvEYQvCsCJ3AWO6f0iJMR8XeCE9xHA4Q8M0PpCARf5U35rq4wZqDPfIOz9P35u+WefcbxsFOaTa4KYI/9Y4XXSDgs/8R70zS+svp1w1PSwMozzGg7ZszX92fwJJWACVQ4iTQyof2jrozAvoUnKxhuesjN6SRTnR1VHidwweAW9ga6zQJgBp4oA1PlXa4mftEf6lLg4IEDeit6ulaIzGvL7RgybIDzrXLemcQBeYUfnL3YE6kwSWcEVJrQrgFNoitcLYNnT2B9Jg8lSBza0n6yXSeZJtma5Lok3YVHdyznKlCB70EX7rJFZ/iez/BKXlaQ2nKeesTJwMOWVJWV5Nj92U8FsM9ZsJcZDDl+bVSHJpl12NQjnitRygS6TojgWdxs1kpydFKmTa6qEFQRcGNyhf3k/LM7g4LOE0OowJP9zQRk8pn4+EmUS3LD9H3PxJMu2q2k4IF5RP079nF0Romts+v2eb9KSMrZjS5JgI57lQ4qSuYs+tZ595m8W23fqVzc//jf/q8LD+qKDL9e/0WB//8pMMEcGfzQSDDg1PrpDa1nXr6NQMU8khEkOjA4iHGmWBrL6CVFrQQXkwglsXRYW3o94PVHgKcRstN1lvPfaxWdKMgC0lNnxvnCI3T1gEqB06YkNI4w0X2iOBdA1iIHjuST29ZE8PFzzrbYAxUFbQT4s/CaWXIyzLsyoFcVK8Bq3sADDc+0m2IJ4vjG3i5lYyPcC0Idhjzoq3YWrXy4fmZAD+B2Gtvc8kEvISK8iwoR/N5wZBdZfRGogFtBpf3wwPJtOrfPyD5Lu4x2pnmvtMahsdxOdgyx79++0zD57ctnBRQISDzdvnz+wgzHZNLwMZPN9/jAbFbykp2WCH6Veaq9gMqgHZwQ86FDmq5rZyktCZjRzjL1kQfs/S7eiIEbp3CQnhmWbCsRhfN2e7EhqOCCaCFwWpu9KsfUdA+F6ZZCWIYyrtwCjCXGATH0vQkmrKB384Ac2gbmjcyvbXsGH0I+qEQ3FPB9DHBQVlRmvFpxXboHG78F+FHQMt/qMxJ/jV8brbvwN8uBn5Q5gwwt/CiwNYKK+1k4iOkJKhcwKYZRVZTPHO5VxvBw2OmAOcNmBTu2NkGjwkLBDznYyTKqKhha1l6oEggjUC4rGKahvARqnEmp9iW6psr10/4utG7+eKu2bN0SqIBTM205cwaRQtZ5b8rlWZlhXtdrAn76bIrHJMtnsMPnkPsYnbPJf8OdFdsYTspHWjmNX/As4B+AFvgfZNHz68vtKwP4cojrzuB10G9UL+gQN8dHfkTbErSp0m/sOXSWAJw9oHVa76rXrD+nvPaXQqLeg6aTACPBR2ug4lTJNDXaMJztFN0bx/qMtUrvefT8CFQESJa6OpnZnfmLK8ZpXem0Sxdl4y4yrdrohW9WykqkBwDwMxqED3gsWSB9llaCDCY4GMP1W39LzyQjuQPBCuKp7VCJt/NjW+/IkacDP9qzLYCKv4/qQ8rkKctnSfmQqJU1e5J/bulDGWZ5UWAEnq/aMomWnc3ZF4vMpajany9C/l7blWxNcEIyfIB1qK4EqE7QzM7+FrCdoJgwDgWNIg8I7jiYD90rvajge4MuI6ni8fH27fvvpAVbKBJYeWDbHgbgXTk5dQFtaMsABquGcwo9hfYm+FH2bNs/VYEz2kHq7daFOisCx2UnJ7Bkm+biHOnMlGTW7yXSzdNv77cvXwV4//7779TdX3/7SlorO1Lt77Ac2XuiLV+lGT0qe/tWpFGpLQv06BVcDOdawerX29uL2uCoxaeyrNn+JoENZBGHNw36J5uS+5d2fD4zkRUBMhIEmbp59Uegv922y9n9eNbf/vJb8Tr2HZWb4AGsF74S7hOAe1Ya7LItLVsAsrFFnMHMygi3/Uj7DkC8gUiBravVqexStIf5fvvtt79YNzHttHwAfU3fi18g/kS7JAXTYDfzrLktVgKkDCpYjhXDWI4LWJGcBRiO53p9RvupBKI3uUzXUVnOOMP0g9iq9BN1rIJeapMK/v72LB0M/lZAT5UgBPke0E5NgDsAa9Afn0XbGzxPsvJBm/gKczWhAwJwv/32mypiHZxTFjrorvMC3gOw9WgAeAYWGnDurRFQ1tnIssWI+o2WldIBe3cBVgAgIGf5FrB5AZrjG1t+dgXDptNsX4G+z0jgclCKNozbdnFlo4VpfH36ybbn2ZLnEwI4zpCmz/pwe4MctGyCDZRzJmC4W00u8iv2YlpZub3Xt2+/V9A5bf5UoeHs6flow3+Nnol8ZKCY7a7Q9ug7Af9UlhAbOAB+01rRGWmFNX2xJGd8FKgALxJUT4vYLcAUfpEtrJ9K6rI+wB4gSBy7EedEVVAKvMkG0XcT9GNg+QkVcN/pf2O/o/Moo+BfuJIgCWvdCnPql9hBSdJovzRbMJM3wpexnazKSrOnon3XO6wgY4txtSfG81VVOt77/p2BjAQiwINpj4Qqv2rtiyosdihQ20C2cHOFCeWSg7f4Pm21BLhfXng/ym3wGN536+qFXwPWr0dLstRB12k3TP/t7ivUjV0Jgi0Ef2Jd3799E99YnyY4eRWoSAVeZBttMN/Qkv+w4vY7uP4fBCoIi6Udoa9Gnp3uVr2u50onh/AIkzXYdtFt9GAvggYOsuI79NdJfyVCTFmXcx29gdvxOwlMJkg+WtHN75x8JZ3xjwMV/ZhDAlwFKo72luRI6ZwtSTeylPeBPHVHDx+c2jsFRLTiq58OVPz3X4GKSyr9euPPQQHz8ZJ5ylIoz6h4ffaMiu+31+ffb//jP0rhxbEuwCCAXDlH8vDY9uSrnCv0EiVQDgM6GTwjuRSBCgCNowBjCcjvGbdy1BrrF0EbMINyTuk97ikhjT6MaavjDENE2in4b+z5iEeBkUaguPqBu996nq96MDYAwcwxg2Qzs3wKERrPWNfnzxSuv3/7XUa+y1cDarK0zVZFGbXShHpMghtRXipdE4ivvvsBR3Tv8R3/HSd3AbdXnMyBgGbTHdaZoForu/Gp+etFuwfa5oNneqnuoWsABUZTgB6qLoO/hSNUqaBnXyxOugwqGBRw9OXAPGsmhTM/o9DKEExWfDJDyac2fstwT49k8+GdXvC8AYOm1d+SgFN6Fk9FYma2epnK5tDIwWwwHVCzRmtL84GAgLRkU1n8sjkFBc7dzjkPI/Q3kr0ZwGf9lsjg9mHJqqKB3U8x719GwVGnduYHwYyq3lB1CY1I9/zHuYphvgtX9cXWHuregj+S292GwQT09bFlhwyMNGAcgK8dLmb2poVAwHqWDwuEzLqzxuVcjfJ5ZoC4TD4G1smAioNbcmbBJFai1lsDEB8o1AKUTxqy7YLPFB3LDWBPVksyJSHnYwidnLyfU36izC738106toMfBPjuEu3iTpMvXcE1AUnoAxr9dtojR7kit/MYx6wAQYJascknjSOzYmAmMO6/T6vMvBJ9dVCRoI0cNTgkyhCUvkjgMiD5dPT2eyw6YrypM3Ft4J7Wun9eOqsz6fV79+4myFFtIqKfBihpvZsKA1a/MTgyT830fAzqDLnPYK6TC1TtIPAseHeCR5WRBbBzZAVOx2V/5gaa7rSij+H59QR3qa8jgz3jQrig+obrp5/pZ2ge6a9grJH+zA4xSA0Ud9pvwsHU0kDgjeyZZcZSAdNamICX7CWAYb/ekcFluR85TFd8dnWKIQfhnDbgIJBhMRQXwXUVyOr2OOqjbuoFhU8gTpEog+3i4bQWSVXFlSzjPJL6GefJ7TXwFgAi2noA91xxoPaOb7evAEKfnytwlvYm4T3t0f3d1fYvLWzW99dJCWN1ORTFd1IFkh9iKFxXc1NgV6tNEcAfJgHFTg5I64BLeAlASgCueztyo5JlXbeT9GlwQEPy99CGzZdpSpvz1C2vWoTsgPDxbDFBW/ZdglFpLZgEEdoTtj2wHgDVAq36nFQlHXwMAH+vSszB72lL1kHXgHtn2YuzAt4AeAO/JuAqKwnQ7jCBGScTBLgp0Nr7l+qDn5cpcgwUZBKYi58A79T1nl2RuXc6I/CH5HNx/llmEOwRSPMY92XYW6mArnVW7o2DbLXfG702AIitXO0yKOM6vKPWYd8BVGZOCj/oqpxxFiz4fB4A3mIP0a5P8zEItI2e9QLfApKiPdtFWxfr9hlHSkvA2ItNhw7uSoa3lAQFXt/wHLIDssdd5Zdz3P8y2OqATGisigJVQZ1+GqbLWuArq4XpkZ+WrWnDNMEJtcYfM2sgN7w/xAiGrTXSTrQd1nOyjewLDJ859mBLMDGB2sP28+WcxI/IKlmFaKB/sZGnnDmBja4a4hr92dytKlzujrhaUTGw63k/oUuq1PBessJnVr/0k+dvGmxPwLNkgAOosnleqEPTGuoCL62ZTHp/JqYIa8A9GAyJrexKRM6GIaA9KnrKURdBYiMT1A52ZIVzt2+xfVMVfWA0Bg8QJPPMilQ7BDBnEMZBB865QMXFmGs3L1mBpbEeBZMtO7x3sjvWjiHLdbYgbz337hdsPJJrLH7n9LeimMvRuCfI5Sy+6Z/wYIgzr4IUCuD/nC8wzdb6TnR5Va+e1nq+fgXYnZBAG+SVnDW9suWCi8VV9O8ZIDlT3AsmBiogop9U0HY719NqZwZNgvk6Ig1m1jo+IF3J9WFfSy6u8xXjc8ZWjo2eZ5i+YdsSzUVZ1rRL5nM9/MdfgYqDSPn10p+OAj5MEdA8uBeBiv/0jw1Ozgi9yp9aoQlkFZjeA7ukjPnjzMBpElpW3AGDZ3rtTuDWHsiOt7I7OjO9qyE84I7DpdTTPcZT9AAzeOBQ4LnenOmS1gZWHBwIN0pZk6mwRFvGUjWoSlnbnA+QvqsWnMksE5jcP60E4lELXJhZt1VtYOAjxiyvUuHTKCY7H50at0Rxdee1N+e9g9mv5LcVAB/rj0K8U9Lr0D1myI0s1mTCyuCy4Vg3890SNIq6Gfci1DN8WjhOn0ZWeB6TWV5wtioO7YxsG1FR/Nnf6tVZPUzjnHoRBim07oAlba0tODG9s7Nj4F1YgcNCVRZ1sxwTPYc0oGio6o+AHLlfrWPpAe9MmYAUXNrqHGLABJMAACAASURBVDJoRKB48uj9MySwEIP5Hmgf3zkq9bVElSuxgxaDNr2WuyfvfiEPKqss0g5VyHEZj3FhRC7ErayOrvhgNlsBr1ljA/p0QjgXRLImPwvFNueJfXzdwikOykK/a5aZB89HWfcsx+lnnnM+9GwPN9u6+DMBewNGzRYsd/L7Yt17lqC+dw1IaajaClrlse5mVGyLiO7S2RzBBWebdaBi11Bt7umSQ56Gvkul2hggaBm8nIm01LgjUoCy5pV2oOHMgpcwiDWZ3Q5UFFg8WtDcd5oa/He/GQwpbn1Si18v+GYFnKd7nsGk7lcd3XQKVCR449J1gHHIFK3WJl5qL4HSfVRUrABE2hsEcFBrEgc7PTwxtoEAHQVDAjglnjkdhONrh727eklVfXoXFZoS06kW7fNZDTv+jnMqR2rIQAcr1FIx/NxVTnjuzHqRfJWskhPXl4p9pN6XDkZXe4+Pndmfc3UH1S7Qk9hPBJUMEjCz9OMW4PfbwXPfrSpSrdtOuVYcsLodXGc0czaCwOHSqftdLoKm6b+sYb9xihV4Z7/xyopWK47Ii9geExQ8sce/LFAxbLrOmygbRlUqaq+X7M1k9soe0HBiJOCALsj8x95US5xTSCkmbehXwSLZSwn4rPjMx/ZSb0VJzQGOrW0Zj2f1XfIzFYuPHHbrAcCurKXuMbiY1otsK8QB6N3qMTomn0mQeeWbNdv5tKaZVFFP5cxQAs72KVI5kLM790ftcjA/5NwaJG107+7vtjQESwnepvUohknLppG8dbDcM+Bm5S54QDPR9nZEkuP9E53Z1ailf4a+nWkvc713AQ4HgHWWmZdbiUKaR/Bye0egYnF3wpSjUtRt+/C5tzfPRnh9u/32m6pbkqSBZ0lAT1naAZKvbZkk/s0EkKdPSqjTPIEMnB5Dy5fDj/Zrz7enz6poYBsqtv5b9eOyr+73ruzllncFph/kGeyCZJTjGfHMCLyFx06CdhXlsrYbAPVsFc9fo+7lrBSVq09bXwky7SqVThn227SP+RxbMEdg4v0cElyr5/FJJzdWcJY1H+q0MRtm8S8u9FrbdiPg4M+mVVZhC5nTMfyNSfesO/ujc9mV0LPCSrORDu3BrINYITMq+zLAPdUWrFxwoF26sJNRkkSkve45EnOtV4GKSTPSptqFns8QfAcEHxI4zr1pQ7pjQyrQeOYvAmu8FXWOklRTtQe9jOod6Wy9L5ziYn6JLsSfnK1pFR91zvbi5C96khPDKTv/6koz4WVow8F/C6Y0Db1FmKZS5mdWrM+oSgdySK3xQveZ2Lre4nySZsJUJe26gwB17w+MyqlfiVeM6gxhnQnU9M6Ujri4NtvPjoBE8IM7UbnR8CPq9Tp9003c5DkTxMTbqRrrWYfLqeIfuUw9XVUQrw/38B//+//9h+3zn2eHX5/8RYF/DQpEmiZTzj2kCdy+3N5fPUz75RsrKjSjQrAl/x0CIwolAp5Zd8hofH8h3JSy6I7Os9OTfmJ00WZdjdY8JZXD8b02snwxZ4MZALAxr+/LSGVrDii2B2SEfOHv6V0sY3pkUiFD7dbGnMpzU8Vgpz7DMz2kuAIVAVdMLw1MFOjL0i1H6meWV3rk002LARkiFEg9AxVSmjLkTIuIqfr8lm0cMH+Ugy77wD/+9QMV2uq5vy0i8zp5xcPQOBLPfX3Ze95l4LI3O1BRgLMtnAqYsM2Rq15sLD09CuBLH3DqLBt9NOI86G1xqN7R1kXVRDQAq23Sw+2FpZBrNcQSeIhChPHr+3wcqFg1FXv9x7kbXyxDaVFLYhQW1zt7QpUcDeoJjEkv55y/A4LArQmgdQhUjMh/ywOtPXybrJUdzFHsYwMaD9qSzX38zNNQm0GBBPXaydsvNMBkt6AomaLFNhEG6c9BhH6+ZHvj2TMXYjp8ATU1xFPARcriF+dlyj+fjzgXdb0ELeZQ+pm5eaEKlrM2naQN4Sqj5sKRyrmtYWcOoMwAVMrWc8/ZT/XAoncrvq+cuAajyOPjTOwZgB9lageIbpzY7X4KpFW1Ap2yBBBLXjq/OHQqY3eDWhJM81NW1svWXieZgD9jKNZn3EKMfO/sdzx/g2M6Wxpiu+mDCz6ZL//LAxV9tQC94YkCfGs4t06CQEjrsDeAIU4uYDs4ZMo9ui1bn5zItAAre5Y1z5DnRsCxBujDrDgDFQGaVd1B6M1t73rOTmTKrJCKavwJUt59RDU6Uq0IVESGF32c2xZQ8rJS4CKnjKH2Y5AppacjUFGrQwa+2hTiR9nxTtxIEH3xevS5Cuj4d5oLV4Gsq6P8A+BmJyD53S0uwEv4XbJJWf0//+Oht5a9SaxJoEJ8yjf1rPW37lBtT7ZWS/P+4c/9NVZluDUOM+ENRpJ/bdMEbFrsEoNpCN7BdlE/ciW9LOd37sMmWPDnWdasrTpOwcACXDbaqIWF2rvw97HXCeRIhw89vBBletXmrbqIAhW9F1nntW44PR+DcaOdaNthF9ex7ROQLa2q0krKXEDME61KBdTCptf5AYCXQE1akyRTHq9n0HuCGGLD1U69433Le5w7ZjNbB4OHcD8NflX2vloPqo2L2nuoegCv4+9U197xzgX6wzW7eiRJGao4lx+T+VhJlmIrooeH21/+4R94RrE+VkJxwO+aMbpWjvV+SGdqGPvp5zJQIYPeMkrfjG5h2zcHD6riAzMYd/M3ti+v0yvQZdGySgEO+I1IZlurByUvkpiC964SJzK3LHu/BsLthDpIhDtn3/YkNM7l+PR0+9u3v5E31H7yyw1dCtLOdA3qO8mNSXxqS4kftMlhMOcqi9rD60EG8L2Ck5qJJMG4C5ic53UHU4Xx8uxkE1epUwfjHvZn2W75GZn7qiag/DI7tCVw70OS/rN160giqWzzzR6OT19VumKcI++JC65+NutzW8fpW2nrRj3jJMVKiqM91O2O0rUhLd/Y0sZtclX11bJOVXcOqjuYhvOKijjwLvf7IlAxeVH8JtwnsgZPidmOoAT2/+mzB0975kc95xZQmb5gkmPFO65eHIGAXKOB5bOOryqJYX+AZjgDsvnUvikBvN0f3TRoVfnkdVUa6ayoMkx2nHTeRzrkfrc/vnd/fvLXbD7Gu1Xy4xUPngMVC8g+v/qvGKjIwcA60+qUQfqL5KdrenTiaNkPCPom2eknnKbpj6c1fRJuOkWx29fryH9wsvkMft/8uu6TiVq427UMCR5ZPJ527Bs/RSUzqAd703aW5gEbj63vNC+2yT7wjVQATRzpV6DiUpL/euNPQwEzsTPknDplY+U+UPGf/6mj7xVbMFhDJRsniYdYYLpaEakHYEpg0z+YgYoBAhHvrUM0AcZdgNwrhzgzq6+soEKcBEZWObgOJcnqPwhlpioHORBqSZHyRj3v04N61k+Fmoy+OB1QYjH03ixAZLv1WtOnn0rOgzIrsmtfjnMOYHx4bgDpGn6ph+t9oBMRJ8e/1zolef2ns9M33osR0rcYqMQVcBvDInK5/j1/YQYO9NUAACMDw3ZujHZWqrCvYA9QuwtU4LldnkhWGjK5FPqDjPgCz90XlcBqW0JyLpy5MHuJBwCDAYjLp4omChPJP6ZwO0g1h8W1CO4hKQPaym5ouFU3brzNM5RBc2ZB7aif6WAouaR2BVzkRcgm2XrKN46wWUofByomb59AqglQTrbrzzYQdAfKma4VqBi8VrNeDAjnekXbutmUIQ622MDg0RjnY5FDu3wePb1D93oGV2UFVMqZZ29fO0wxcBmoUGlL3yHyL9vIgYM2ip35UcMr/Zn9PF0ZVw2A+nZThs2zuweDtud/dwuqZGLWs7qqSwk+Q5eMqgKz6tISYycv/v6jgYpcd5LyFNAruWZAvAFZETOl52kBo5kl6l/7XvOSmjt5injTwVuh5dRlw5ktkG/IuMmiP2Fz98fZxqQr0VKh04EKne09eHOi+em1f61ARYIUAl3hTCtYJ8xyq7DgmezB6GyF40G8oN3Lqwag3suQOevg7DBmCG2G5cYhZqAiw2CHXJ5zAua5SmByWcQf2TiK3Q6KqUmMq70qIOxKAQebrT2OW3eKCQjcG84Uv5lAjHj2ni/SKmh32JK80pUqcvYGIBXQKD2JL5z2SzL9wUCFZh68Vd/pytpki8if5XBJ/r1SRqC0+FPyLeBxJzLw0WmfiX8/vmkr1dIVppfmZGD4qdqg4l7pmb3wuFtdpU0HW8qkb7YDBORRi6OcubrGRpPrFed5W1rmNwUCwwMCpWL75N5x+rG+b9+/qVc67X31+o99GtaZz8gllsnZBlxA4QQq5rNdYQktlccd6OBjeGm3U13ajRzYBhnd0t+eZebvphpm2g2q+FLQGHJLs65eCGiBDqo+iA1eiqL8DFXV9EZdBvv4VQE1c3/DiwlYYC2Yn/C3v/7t9gkDkdnKR6Caqh8+aG1RmWMrUWiPeA5WAhPThgnd59wCgsucFfJ6+8tvfyFNmIH9aQMb76qJp004gp/bpp8bieooTACUf48KZ83K0fOxlRyCfVzS1B9uQ5V2ePM9tAb+gkzt755T0wEmgJYC/meWelHn5wSU5Q/pZ5pzdR6cq4qZYbAn2xy2mGmr4Fi3INXzxv7Xw4NPA3pVQHHcb1/sKwLDqKZiIp8SoQKSZ+7P3fnTQWl29a+pSNdMD+k8BD4Y/LZsxZakOkR2nXyRkmFlC3e2+fQ35Pv0nubMj9nybmmWZCjRZ/4oWeWqkc619G9beL0e13PQU7CNuK9zOP07hkc/0xbl9/wsaQEVOyZVI6xw22Rt+bxIxnBlD54vgaK93dVCAYPy2PMEO3GvnGsGVNwSjvdGwN399SkPXTU7K3TWIEUn4MmmGIEKt6Octopoeg5UiK76BOjDuTOYn2Na476ah9N0PgcPxUu80xaUkLzILMBceI9wDu6Z+zxFy2H/862dPjm1BKmD4/jDpfePUuUiUHElgT4KVPykYdXuq22UkdBB/XOVIvFhMNDB6sg7z8cgXT6g4+kxZ6CCUsn7HDqOQqtLOS05tJWon9b/U4GK0cp67mkNluxlgH6pTlSrVutIVy5eJzRFNo4K0YG/kY6/AhU/p5d/ferfkgItcMu4c0T7VFHxX/7dfZkgj4wvA9BYme7uSesMeJyrtCmicrPRNKGeympbBMEF3DIAoXZtRtDDxh6NRpf+XRnYHMQqycW1L5lCr2/MAsLgu0Sjs37Qq8qqOTjNMyOY0TBahsSzNw1wKw2pUqk8jTED5DT0kvk1wL8JwItbylxTrz0bsczeBrg259dGwd2Ve5+VbWXHw2mZkdedTQ/vLbs1lPPV6wXxF1irTyajvIat1WtQwPqM+CzGt/XHpgwD3LAaw7QN8L0EKkzSVCLAKMdPl81nbzWwEWXsdGLTP9NDvssud8n1zFJdjOjRPkPbGcTnztTn26XkFyxuc6wWG2kDYvT0Nnbacbq/nJ67/YvihqWMWopxyoLyGpo93auVOxQ6LXbdcLYOIhD0FZBokGQYJgETd6f+mE08h2dXFUICeOu6Cy+xPIgToH/jQGuxNTTRlV7J3g6fxbelo+PWTzF+16qxvYhMmRJzKK2yViNkdf89WPFDLbJgec4at2wqu+rS+OsvK4Oo2zPQ4bWsYpDVVWJ5flIuMnBWQmwL/qOBCgJXxa3aGzlFGei33iB7WyXArq4JXeMMJkCqGRgGx4tNWpItZ2d7ljikkesdSBuzW4bP+pHNHWBfe+4M2WUQsLUo9uXNXRVHoGLL76uVXq1fmuUPegHz87XXAAAw+FeAlYJ07n+dNhxWMaKXAhXkrgdlYFXVyOuLbfGudohxzv3bKqXIn+6rrH7pAqfEi0pWSCAxGYqqQOvnFjCqzPuSmHvW/kdEPBxItrXI4Oq8T+fLgJzbDQiQ/OGJPknNew9uzKmI5JCM1w3eXpERjkHTcmp0Dp3Dx490tWadFd95CRB/VFHxh/np/OzJbJznYJGN+9cu4he2GqzpEjASKJVKG8nxDsqIFxzUcTA5QM1xq5bONdZhuvHSFzk6K1m1kUOZPcDMV7YJ7cG8ZXpVUMVOb2RzmGdbmLfzjrgJCkz+iB4rsMvZ+snATnu8AIKRxwS13OIVr8G+1twNLWY/MuLDXqhsj9bEyYZf7KeLozHBybqPMxE74aGDMpcBD8oHZdJHVsSOofxwcAj7EPnSZ6Zb3ApUlH0fevLxLH+ivhZ528bX8pSwSSk77EekXVm1qMFQXVR3fHpi//lvv3/TPR8fNEAaMpQddVThefqZQNl8n0GOT+ihL9C2QLOR9MFZNULUtEYnGf3tb3/l/cseupMF0d1qQTd/Si6SaKtWmoFGqZzBWQGhdNhYl1E/aZ3joOPzq+asrDe2rcfZXBICvHzYlOdOLY/EcxkIi579qlpR9axbn1y02tqW7OBV04/AsKsdMJSbthWqyCKYQhNUNHlNdJ/LB++nal5PspKqPhRMc/LFaHl0J0qZRGjfFW3qPJsGwchLW2iRP/OPBAF7Xp/4RwICiX6Qd6wcq3Y7eq+kRdlkoy2OF70HKfByAhXKMZE8nuuegDrllpMl9sqMC9FTL8cmraedcu8iUEF9P+ZMhO8Z7Pz0idUPd/sxBgIvwOWoyuBzOzEKuACPp88/fGsED09VI7j/S1pvucpPYkkGW6owcMbxs7dSartNMzfWszVkfWgzZkJWC6klOcx684L4sQfwNoJLkH89JFszKcATafsUjOWOpraBcL3YFaSfbVrZjuDNMQfqYk2xF8pHbZV2yUIfBSoWP6Uqhmz7b1e8tB3HGtp34sae1zQT0H7A+MtZcuVy/F7OarqYCXJVacHbMbEnot1VwR/YxfV4G88Jf9AXe/aVXlOMRv4AKUH9dZZoCVTos9NG6bMRMpW+uCLtRXLCCcMQXBRjtqtfV/xj3VF+wxhV2al+1rmVvwIVP5Lov97/E1DAp+gnKyr+y793Rt1mTHMQdqLpNqKSHRHwF4I/GRJqyzBA0EGJao+wAOFr/+nFwqBWp1Qr+YIrs18sexQq4+kLKicwRNnBCw1DVIY7nS5nDeNKVGjPL7dv377d/uEf/oGBigAfXcauGwdUh2BIST9XM4XdkHtpP5Ehd3r0CQzolQzio9FZBvLUdhFYHajg/WelQAxQZwNMhjtmfUyas0VjL/xOdP+BQIV3p29fF1sduBiPMSrg9CgghECDBe8YwF3ri+PoO0yXBv2Fs090oLxn4AcpLisoG/0MVpWRpqGvcLRxL/KSMwoZePOQyZpqmeOUDh9DSWmtMOxWQKz11ewnu4qGMvbKON93Y/0bPM3vJFgQMDk62EAAT+C2F6FdsrBiCq1KkaahFzl4xL/GuNB3Avg1MZp1psJfn1mBCmdtBZT2hQMm7+DF0b5ImWz1Uw+TeD0j6JkVlFGug1zt2vCnHBdlw4JPO9uoq77Ex+YrZ4mpH7746TpQIRlGwMGZVPsQN4sL/+PduTCsKEcqrajpK1nd5dwffF1nBKW7HASqoZAZlk0IwMDNNN6z5hmkyF4xAHD4uZ9Rcc0b+TqN3HLMOxD3URsYOkIGsUsDhQc4fFlnnC1WGEQOm/vTHtJs1tjOwNpCJTIrgRo50JGrXdB9smUFWOry85xCL4V/8Bk6heE16jPLNINIOxA4Sb+e6eO2LC9eAVnFY1kv7602eapWlOMfh1agZjshyr6LowC5ogoMzZVQGyhVRtZmNN0dqOh39KFXAknqpU8H0wkEqtaQHUM9w0oNz9zhgelMJ+yLesMqozMzk4ooZ3/m0u9DxisdXw+nF47Wcw+QNVugQ5yoi205BZN4Yu4V9bhCdF2/9IpqFQfylejgQEUpphGooBPXsiNnVlVim80z7npaK9++cjqv6OprVmXaANiOvPwjR3vIYjqzHkyc3zsZQsGFBDKwjPSOP7fa0kwoPaD1x2YP8gwEfDYxMrAazMmBp581qFdnAS3pPnfbCdqrXe1BnePB4tXOY8eILuh6ClRI/LQtBJkPvaRqZOinzGXqhA5VTD/eHjgcXCAtwMbZlm1fwpRPDe7lU2n91PZ/AmqnY1GuwGZ/x5bmvrkFRdoYHq/zhmfq1nqlQg3QVhUbbUXJC5zrL18+337/XfM5kOCEp1hmihisme1ZdtBszrCaa2sZlPkssvFqzp0DBJmLUK1R3ZqHFeTO+J+g7LzHR4NT095SIrIDY/lOMuGjX/Evh647aAG9Bfl332pGex3Ae/IK75N5Rl7oLksSfJae1E/4KABVtRUkwOcKmwfop8+3F7Q4pkybAku2B33C0X5Ud1DwOrYpB4xbfuIKqN5GSxz8qwDd2+1xqwbMndL6KcAung33TEA0VT3ir3cN6Oa9erV5RgzTTkAoPMd1mRgqACvrntfQcHSBzQosKeBydbYQDOGwbgdPErQ7zxfb5Xs5sbov7duenQAZJ/mR9oPSk+nDnvZrfIyx2Uv/fi88lQXr+UnkWAHIqpS3XA8d8mwJyPJWPzKQJ+sMDuwnbrviirYF5tqngJ2CM/vVw9rLFrVejqzLWU4VA/gBshfvS/aajz0DifbY+42zVf76178e54vw2pkDlZbF1e5YVQn4jFq/iZ7cFw/QrkDFoSJlqiSeb9M3+jDVPbJ/V21xZX/iOVWtBX5X4IpVHm/vrC5LtQ5oCExnl7nL0R/BimkHZLA6kxQRqIB+WGakrTsrOejYW54jhDqesPYfpwyLTbcHKg5uZF31qpvX/pwdeL0wxH5kP40Lzp2qiu9qdX01rnu08N1oQhdi+Ai0Rn7Q8mpZwwgExE+kLnKyUemGKrHqqoOrQAUxD95k7UihoFQ/QLFtCav7DU8gi/xafl7LpfmN+Crx8yr46HlRE8vrZfQg9BlYIR/NIMmvioqL0/jr5T8RBYKsJmLnDJSLGRX/5Z9QLbAeIQgPGbECoJJhy/ZO+D9HpMvJd5n+4rctALlKy5WpJAGnuRHn9DgewjLGBNSjPD6KpVY7rIY1l+IsbZfPBNMcJfCdVTX7gytqf6VQE7XdGUCPppss4ZsAzZseoTFH8FDDRlPKCUUdw+Uvv/3mORxqVaBWGgPJSInjyBJltvQcujP2et12/ZXXyulORqadEygsBIfosPgLexR4OjozUBFeQkZNBp6LrgJ6O9MeApmtTZ3toeATgzt0zGRMxYFKx1l8HAYVjHvclwPxUtrsB9P9BDrXsDzvVSLxnCFh5bXsK4J3VIKmlekKUCd9ZAPeBcSOc8fWU86647pLkXUrpii63olWnp0/sJ7VUvzk45lFdqVR5YBPxygtcgLQwNkTuK5+2TOolGMdOmo1pukSxOj2EpM/lnM0BYYNIF7JgQReebRRyOvZp2LAhSTjlC/Xzzr94UXoheLDuphgstvGgSgx6OvsuFRaa23HcfY5XZJBVjt9Ya+fkWH5QgPyeqXAkMlX/nBnnshZTwA2skl07aVEDirusc5F2HVF7/8uAU9/5/6dDVc3DpF8z4UHJmAxiBlw5XSnk7xWIY4N7AQy4nissMYF4rpv3skZYOSUYFfK/iuzZxqT8341DmfMUnhH5cIzjXBW1wnB7AqqEdwtwW1gWb13NQtCuroz5sSnve4rh72SC4q4Hk5aDLA5nCeE+n30ud7pyx74AGY92wn74n613R+770F5/gbARY56PTOe53WWQ+s9PuOM2W5MUlI8utHZjHRFYxtkRtSFz8f7jNZPT9h4Ha/6wY7mT7VR+EAAHI/QSfLrGrHL7pIi7mroo/xW2dcyJP2/ZffgBzYIwbWLOREJjGYvkh02s+nms85uMJMCl6Q98Ggcsn12Sci2J2oErMf5OcqIy6jKWZYFhCTtcSbdCvAjMDhXuuNZt0+rtccOukuMl8xsMLgD5mAl2Zlq/ZP5AtIHCEJ3b/P07wcw2vaLZ4cxWH0G76TSZkdty1AHaH3MygbIuSRAy1kKsWtjjwigVdAgQ5CvMx6vtIr8gcwx0WnO4OcZTGZyBOfIaZDqT/84qWIB1wxe9Gw9yS7xhZMWDje4CiJwX0fSDM+e0SrZzbq+AkQKzqadWIBvgOCY1wPgLv/ivTVp6n5R+B6ylEGbBEeYpMD2KG5n53kV+VtJDG13w0fBvZJAluBOgEnJKJ29PA+TBthGRpXuoFsy7CV73/m3qh81KyEAlED5AEjSA5Lzmy7in3dTKriOV85QYKiiv4a9vmHO4afbP//zXxmQyLMFHBXg/0yQlAEBVLOMAE/JfVTkoOLQzwjawddF25qsshPqRE/o69jknEvy+Hj753/+f27/8I//eHt+/lYJAWxR65Y8mk0iuY1WQsnQj18t3arWaAWgbWzw9tBVfq1StUr6lqn6TcIX2/LOi7itDtupaR/gF6YdcvwrBiuQ2BC/3j5YZEWqy+vSY2aXWm4pSAgZiMHx2D88p1w0zLwQiJ+/xUZqTym95JZRlegBwD/VoFLXCTTy7Ix2rvS/2Zrr/gyVqrdc6GqExipqTWV5X0ugCr66yobn3djD3EPKJPsadbVpF4sxKyDIpIMkkvgL0UesUhjVDxVEXJwWfan8UwdxwWOQOVhL5j3gecGLaQWO77AaIkj7ts5UuWQ9qTa6sksRUFfrLLWgqyqZzBLd7Nvs/4nqBR8t/qYHhTuJEevAWUMwg+yWBKIB2FNm2lclnTzUnrrvoupgz+gIe2kWkGRTwHJiQ25rmhbCmYV1hUstyUxbcOJIW+yhZ6GopavOD2ReKumU4Kl5f8Fe4oOJT3WOOF/FiUTSKapEC84z9yKVBcEC+wzrCfD3bPFUfOKAGe/vThzSEyO50PLh5CdK3mkgb2FQCVqPiuh7f5fKos7D9Wnud/Y9yl5Tf3lGhZInc91uqlX2dYIR8VtTYc+/t6DKr0DFz2zLr8/821LA4vdnKyr+SYoqP/wNgYoxkCslc3wPg9YyEC2HixKq0aRdEFL52UjAv6lYiFKSQepMUlZHyPBItggMyKthcT+idT/azeSJjQAAIABJREFU+ozu1NOgqBUPyrHxSbYIgiBx/9ArxXlV/tZitldIl9MCcscS5PgLwINg+8zhr8hec5DENApdvE1roCJGyLCqAphSiCPLaN/r2njRZwrRjs5bx9jQhDKFsZAPz2tOYLkzg8WTVHgD+IiuiCKJU4h2Y45daEV2UGgksDWnHSo7yxVRd6YtjU0ObHWG/HiwUogwdNxDVDR1tD8GWRY3GSyBa34hA2OL6KraqEoaAYXsB+rKHjga+KoyReDAlalUii9KrUrmo7yOzVtGFnMF3IIZXEFAcVy07jiQ+qPLthlMYkZWD1acgbcAgVq4dT7PeFcSJehAZ2kzIJPFMNR5BS7FB2NPRka0xcLYldWDWP76qUBF+N7fnBeIKI0xhOCYjTkTb/5zCFRsRsS4dn5tDlifYxXIfS5XjrHZPPqdmjOXs1z75kASoa30oN+CFLlvqkwitjcx0UxfDDAPytXvlICVARsej0ysMtwCEa4IdpnPPdjpnv/Jg5MnfPlHtxK72IEjr5k97x8UrMszI/BwzeD2mu5Yrc8MjddxpvirDWNVYVBLOAN2Ls187GAaoRgnG0gO62fxP0d59HwQ0mkEU/XFnTrb3yfifRSoYAVM83X0nuS++GRBBzwbK69PvR6HbsqzAOe7Q5jP6DuZdaWnp3OVQMVstXVw2kOvPxKo0O7/UVD2vg1GAc2trdcqq6tAxRAqa8DEwRAGZOUkVy/vK3B3lu/7ueRL9bkrx+tO00V8dB/q/SBxTpWvy0B69PKHwZ4VUA+z/zCw8TOii/whEDcJNxp4Knl2Fawoq6oMK+s1V/HNg8kn/lGgQkp1hm6XhJhkbOORAELHjg14GiCc7S5oJwkoDVi1k0J6ewSrDZLJZhsbW8kKsWH7mjIPLPsJjGsuWIDtTuk5bcTZjiE5q02OmFEAnvkmAHYqJEeV2i7rTneVPHKyxdYWIsdY4rgMtMtkJtnEp7s00C7Z3mBgzlFVbJr/WFnrABD1DAIVaCWDTO2vXxVgNGinyvOLIJ0XxCDD45PAJ3CSgxSy1SUPM+ATT8Aqeg+vBqUxa0hgXFfToaUR9jeZ3qqA6zkwbM3kFkCsTHgXuCk/U4GLV1aC9dBg8qFB5/BkgTg7igzw6a4vuMDdVFTsMgFzF1mNgQoHA3GgH0BWPAfWlmCC7qtAeMC0oEzYN9iI5T9iL9wFQMtvAJnBtZoTon0iyOtKCDxDqryQtCBfUCA8W/sZIG7dnsCB/DyCxazQ0Vm8P9tNpd1PTuXUZFt8JrNZdK1uRaK9cwDANjKv8VnJEnjuiLYCe10xNAMVGvztqmvjBvLZWg8moS+zPZLEQRngh0x7p/jLzSv6QHwz7od1PwFVzmGx/WZ+B8h6h2kMYtJmG/qQA8nxc/C1r7yyer5Ue4O3Rr+fY7BJLLjIHfqXPkucK5Rn8bzGpcXb/G4ElNd84pkZqFh4abQPSwUj2lABJ2B3iwR+8qVDUGWR3x/YW0q6QXBUgQMEEaTrZCTvoHCD0PfyV3IkMzXFnbQJGSCWr0fI4VGJspAL4LkEB7HvbLU1tDGD55a5qUY5Sf6rQIUqh072jjibtgZnrCr59/on1lOc2MmwF9+Ke8KKeslfyP4EqKOvEwwtPyEBbso+JR9VwHsGvw9TLf6eQEX2uKrvxzmjJXtVUTFt07TUXOa/icaRNzN44AMtuf8HAxUnatNErwrcyGfplZ5J1/KsA/QDQ4yMGW2w+NKvQMUH5+LXW38SCrRgqmiyje7jjAoGKnrpI19LBjGrK2RECZwUWCy3IxmEnYGzEkEHL0OaYtUpiq9WELpwK5gIxRjt9N08MG4B2adw+kBgXxoYQyjL0LCRZ6UXYzEKEL2ojwLnIuPwDohV8LZ+9qvxEUxfGujbEDSsEUYsMksWo8YOzGKrG3RPRhahLV77jwUqAgDJ/+v2GcmIk5wsV5y8EQdYyjvZsnYQ0FvXrTDwvQTAGKQJQDXoxCDL4I0A2DQm2aZA92eJr7ON6US5JQ+u/4x+3bhn+hWWwdtZigUMTjVxx1NTiTUoqJiKNjZGBl559bDFBEao3J1lmDLaaVS1IdqIxgr0nMDZBCpw/wFG2nA6z0Ed7aiqrMMwgo+jjHW1dUubNZHDkENlgOe1AS5udhF5wA9CE+t8jCo7LnwWeZOzOXlt3Zr1gstfPxmoKHPAX97BJTna4jM6ftPm256nAmEFbjjbYZOxJfjunGxffMMzs0Y6YIdrzSASrzDXFXlAJ8izhob8W2mbp9O/+rxhgjuMtVzkn9R90hq+sMusDejb928em9feBsWHRPPgbis4qgSOfEgIuQm0nJMP2t1MOl0+MAMVyTpdA0wqn75nng5uNnngP9ExINAQkrlFFyzl+YDjmrP9Cb/PoamPt4cEDQb37k7dfKZzKGi2slsZX2MT9sOwPOxCsv64gqNaS8vVLjnrawBMWvXquL4LIZJVzmGrIdy2WZQpaWng7C/Ns7DzYBoVoLKc+PudD9jBClMdFcmzgePm94c/OjFwYsG5tRY6GWnn/gN7zsooz9vyJdr2kY6fM2qu+DzaJjyko7gKiDrBth/qWlfBj4UBmaYrjZMWf30QLpa18sOPhNJluPPCntTLTqiJTnOrust7lZz1J7jEVGbujIm/u9rSp96fj3d8x8x8gTZUZWLqMwE5Ub2A1jVm7yXDOqBDA7Hr9cW3fe4bmB9acNq1PgKcXWMbT1UcqHR1izYD0AI+BOr9ROh5WdhTzSVoudG2Q0BzKZUA5ZfGx+F8s51QgVixYTqyumT+GiC9kqeXr5Ou5u/hg1AfWOdWVngCqQ4wpUULwWC3P/kC0C72eADKc1dGBYmZNYxBtZ/obwDgnIBozeXzsUrGrfjMrf9en+9aUfK82i9KRYLu5wx3PItbn337JmD+629fVZ2B50ESUQIV8D3tezAI4ECKAqnuO39nQ7GB64YFti8heRJgss+lfD1VQDTPCBTtwIZkJALU8yd2anRZMuGZ2EL/xDJ7gOm2sMT/Hg7ModkZ9qy+KLyfZkF1wp/kYtrYjsBI/BvLcVVgqMJj/5ngl+Nk0isgFWc0qn0X1sDAkgMfq5jWU+B9tUBWYEK2i2yPOVS6/Dw88yFQwWtFhqTNnJMXQZe0Pkq3Bw4CN09IviloVvMrRFz5ID5jYOdUSmD1kEGoysBr4l37Q+ZxgdHrfns3y4et9TwhwQt+0/O9PXQA0ouWDmDl/MXXyN7VuWxxtwYosjwGk1SppBZOOrzskGGbZ/pYSSCNjCpfzcC/7DRdg2vITDW8XnP6hBplbhHkCeSK2pCpe0J+dlmIIFDxpnn2ugJNCRRlX6WllgN7+/f6Xvd7F2VYlYpboDs2ongKFVQ+B1XF1xwR12W2jIwMv7axN/lhAhFDGEFr8Zn0RPCSn5mxItf+Xkdf6dnpg0SWySaIAhEnpWKCwXDIyep40LpW8kCJmORFt+XVvbe98J/lN4vgi3+z82Z4qfSzMQbxp1rKZt/02VFxMG07On5aU+vhJAvom6up6s//4UDF5hfhuvERRmVOzpgiIfZTY1u4fZlXpbUNWs19/RWoKHHz65c/LwVy8s3qlY2ATIWX2/vry+3t9fn29vLt9vr8++1/+qcMtcwRWHPteKA8/FaGKjJjLD7LgdwFkAEH2FnUdKaWD2dKQ1NZMQMhMmy7jDpKUllsrfBiTEQcXymEfH8VFS0IY5jEEFCptcqOOZQ7Rs55Vt3WbmdwxYom8g1m7sap3BgI2xSjNr018RHNyJBjgF6MX3/7TQrDAleGxChjNl4QwRWa0Sh8/HsCFTbMTYf0sk/QqRxXK3T2ei0jpwFG7rFQ/QpcibbJtrNBRF3gAbUcJtuZNFErDBo5i5ytUQw8wdnKvArpepVos8/lGKxU4Ep05qY72d5s0/NhYinUBtToPI3S3/SefsGw9vpRqXJ4G9UyreCtSh2Q6ZZBzbFWpUdTOc5Gg2oBjJB1ca8g+zmGMVDKUGtOIAprhsHpFfospCw1DyfLWedI2GBsab9j0G6o0sOyYhzNYzEN6vX3CTmcntFX+SOBinGZ0DI9oVl94NZnpM8FACpDw/zrzOQZyLLUjKANWde/bZhOg25K5MUguYz6TM7bQCYbgX2d0St8Aeh6X/VcI6Aw+Hp9iE2o3f3ZykByQydasrf3VNs2lMbWP3Ry3kWq6vnlQ6BC8mf+rPpveSf89AHLzczKhZeLOVbrN8ZmDPUshq3vrO8IujdzOev63vnSdzJbykOmmaEqZ75/Lhy38Ykzj18HKggC7HRZXrh709mAqQ4RuCXwEkJk62dMcdVhpnlo0n4lDuwyRO/AktGfuB5bSBiwo4xxH+dkODNQ/kGgou7taUUzUMEtS4VddbP8Me33Jd99I6DXOIeLqLuK0n3weSW16NjN/uSXOSB+g0tZgmbWjevBaZk5FvrRMYpcSPCjHemPKlIurnhB8j8aqEDyASohWRnpNgh8zBgmJ/G3L7eyD/bZN2Yg8PjyGJKTs/VTywIiAq4iUKBivsc2EmgB5/YlcgVkW8cGwu+ZU3QGM3FFz1CgvZZ7pIRaSSZkHa8bdpiCE2rxqjZiaiEZ2zADzlO1sPWU+ZEiubHq1gCIABWA2AqOhCX7925DeXfh7vS2vJXqglIOoz1IevqXnTuCA0cWuDxEnRUL/s48mbQUI+WdeKP2Fy2LEqgAbTPHgJn83uvvaJGCiuKLQAX2XzMX2q8CIJtzJr+iATK1ctHFAEji97RHmpXaFUwwkDVbpQYQ0hw47RX4I1nS8b0CcifJhQG38F1a5L6pVYnO33ruaRPf8F6/rriC9Ncy4FsC7Pb569fbt2+/V8KMZsuIPhmmjduoDQxayiqgwD2qoGXPN6u2cPZ5VEEt0F4Z+gL+mcX/8sIZMV++frX+A8AHANfVWq6gYDKWWyylWiZZ3qL7qGKKfDYQdhWomKottsjk4QRe4icjgCR7v8V+bHNVbWUYuQyrDrLYnuGMiiGQbZNpF7SVAemRxU4aeT5O2hKp7Yx2N3Zk+wc5/048GG2rIhjw3cxhY6stJwFSLlp4lD+SWViHrK8S+2ybo8H22OcES/JMk55XOMUMSCQ5LHJ6tmOa3w8NqpmFnzVBo7wfORIeyXrYriny0i/mxAQMnycru5aW07xPql88c4XYBSoNEBh/6Bbfy7qHPEwbvVybttlFBZD2L3wi+zYVDh/ZEh/ZbxMED6akYMjAHWyH45kgE6qix9hMVQMPGk5c6azMVqOk6D6SmbS2ThzJNcWiPUfpqHN4wYPh84E9Kx9ErZrwO7CeVJExMAFbwdVSZSvfBQU6ABlbnngegtQUwtua/Gf8n5JBwbcqIaEDZnleBSaMFY02gKJb2yozgBT/PHoDiUNy2ZOIq6uXT3pni/09FRW7h2m1tc2xlcxxZVCS0YKraJEl9/Y9/xWoOJ+yX6/+aSmQk//HAxVxMeUaJSqqNhBTOKaGU30+O/snxw//5hoF1zqrLkEJ9u2kYQhjLcZFG1tdStqOB4314RTk+EfQ7FtyF6QoJ7Gd6wm0Qzgls6ydHIP7fzhQESq09vqoogKfghGaFlhRBDJamgbKxqf6cu8+WXdX2Z+ZI/L3Bipo5CSreoK1bnMUX6DpuJYf8/WpVD3/JI5H9Recw3BjyNBqGYNQPYj7AQP8bLFwXoWH5MGImIPraChn2DENqAwHk7Vzwi/0mkuilw80j+qLHkg6DGFF5VvJUeGnVzSqSTDXw1ljpxgC97+CcY1+SO2ezC2viQ+zrgffuA5UND/lzOCVT5/lmCk4oV6tEzCWMr8PVCwGVM3jjlM4BrfOm30gP0umjCyj+fEJau8w83LZnw1ULODZappTHlSALfReVjP+WIMC7cxtWfy79e+/V4hczLdXeyxMe/Ii6rW+Ws7KbFNXAFEBEjEip1Rtnuqsk/ns87M/oxClFWRgylkMv6sVVQZgnh5slacD77u48f3pzhNOIHCvQ8qdKbd8BGeQbEY1TiENJvKPqpuiUITDAp+07J5GtyTQ2Pua39BDOSMmplSQ/ChE3PIO4OqnKlcWsU6SbyXjVaCiPrUNHSBtV3t8e+HuTZPSfD6ycNXmsalLeeBesnWPcnBUcUn6oYptBL43Dbw8YBxUDbRM5pfbdo1AeRyoS+4GTmzgpUwEVMOkGhB7x0f/OFD74em5AzpX+d26NzSeQfKmQqnVRflQyfa2bsD6FcbKo7HxuQDG5q3i/VRU/HSQwlzKqLfb+hS3fMC7c4Khn6iz0+8p/BGAcd4P9czHT/qvC5jK3Kf7by2J12s0SSfRj0NdQaKeAxV1bA/9pnmJIV9yUVV4KuCnfzCg9PtiQ6dqklxyMEq0vM6Ez7mcwNM6VlOBUoLake8GXBLkyDN38HsrNx5kvAL2HtyiI88WYCGyDfdY2p7SPjrv6onHr2wu0CjtVApQ+4EyunoG0LWDHeq5Dn2o4IToF1uIOih2oPcV76UNK/uJs3pYYCuuy/7tz7ssyNkSEJ9ElOljJJjFiuSaVSO9XZXBr7o+1492rCPTOTZZg4CyGVkNEd1jEBufCWCKs/WCdmVVeaENS2VQknvUFrd7qt9vLNrcjue2vS6FmDlB0ZMGJElLzQbEOrOlHH789avntaFfvQbPKyVWtNwDFTMoENCYw4FfRLO0QoWvAvqmqolZ6ej7zzkVGowNfgYIrnki3bIzSYPUX0ju27LLG3gbs/ju2L+DpX009BueG88amzEViNLzs5+6Loo1s6UtkiJGKxLy6JsCYEwiQ+uc9MJndb2qXCnCrFMgA0nDUamU4AQDdPif21mm2mXyGnnGFTlrQt9qnycgkOoXrhU0d5JikgTTbmeSr+jlVj2pdIYsUZWTK3bml7Zq7PlWaNJ4igOFVAn3Z5hnfBFc7dDmda5htAcruWAZgQBZzcCwDokOSEXKxFDuNO9QXtxzzz7Md3Bt7Dvalu26JfvFihvOUnJQqyqQznqeQYIXnBu1Y8N5Bd9F3oWmU+Z+lJDQfOPEmHTWmIEK81x8QcrHYQdQd2ZOglsP/ShZZrfB71TT7IpBYSTZEP7P+ZbeO/k647XhXyqx8Uzb8FkCFbOiQu3skPCkSh38q5aRK/4kEatg5AzW0EZyy9rlHMWONyDDpY4o6KL/ElQLnpQgycBiVDVVIIRvJdxCzz1kXra8aDIDsN3KsNdrh/BfWFFRPuZWqZq95OOnvW/889h4ZxNmhQV+tX66oNKvl/9EFKiTXz09FR3+uKIiDlUUyuuzjLYMbY4BjcMUpdyZKWtK1Z3QHcNu0r/7vm+hEBwaw0/IstFAx6wnAQTJMd2BgvAHsMuylulQpF/oyJSK48FntRFePen/jkDFCjatkOrJZ9IA5sw2eOOcigxUBc01YBtKX7MekmVVVvXMHomD7+fTsxlAMbeeaDOBumlMJAAgxTGyLgMMxWjPgMlUomwGkCxSgQ9QumzLZAes9jPK18A4K0o8tJAAmu+B73EoowdjJ9ONfOssWZadZo8zvIjZ4Yf2C1GEjrKX9VxMZkNXG0vTO2CNqjfiaIpGCYZoYJ4yvNITehoqc4ZDB8hapFw5zcVRXF8YNINRDVLcSaY4v2sibOyDOIUghbLt0uN4Aoo950Ik64oKVc8nYjMYjYkIKcG+FpfTuJnG2Gbvy0e0AbdcbRphXlvt45I+NsyFUY7vjdVXkhW4VxMMgyn31iMbSqh2DqFxmsl2+n6BeGve38DBzWRY84awLE6ln5FG5jjQd1UYqWQqh3Aac3YUx60a9+pnKpIXwedT/IwKlMEdYA9Gs2Q9BiJicHSy6nUtbeU2KGzu6Ye3PBnv4hlmgHaEVToEhnXYteSF9FGxzU7fgxDHx9M7FXKqKJTe1AfZSznigbjz/JcTNRvXi4QClydoaX0W4F3AloEP0HiciwVkvGhd+MaM1PljndtUqjdD6XuKf1CBwcV3ibaeexCU7L8SmE5W0rdHNpIGDWpOwAxiRp/ci0ABVqRDnCKDH7OfvIINh8z3ccHKfk5ww2BL7eMYpj1Bup85LU3gnbKiyxp4mGfx+vOR17p2fyevx5mbcm1f64HtyylN7+hl76w/D3GEy5AZ72G7tRIxSg/fU69AroS45iLPfvllpUxV09wzTssD2z0/CnaoF3HTepGYg7fC/sch9iWtsu9t40M0lIyKLrC+gm2Es5HgBBIl0N5Hw3wFbmYYaWyQ/ZF1p9GyJwGj0Y6nAxVaH0FCnJ3RH10DQm0vmXGl3z0H66JK8QiqMAjhOLIBWtpWzABNG9r2E3SNTb7cSa/1ycMy1eox10j82s8Qe4XPDfR8bnAL/zOfv7vFkYMT1Xed1bcN/EE3MB2HAKN6+AfEZaDCvdNTHYN/s6+3t9NpVWWNvgfwHLajAG3sWwZ3ByzHHiGoAYA+gS9yBT7LgNTMSIVdHaBYgRglV2nWGQM9T6ri4alwi6DII1yP80sI/gkQk7+ZuU8Yev2Fc05K1sgY1w+3Wm1u+8dv2ibP6w/wAQIew98sWgLATdWUAglpkYVnIJ2eXLm4+Y+4NudzwE/zgHcNFwboL1u6MtLpY8b2ajsDswVwZkFIBhIdQHlFlfYA8fDNBFXSBkqV4D61zni/mlEh2woVUdMu1WmullUbsEkSjkBFbof9Uca5Zwb4PFfrJ/bVtz3gqpCkB1eggjaqz21aXr1qlg4r0h2sY1a350gm0LfqQvlAGuQePggIqWTI6rMfPMPXyzwS0DNtiVYeXblK1R6oktHZCZ9WNezYjws1pHPA7gmqHOI5ZsJYD7rmeRj2EPdo2nR5zqiGyOe0G/ZMRtASuAL4iIGKqrZr/650abUgW3EWNjpg0Ex0JE87UDmB/xPIPKUs1/Ll8+3b778Tb+Fzc36jK+8OgDpkU+6ZQBNl7+jCMW1dzRy7oHwl2cbW6ETZyCbiXSNQxDaqbp8rGdiVZtVW13JOW3+16+vrd1J6BirIV5C/qlJMxRHv7xaju9pRcG36OS0fzymPXYktuS6dk5k94PEM8M5z4TrU6yPROHRTVxK3q4qMO6RbRkxXMp0uUHt2FaioNdCvUrJq1xvMIINkTgL4+36oK18HgJs//78PVMR/W3x19vwVzy7pjcNPqTUuWEdz0K/WT1PK/Pr9T0qBdmJ0+M30F4GK/+XfaXD1FJQRDhSK7CsLw+DhhpY71fMaQHnA7+GAxCebQNCVsJ73aaBCQgWG3pfPXyrDITDJslDvgEqEaUEVEHZWEgcD1g9ujFGZvs5ognwlEO5Mi8qSsKGF54oRvlJQspblzVBkLwr6nIDXFVC8w2ZoZyEj5fPTZxqsuB+zV9j/Mb2mx+6xamAYZ8avdZ9u8xJ9ECbms3huCPuk2giJ4zzXuSvV+V76Ue57vhgw2TcHK8qYzF7YdJuG2QLgDX6NkqTSNijUSluqGgo25ZxrMCQ9F9E/WdkC+AYGqieLvqzIgVfW8O4oCr7nDK0to3e1U87oyTRZVrq1cX2XreyFJbNKfVFV7h/gl6X/KZOuqhuhPVgXnKdkfHG2SGbO3Ek2fSdGSDud/cHFiJalK7nioBrP4xgCzGCX+RcOgZwQn3JmYgq0rh7WrqaSYbi2MJtnnQ4bAk1u15QsusrOkiTrFhFlyCar8wQuu2LFTpQyvoM/rdll8SXatDe4BHCcQ0kd5OoOYksrguIQI1wwFEErBHYpUxJMICCuYFTa1ejSqyxY/h77KgO+W2Kof7R2SYb97CsLsKAzVCPrIuubxztbB1dAZuTppzNypFeS1XVWqDJaAxhhxg3n91SLuY/cv/srpnd6AUw+FwWopC0KaAsgAW0u2FID2WFyInFvgRUO4i0BgxiYyQQvTjGQ1T2QG8w9gCp0QjwMc4BiMWCZNcRtMqfNz+yPPYosaouH7tx1l013Af92jLBnAEp4vA6gX7JdqdN1IB2v1DmecjAtnKrNXSUQOIg69Fc/imk0M2Upc2fvrlUzKcY0BmYPcDktSZZvJAGi8K6cXfkO1AloVxK5ZX1xrAQa53vZjvuOVgqeXWTGJdh9dTZar+oTWCNkBbnQGcyk/ZC3+34LrLvP2iy76qgPxAdJPEk1TwF/ESXRGxNMHHIqySGxjVgV6TY+52fejNV86KJCMvwegV2O7wQ2thtVRt4WKIue0fwY6bY42D6Ma2albW/yh0FXXANgXtrWFGiQ81J9k+eiwqV3cIZtd1nwoCUAVTxjbNXSfxRD5meuGrK5moaQQTAEuTIseL1X61rXndleC1nSIjIVmAkICBTIuROwmxZD1RZl2CNsBVTyS7xa9sQm3tsSOcv9Kzu123N0pmf2s9pZmURZK74TgIbDdwFkB0SOjPA2cTUFyDiIYlZNixSC9Jw3oNZJtFgPOlLDsNUeNEEz6EiC19zCe30h+90VDvFhTpnYpnPOHQH0B2TQz1mF4hPYHr/95S/Uf3gfa9A6kCzlfBSDszy/HqIKmsF/+/zpc1VgAMRmy18M7v786fbXv/3thpkafD5UDzw/M0CCWRUEUB+fOMcCr2fG4aJDnJjBFk2scnjm/L6X7y+qvgsIH4CXQQkHRnj23d7EQe4Mnsd1YEd//fqlzlRp8Dbuqk0h/LAkWGSGh7K7AeBh/aYraPOE53xRO1/QkoELZfFrULYTuDyTQT7w56qWSPvctdox59gzImiTqEJQ7aZuPQy9fN22s1m5Y3MP9k3AX6zxM3mwq7yxPvhG+EnAipUObwKcxRdqnfzl6xdXFjS/ZIA1B+4OkFj724kpAftJdw91p45EFrfbfcH2msGr3qPITfm7WBNp6ExwdQeQnKRfSF/3nRUre+WC9kNX1uB6BU2yWEld+1MHDAX3VLWA2u9J3qzVi1ktEkPgaz9mdoo+LNsf+uLlxXNbNIMxLfVgzwInwc+3798qyXOKiOgYzB2ZFXQ4N0lALKoNnbdXbGQuC55YfqPnRRgv6ax1+zhRuvI/oW3+AAAgAElEQVQ4h08og1QyS0IX55zVTA6O8CzZzuJQeybNqvoiOqrc71HBc7IZRh3XUXbu3wFeQ/1TeISDd5anaQmupKAZMHU4fNBQiSxKeiua2dWkD0K+Eu6Q62Y9Kw59r/vLHhkFiTSHbXviG7O6hr6MMak7Oslo18v1T7DDgSeVKZIS0O1Ko6tEJSw6YIN2fLvW/uHItotAz8qb6xpK9meuJOSTk37Vnk4YmuwV2SdTHql9d5/TVEfPNngnPpsYyHz/mMxi/qdt6G4Y+Q70RIJSXKcxnPie2aMr3OhXoOK0O79e+5NRoIXNzwYq9geYhxaGeRQ4jZDqAysFnYxrOdqdpXt1aK+I1UC0Wwe9vdHYgUHBFiEWHif3RLougjNGWMARe+m0N+bvLfinP5r2OxNYl3FicNSZCjJ0p+GxgnLKzJSABM3gEMjo7vYBNoGaJGddZCGqe80Ic9poBYRtBScqRdnOoNF6C/2lqHwyBwISuwfku5SL4F39JKhT99AH+p6HTZ70rO8xIj9cywVjbUSnXuYeO2kq9xjZPXdguWNXUE4AQASIKnOFhnwZWJ5HYh0tUPSe06Izs+LlEyOSYA6UPlk+NKnfb+x3mqBVncVhOE2G6SogBxRHubSqULqfK1BGnlrfMGdXQQpsIfpIHlVwueUCeO8zRWamrs5F8yCyQUQLG/rWtLi/AnqSG/hbylitI3KN8Kf4JiWcB9DGzrLude/MS2JtgQp+zshT+DsBk1HFE0OTgdvR9iw81wCKz8GVoKvX5/p3Xk8LG53hBcQcGXwEB3zOlxEE+zk6ncdRhhuDmZmzBa6tA/AY8hugyo7hNblF9wQ+T2SQHMswS/0+dc76nW5/ETB09uxdQZuPiU7H9t19zMszdmsUO8UB/HBIcB8416qqUwUbnPKWu47rLF6hZEfLLHKtaILWRAH6FwLe86qPiDIu0xt+ACWsT5pVaz/itwFS6tob/y3fH8EWA9zKMFSW1ClQoeBD/wS0nLKKEmZU3Imn5o3T/z6vHeTlKVBxPFNyjnWP8ji1FyWfpu6ZUtsX3GiUdmkBuQg2GlheHsO8dbJVGgRvoD97fenQXOytzgw3s3mMPNFX0jmklBhQyi47NX9m/zng9PURd2rj3xVwHr3kG4DfrnqQTdIBWoBmYAG4PresuWTzjwIVg0SyE7s1yOl6ValabDgWPSpxbD115TKA59kCIhEiy2jqYiYIGJQMgMP1eQMu9e/pTGhL2U6l9lk6MsDeimmLB4YV/KHUiN5JaxvqCXzDNgDBviQy2ShsHK/1v6qxpccS1JAdIf4lTFMsvIXWB1+GNNYw9WirJOu/Fulhmy5gtWSCMinbnpF8kk0leafKg88G+JQxnvkbO/HCw/vr4Ol+7k4uejN4Pj8v+iprFqB2KskRfHx+yzzBe32RNScJA7TGAHW075k/0y6L7Ui9CPCY840EbH/5osQqAMLfv32rYcrSORpYzBY3nkGS85rKezwHeBKAC76jdkaokFArI9AD/l1ahGCNTI7yehNkFbvZLvUZaftSfKPhvcoODzAsnhp+kKsndNT0DLE7NUNF4G/OZoFS5vfxjwMYoE3PMMStwBexDSQTlZGcgCbJFj3Mh7D90MzfCTQ4F28vpIcARgymduLRBXgH+74TBsRnAT+R5HbyyVlB7ap0+vcvGoCN+zEI9PTphooQBIGY+W7Avc+v6KyABfZPfAOef/7+wuBMPssAtAHotvein2dbJgOssW+sT7k+BwuSINig5BQUwgLwec1wQWDY1QlJMnBLM+xX5gcyQDls3KmPeUamLxU892ovhkhPQiECCQkMTpGfxJC3Ti8vXU35RLupW0khaMEfJ8jwzKFtmls5VUWvD36eI5dPsEcgaOvayPbIC7Jn2ReuZrXUlZwMLtCzC3Y9tiRiDh2H14MZxXfK3BD6WmwbpR8mZZr3E8TWGTYZPqh6rZahJQQvbO0hJN9rgHRsXW1HWjlHVuWshyclIzrAAdoycdP2ZoISePa0JpN8lyDI7Iui/4+XekAp9G0FEjVPiOfRVW1M2Dz91D5vgQr86ZZeiwwsvG27WDCx2usO5ZEP98hEnvFkLK+HZLnR1cfTHj6+ETuPuJtFcEy2JLMs0d4pASF2jqqNuqJ8BirOxNOrV5jnR4EKWWTTP9G1IPuhN6Y+2l3Ge3/L6/jV+umjbfr13p+DAmbfZHkaeLpq/YSKivysYKMMkFQC5DPdi1FGYoDFGbS4p8PB+7oroe7WNVRcLkvv0tZuN3N/fQl6lb/GIe/rFZjFYEPcHAMT29JkGPjA2zhghswnDS1Mhgnb+TAzJKtZAxUyxNwnFr1jkZ3iIWpz/XsG9BUPJdMgBstshdX7d0XnasbXWmgrTZlCMAqYJbZLRUbFIxwYCqHGqq+Ua2MpC3CEcuBa9QHECIEXp3PmjW+BitVulIpIeTt51covfXCz39MJBq3vI/ZD4QZTGES7x1X2vVjd6Qmw7kr3LlBRG7xzh64ZUHCC2uITtQ9o0hdnL+Awe26yDP1agmWNs+/zwsdjE+8DFQZISCSfv6pG6nYQkT96nqxa2W/9nM7ku0DRSIPNSV14ghkfBsYr6tU7MM8jDBw62B4Er0zIHlgo44T/XdbXpChL+kDY2TAjhoplktcP5woGVOROjPVyEi+P3UEObCsIiJvVqzLpFKiQG0GA1fNJjFb3FQcDzwDRR6uYASnR8aK3nqtf5Ay7dYTbiijj7EeA5tqbHFWBCcbMXafja65TlpkqSLAuAEYADOj4okUV+0zPvu0hRdDSCIj14HZgYYZ9CZcd+YP7TiemnX3RXudjBiom3e8uNniU54hnaw7e3XdKdK0gnFtyJfPI2nG5ja65SrIMAZ/yqRxu9iaXM1DLi+7e1ls3uhvG51KRuu36HAuPl7yYZ3I9d32S94PVvWt19nROlPW3UXvIpRP/FwA/dV173HdbR6oevbIO+gwBr+QJ85PIGN6ZWWL3+/1HAn7Zf9wLMgo2ImT09+fvVeUpPmuWqOzw9UgYSFPgQEGVADI/oYzuZNrhGI2j2UG2gJXnz88gyaK1DdDGFpPwDz9ZY7lSQElCXSGrIKmDi5vttTiyxxTD2UJtszNp38iGh67AagACl2xY7DHZgcFIP6CW7TuvbAK+I9yVQarMRne/eVUbroMpI1cDeiWYEfmixJCVJ0sTJhi/HcnTkVj26sgbs8pL56qGV/oZo5eS/UqezDDV5+9OprjSbOfXGxh0exO3imECx0HvRfy9opWOhzdD9yPjGoH2+x8BmW+vAowD4jLJ6zAEOL4V1rXoVCeLqFWYZFwGqiYgBcCb7RrdwigteTKrhXLxBdd1a6nI+AD0CPSzOlHZ8qi0KFDJg92Rnc92Oh7Y3cG13nVkh4s7XTFt8LZawIx5OQpOam8UgOgEEFWfqfp9TaDotmgLvUtWYzaSKlhir4pXNEh+JmJo75gKVkEeJSBEhrvNKtuo9KB7+Y9uZ2a7k77BOINzbS+2T1HJgqAN9jEVEhNE68A9y+/VcqfAb8zh+ExZjrOcrga//fYbAxaoqJgBoPgc+VcAts5/7IUEAkF30Jv+VQ1Mnk/TNk38tKo2NHhNm496xRWrfAS1S4nMkCGn1r7iLVXgxm6GX4vgVp6DwTPyKwJBg8c2eyZyP/Sbftp+JiPjwmsAQXF22oOeignBWswmWssw891kgSf4PKsiBMQ6yEhAGolUrpLxLaJfMiNEZsFIRFpst5ZhoKhobb/NlUpKnEmFEoIkmnWjHADRr/Ziym0+0Foth6AA6JhgEfiflSveY/lzSmAg6O4gcqrB9bF723NSl/q8uwldYiC11INPEb8wsjxtExVcmbZKPzl5L7PKMv/Un8WcjQSkoxdn1WVYvNZ0oXKOpuEIVCTICToW6H0yKKex5otmL3Mm7l3ug8+W77IacAvMOlCxmCTZv6sHuQgEXn1cgYpeF8gv/CfV7/pmBfMsP6L3s2dTDiT41PLkSv+fLaqrQEWfE32vE2D3BC4lo9Briz7fE3MGnX5VVJz34derfyoKlJTpTK8PZlQkUNHGix5mGZwzehVGUCcwwH6BHojWWRIrQa4ijVEyMSDyd/r4p18+XqdD7P6X9+SO2JpVFVOIxnmCNNBnmadQ8mYKHgAQMmokFORmMSMsypOgFsqzlPGk66xC+wkGm5UTjEAGfGycJZNnCidLqiMnxfGA8QjDJL0CT3RdXqv5EQ3OTHCrAFaXxartQldtsGemh4JFiK7OYP8VWlYJ/x4lHvZoA2CK/B+3YYk0r2bP6LxY2X0R9fp3GJuwjZwhlEFQMJbJY86Uzv2V8aggBVr7VoLL/J1lnG0ky4my8f5hlvK1cptKt4xnG4M6G+oqcK/wuj3Sywt698qBlLOm+1U5szNJGySQ0xxehENMgOPIgd2vUXsX4MQZEsugylS9TFCgM3+zLt23wTb27zWQIx5FNgGGfyJLrXscd6DgPjCYpe+BilipMaEr63AEKo4Bw1kx5cGgrO4Y2SILuaZRNa26o7F1gFX8HSXDKBsRciPOGqqz4CzKcOoVy7iyITaB0qUN3LqxAZZ5LKtKo0F8taVQNDnZjYuD68sFhDqyzVLm0Z8I/QJeMgjg1iX3gLv5mDQ06FqzA8Kt91y767OStdXTPfNS1pk7E8QTwPF++/b7N/bFxl6wotDC+mSAerWWQkMvFb223j8DWN60ZgWD47BGP2oB7dRH734crNjlj0HLkS01dkiD+0aQmkDr0nJtvV4HKroCZjrleYZaa1XwNZgbHdoVAJMipuUEcvmS1rXK/2iBtG6Y1xnrFvNrN/3ynZS2TJ/BljjpaWG1XGBc63gmStmYYln7dODHFwWmHq9UGb2ighN0qZv8pXo2Bcau6PRxkOJ8c8gb0AFAI/QIbBKCYnferB542jwTk2ZmZeRwdpHXuNREZ2LwSHykY1v6+/Rs0Hhf9hioiIyMThgyU8tvkEngyti4HZy52lA+wmkQ+hwQuQcqGvQDOKn2KD37ZVFJNdh9HX+dJ6eN63ZvFn0C+gbFV0s5rXQ8aJPBu5fq154Eg7Qs6OqF6BxdeDRSnCLIv2ff1m3fVctBuq3XUp5RJUDM50sVBd4P0LrOu+hKC80f6OSua2bsd2RnKSgQuc3seCYGrFcg5xsMfnt5ZQsiBRweHajoZI8p85hM4QHTAf4CQJ/0QuRwVSnarknyVc9lUDZ6ghsMRHgWW1bOhKbiec3BY6AH68acFIONpfcxi89+BXfEbToBJv3tr39jG57IDALK4ZFBrPTIx+foH7l6mEElg+Rp9yU9LpmiFktauYbBptIH1TIAr5Ok0BnqJz9Lvp1kXoJdsFk5y2OTg2zd84bAi+hIeW0fMjQk3ZOUYXmumQU6q+Tv2J5X4F2qlJwlH7tO/LRzavxgDQZG9Y1kLgYUZ0aA2pTFH2d1xqjwDV2mz5LfqRNYbaWzEv0pQFqt4KJHO05vn8G+y7x+dXVwZngFCTLQN5WTRSwB3gJ/XXnshCNUQYIPfv/2e1X6wK5WskpLkmnfzQDR5IdFrw0SR5ZgX9NWLMG+3ovhp0JjeP4WpYTtXZ5hDG83z4AOsEU1vwL+s9pki8fdtjptQUuCmufQqclJabTnmJCzArvLM9d8reiklj2cXfrixCG2nBMov7fPmlxXQYwELTkfRfKk5uy4coLyI5lzAfntnydl0FEPCvYr21fhwXO7rSvZjTVd/UDWZUh5/LCaD7h9bQlUuPsIWy+BrtYFCUyqsmy961zGB6bNean+slSeU5PsNx5pVbqxTa8jwO7r6abnQEVmu9XCWMHqAPspEWN0YLh7mA/24vTgr24vKAxAcpOJxtYLSv5yUgxliao855kmLyKAZiMj+/wRn10yTCWGbZ8Y7S3vSPIgvDE6bsrB4pEtUMFUj7hIvyoqPtqOX+/9OShgbv3Jior/+u9Hhs4QlDDCUmJYvdBtCKlHeLIuOwNkZktOWpwMvbwf4Hwexji7Afjx2d04vqe1LBQpMZXdSqbGabPUKqmQh+2HLrA9jp4NpgxDLjDDGdkJaJwCFdX6yf0xYcCqX+mqjWbZ1xWd6CQQpPxGw0RDtXsY3U6LAIw0bpTCICDjTug3SJNMxghoDbdSWX5d5yKTJ+9TKczPpwoyXuEATrJmBSoiYReuGSbj7EM+V5OM0XxvBTgKT3bQiJkgyZx2qTt74boU0wzDf9buzQ25QXlM0C3Z7jAkkkGsFeq/TfOPQJR+7rlH6X1LY+vYjqpBoNdXVD8p6zvGc8ZLcSUjUJGAzRwEJmfqyjRpC0w8GuDEZ+oHgYp51jNwbmZeZp86iOFyZFdV4ftqHSGjQw5YG0nLuXFbqkWucDaEgCMFKD2jwjJy2ZlFBioLuYx5v7eAcaeAhLxKc0Ayi3fj1xczPfsbAr00FwhZsiMQbGels8ki42Zbptlb9XTmvRtpDzPL62lAx6jvQIVI50y+BbXyH4fADU/iRaCCGYaYMeF+w6w2uyznGfI55e88gw3GnUDNzK7ZA1AJYlFLuLy8ANw5x8W3hXz4/u07iRZwRWCHh3zuAVkqnRVsnDuP9mol2C6DFJZx48wWwO/sOWWIdduEAGD3elGvTEdHNGneOWX5VaAioplO6CxvXuWZKm6mHJ4cvf5eIENZ1jkrWlefnPk0WcjuDSohQD+bjA17Rr/wYzl3Iso4qqcrFOGi63MfHXvIlW4bd4fRX23GkFGU93Za5ryl5ckv/ObwhBbu/eSZE/+tVJlO5a6Lrh3zq4BBqtLguAsg6UDWSgfrqHEmlqq1DF11tVZab/6In0+kvfJpZX4kEzmlvJNC69W6PdeQPbSjRFTxenTIbPVg7phVffO5DYQRrJiZ9GM77qurfFY/4PH0To8efPqkygomFVn3TTuzMmU3IoqftjZgo6Jgp7lwDw1fTpAjmcnKgNVsg+juJDe59qRbjkq6DoRk5cedW7OOk0YtVbSJjmDVCrw4AO+9TMJG7LrKyvc1ov/xXfW6/mOBivhKCbQH9MdRPQVcItff3Vqp2hm9v7jV3Hw4UYe+0qcvVSUSG2fq1Wlbtu4Iz6p3P3eCWf232++//+32l7/8RQFJg+/4nrL0kxiRLM/VRs8zAgBOSyDO56g2RrKtVF0h+wz35eDpR7RpRRsjvUa7bwT+COQ6Wz7DvzVvoIF9gNFlB6dF3vtNbYw+f9ZAbmepyrdUxjFbVaHtMOZd2D4pflsEjCo5xDMKgulcp5KgZzjyupg1RvvNs+Ec+I9PyFmGvl9VVUR2VFWcnvvKVnp2AAm0x2cyNDlJQc01DlLweTSfIXY1M7DrXDwxSQPVFH/9618VQBqzdiJBpcO0V+q4kMHsmjGCJCj6v5iz4Oxm0KwDqtalXk8nD7TfinvMOTf4Pn0iVHO50q3VoGQmngmzDZ6fXbnpORM3D48PaCx62+Mbe1zekFsFRs/G/qfdcaF0WFHkGR/EUaryP9Ise+BdeaRlKv1SWeY6U5phcON+4roylXumgQLronnmU804fz0HEzDdntABp7Q1rUyHBViNZ17jzqtNLitEUBVA3a9zoP0feNJq+HaQbiT3fXbrwGpV6FkknO8yAn7lt9tPyLmLUr7S/aJqKDCxsSvjrCzjMn0qwOJ5MmnnRMC7ZriVsWnbSzPCZuun6Bm1hxTPpY1ez0Roov1LAhWSj/aVXaUl3XeRSfNBoKKSSVoQhmnviThmVMTmkK8k/+BoI/8rBiqwI9RN1T5UVWOUs2zla7926HZV/0mfSaYo8JUqiwr45nxeMNsVfndsY3oRqLBUiKEZ5VwzxypR/BSosED+VVFxfbZ/vfOnocDfGagY3gDFaDLOXbqWvuAZiEZ3eGndgO9IQCwOxEd9tGPhBUitrEAZit+RTZ2B0c72OpG5hV+cOprbEUW5ql9q9/2URR1jXspXPcnV6kOXI5DvbJoEMKSZUlkxzUENxWMLF/67Rm5lnjVwcinoqky2s58L7Bm0y50XkC7BAQXWK6OsPhvAhQJ6zXRKFhfwpH1tUXpz/XNv4gzeBWaWCoplB45abHFSh5ZrTGxt7XKnS13mx0HhqTKwMsVzqe8kMnz07DFC76Abv6BAhYeowwB4feOQMwYqFuZ0ZcFdVei92z2/F/4r5Wingxr+7qs9g+Lp0b2IY8F5mLvskgyPTn92LKrnAtCgGT1Q78+YERpeK7MF5OTc47Q9R2TFrxW0wWMsZZY2mJdS5GXIc4KU3XJlJ0SCJ1p3smvoFnZv1xCZL2uoZcCr2rkpA2kwy8TF9bNmDlZOGenHwmji0QeHZlZF7BZcHACDj/M+oy3Z5JE+h4F5890rlNOyQGRydtuaudt8oxZEO7hxpfJm0Pn0mYAYXIGZpFsB7N/w84wsrGJxvnZ+vjtZGj9iBDiiW+hwmQZoEzB75TLwZ4M/QyAzzHsGgZctSgZXq+J6ewkSBHzh2javbr6UAIpsbruS+nzz/nVW2XL1UjfzHN8D19xrZCFH3rGPdScl7GeQYEixca43+063g0BnmzIniQUR/S07RLC5rnmAV03Tf63PMU9POf/LNbe2YEeG9lWMSYhfFRgkSDaB6HH7j0Dz0lHb/U6AbK/7IJXnQNKZ6TqfMXz9d1VUXMgOpxaw/YEdv8iHZWdaSS9JEtNeixMHgCW9gSl3Rvu+O4lwINSHdGIigvXVqKT9CNwQ97VtVns2wCn1nrd+zT3SVsbn2cVftJU1k8lz3rZrl1N/1wZuBUD2c8ckhtjhttVrFhUWTVXS4Pwuafb9ap13b882DfQbMxXZ/kbgVAHsnMNhgHmAAOoHnRVIB2uJWqFIZlfdrLdU3I7FBny6Y4ULMeGY76LDYkPvgIRkmWRXAnB5XiVjnc/FDARMusbuT396tjDxB052ZgUyApS7NQqCBfedouTzCMT17BMn5AhX6TvM9WnvUoG7+iX4HPyvgCIA71PVzfvQTlaLI7w+K3NDS86vIG+s5078j6xwtRdKy5fwD+fGed5KMl05M2HzK9X6SckDCD58RWDBlSeqBE8yXZSw9lOZtdJFmZ8RoCqZtm3vzVla646BRXDvtJXVHigRTaBt7F3pCfiyj5/WodHpqINn+/rlKz/DQeoApO0rznZDpKTB0aOq8oszSBUQuz+/2gnMsLev3/3Q3drHiQnYI2bt4xnLNm+fMIET+brKONfwddkY4YEE1hXkXttwyY7J2maCVyqMtM5Us+vaMoiYeLX4In0mEGT59k0VB5z7guog6G2A+u5yENtzt2/neUl2v3STgwnDL9/3I/vGa9j/yp4e9X8lDo1WQviqQWbM+2B1NWY2sNJa1T8IzqXnPl5nVVCiHSVjzLuer6YAtpIfCZBvZlbLjAQqIm17xkCCjgq+qu1ct5kbUse3zt6HpkkYYuvnyARmsrPsQ8Ean4WJdSSY97O+iHy8IWWXQNTVKWoUeNIyMqvavm66fpG3Bt9nUCPyQgmI8t0TgGk5OU7qXPbJOPxICODcVSKY2tup8uPiQkP3hlwzQCPNHFl6ZRdqQYWhgTcqSKIqhr0yREVEG+o+n+vKSLt4drhHtD3Yzs16zc8mE1CVPz2LxrOWomOcOXAXqCjsSIGM08+/JFAxeTSykZjVk+bspMPEZaBiYhe/Kip+cDJ+vf0noECESQSAM4mp0F9u768vt7fX59vby7fb6/Pvt//5H7+XouPiNzm2A2Apc0uUlVCDUquUp1klxBISKqMyWjtL9GbrkkSlx8AqZtS4BdOPiZqyORkokoZboOJRdEmWOeytVIBk/exTamUe5digfwvhgJfMji2ibaDZAlq4z+0etElG9+xrPIzN/bkjCGem0PEzLgmVkdhlbh2EScVJO4WdTeVMqQq8m25RcPTMR1skGwKBnAh4T6G5KcY8Az+yAY0B/o5KYL4Y3kkQRhdbK0aGgkuWT+5JR8RBMv2uIXQZsF3ZWKMCI9cnDaNtveUYglbumAcxlbM5AhUzLINer1f7m9fLIKaxO7But/SS3s1A5Z7j0EBx96rWax+Ak6Hh8bDNtXa/dpnrzkSa+8yPnw2iBtd9cuq5pgOVqgeaPVUG3XHNPmsw8GaFkRzlED1A5AQXqgdEZTktAMNutBew3Xx9395Ez5Ly59nqYKHCchYmNywHpjPy+Zjr+ZPNtZ1JkntkTI8I0RYKHNuyGfB8Ag1+YxaX5QYqbeCAsPz8ysi9ENBXzkQyiXbDbgd6GoQ/3CCO7ZjqezQUB1ArbupKDH5+T4rLwHnTeRrrZVB7u+bgxbnC+6zo8zyIkhrO0NapaV7I+ZYz2MFGgRV9Jvu5vXkbueQUDlU1dFZnEk4elEzhc/iSetbrCrEZqKgZMKMC6g5gjUzLePuS4a6akjXRASRXla3D+NzuoPhylTlbysROAFNhl1MrBCp57+CqGKiyaOlgn/oZL/2Q182gA7QFxHnWapbQw9rSabaaOxyDnJkCAtyCoXTIpE0ifEs7Kz/UxRneVq+M7ZEc0bomsvr+QiMf5fIufZ1ugXBuUHS+RJ+V+/cnOB5y4Jwt498/9r2bfVdVWLaAZMOd8exzpC8F4ChH96giB4NVFZvlcp3bZmVmK9q+roocrCM2wlhvyQln6RIkSbXJdL637N8rAL4OwiD53Otqo2MgCpwTIJtJBBUEhv2175vtGiRUHLZcEnD0pednmHqvdqLVbsgyzMBxB1Ou7a/SW876hm2IbGbwEcDOVFSIl3p1HWzv9rFpp1pHL9mj/PLDGbiJn+CWSNELBF7uZk4MfeFrJ0ko+I/cM4DqayXInKMQXSs54oqszUad4A352a1D06KCPf6dxJV2UQlwhKa4vmYEfFYLoAH2BjRlopzBJrHynDsG8OvhhrZYqbhQ0EWBsfCzZil0ddCnR80kiC6cw7T1HGjLdHP7p/hFbWdFRlcl1RIkls2ZwF3olL79BCHxHE/aK50nyQsBlhmk68dTybgAACAASURBVHkXCZKZh2fWfvzSChI7yID7K9DQgckZnN2Da9oPfZZVo2gpal7mnAACxqga+cTzBICMezWSC2YmDq6Tyo34VwkWpe3ZOt9OFkb2LEdcf/d7el2fSytYrB12KT739vIs0N3tYcufc/srVY2nuZwC1u/oFLC1tFv0qHkblRD4bvh8BuHC1/Ete189yNitxXh2DUpLfMs4mNKHmEpkscVYgPw5W0V2IOwjyCE8i+c7PCk4wQQQVyntdgGxlOht80gHfjYB68XhDCUwq2Qdnx8D3gv+4co9yvRKWlFrSMycAY9zsPnnT+Q3tUzDTKoEohQ4kcvj82dciLN0vF/Zyztt8QGgHT0R36n/VQAf1061CgicwPt+D80lbZ86Qdokr8ZW1vcaD+N3/Czhp7R+yp7GRrl6DHWu88aMYJkFStlk0Qa0TX1fVtm4PfuisXafveju+/hvtoF/VyviPHPL1nYsIntDt05Dss34qKRD0Fu6wsGTIbOy/vJziSGqWo584f2J7irtN5/F8EC3IW9csqvWtLp0PiFdOJNQ+6ZqqWnY+PdR/ZGqv9hzJ3+XZ//U7ioQxREHmtXyruANzjrOh3SIzM4FF/gVqDhYjL9e+pNRIELmjwcqpvosECZgcM7pfrD8PpQthTCccGapq+wsfRkL5LKwaYUmxV0ZO7jGHwTE8KSL00BtbqCDmRYR8DY8JZUsqNQOCNeAMPz69WsNF0tmT/clNxHKQRkuVDmp0zNcWWMqkUTfQQ4+78Ebm4GJGWQgrTx0qpTCoFnNXhjtQVIhEgdDN+y1Dh1Y1RM2F21feYEBrhZATQo/YMlHgYoYbovC9B9LUGzD3FbyxBGX4ZdHv4p0T4WVbHoatDYcE7CCYcrXadwqS5C/w+F5DQ+BbNM51DwLtQBxBhHLp9WKCZkmIvP6BHug4giyDvYJENNBsp6ZIuP3HnArkD+l4wb/CpxcNkprPOM1Fxq7sj8PNZ011H47A8sy9UfAjThPDVBfZYnLGE5fU2XueVBpVWjMKqAOXnCA5RxIaKfItmUttng52z4yKq7kEz6qs9zOSF3nzuaZhDjt3coyiwE337IsitOwg7OTr1YeOwUqsh+gryrmkgWKQAX7YB9+LoGsw2dP9LhSoM0HeeCNThX4bkAh1yIvxak22CF2b14ueqQ1mE78eTlD78nx+aCO2ffooINk4278JlChXsqE7ureOucZbu6e1kPXLifyB/pSsMh+sq0f+VwH/uM5yrBrVzORfO2YTEKl6oSSkH63h/aWs3t/j2rnUYFjyR8CfqZv9qjb2N0/R195vUc5+wNYz7Oa07e91rVLX4wqBeqIQ6PgoxNyxdC+ds5AAK38PZ2uAFJxnI7nbmSxa2uU7XUCM+e16ZwvyPBZ6kc2R0jHuZYPpyuGrwocvvC0P8ARjtQCKHIwiS4pG/14lk96dQYpuM/zTJxU3Af72G+lCuh0jnxeLH8EnnuPLs4sTVcOopyfReXGAARCmQJ5WvctMlNPffcUuBZAVOhNVgxgc6p68FAZfM0eC11nNIctapCt7QHB5BUDnRM4FPgOuXcvdyWu15tn3mwHmkT3Ah0A+hJwUEIC5Sg/8nh7fVd/8CKf9+AEfskOdAY2gVD11k+wtrevbRjRtLPI8RmBnJLA80f8ehGo8HPjylV1krkDPwhUFFhm8EfAGCp5dPcAwVc6u20x+W/Lno5e8QHlZwtPZt47k1722Dhzg9/ZRmq0I5E/oyHOADArw92tU0I9taVUEAM6U587J2hM60YtfmTTaxB4Z3Gn2gWBFdAaYGlaDHH/UdUPADVJdOlxXrRM6xutBba1Mts/q4LDrW1QTXGXwFABY3NGXIXZUz6cM8Bb7EoA8vjROUfcs8FqnaRwf4ixPtLEPdkJQt40u+7bt29Fp6mvrpJVOLPAradSXQea4tykcrUDJy2XGlCfOOxq7bYIUFAliTT45dOTK5/fXgv85tzMAeyl/Z3iQwhU+NwtNp32IO3AWOljUJrDq91WCbSYbdASaMOKBaQqKAi+wY+6MTjBY8wYoUiKPZfAxXjsDPs9603wfJIbZItqnonaJSEYoJkHrgQH5yVQMeSf5EHah94rOyaY8nxJvzw9IUiINnOyCxVw0Owd2a6eU2GQN+3YEKhgYCKtkGqOooLQNSjYvlMqDZT9ruCA7ue5FTkLP2FUyI46VxL8xQPif//9d8lG3yN4wE4R6e/+0Tyo16rQj7pdksNGi7Nk+lMnuL34PdXPynZqEErl+BMW6vJ3OqiP9xlcpG8hfZjq10oc3hVSItubv4AgJoIdqYRSJWkSoEW5yct3yXG5z4NaWMt6HPhF+HCkacWeY1DS/j2lRs0W3S146XUOkq+z1UpPMkwdUrjWvBXd7Jm0PMc5y4etmHb5ouvZVs460xfJ2TrNF4FN0nbQygV26e9ZI2qi+F4LLP2YpNVfgYpL2v16409DAZ+uKqn6uKLiv/4PMt7LiXIP1wXUGsEKnZF2mkoGDX8oRmjAQwmOdoDofLtHp7KPuzS9S2l/lqBaywMqJgKOVqDCipi2rNdMBxhloB7StmT0qDSdQt4DeFSu1w5Ir2oa8VzBJm3upVxaisj5aquEQaGDV549iOFOBVqgGwTj1krK14gSjKES4xLl0vj+lSJuAZ98gDb3l/xvC+IozJllQ8NtUiK8M17sgMS2x6PFyZqdkPXo85VJtwXRrjgmvUTjpDJjK0aie30mMEcFXGC3DL1kqpRW2AaAJlARvqbBimwkGLjpZzyDG8zmPCinO3d2/cwCXqXvbhHqAEggAybZL6naqfO78W8U9wkdmgbhBFhmNnF9bzqO82L3F14u5XWFhgmknR1qGR2cqzHKW5UF1hmpuSOz5zxgrnorB9irD4nWi9yLweIZGQVSXDHa/kDVx3zCTCUxm50OQPG81KTclBxesP7ZgJ76zun8lZG7yygFgLQHDjY7yyQG+fHRr8DJw4fj9P6sdC+H82S9jUBF7dtw9lpWWn5QdlpfLEG6UYWDdLtFfg3I455cl49R2Ym1kWOWwh2QADnel4r80FA6ZyONuSyRAyd+PS3o7ProhqHGmj3kigoY9nZC2PZpXvwQGOUwRfeSFg/dt4rq8wXYZp5VyaM+753dlMo7vXe/CU26VcbEmVrp9JFM0rXTjqgqo+ivb/IrINMpW+oj5nZQBjop2XXchwAGfD22ih63Wyps+mA4lsk74HXu5EnvdQXYcnZGoP9u2TN7YcQK5chlr+5twfPjn7nwQ1L9BBCxsORFmH2/B80X/0cc1TazhenPi6fyeCWFV9mhE1Z7wnv2jKvTTZApO4EEVp/l7FH46x4l5qDjR1Wr3o8yv9MWOvPO/l5BNPVClxMvDvrRjjXI+P+y957LlWXJuRhMme75Rc4NvYuke0XGff/3YZeBUeRnMnO5jYPqFqdDAZA9BZyzzTK50nzpxnknsIlI8j4Wlssh/+JXLmvgclVeEx8rnuFxZbkMyohBVK4z1lhfn9myjbupRJfrp4M3qSxFXDVnGuSdLegBoByaSs+JhTV3B1pQZhl43TUy5izHvDh+BkdMgjnW1VWm0nX0VyLjPZhzjYflkhipHMBpAIbsd9GzzdfTUXy2goAMfNmmsJ4A3VglwEJX7mWiuu7WxTKAZjlV43eXeyJwTied+0GRlnheYdcoIw3nFvbMSF8+HNH02U4u2nKMCrZzw0B09aFwfw7q7NZDLa8M+tG5x9JRdmh7zc2nA7x1Q+q4LtbkPhxYs6w4OSp4SKmDDV4HyadeckjBgHQMRuT2GAnsv/dnmdwv7ZQ89FW2ij3aCvTe1lsXDw255UbDZiA+jyeHST9PxhZ6DlUfd9i75lkuEUSd4+XOJYRyv1SyUqdKfE8RyD1BrfM5R523+vTxftBnA6RN7+zPxLUhfsJ9w9luz7D9yUbMCvZpDoJBBjkAAOfD8mOVLcRaizG61Fp8BLBWrN+2PoIMWoZWnvq9iOB66TAx2yiyfsIeJgAe5y7OlMv5IaBJvXKIn4wlch1AYVs69g0ZQHIGYYZaw1hrV+KwIy6+g9MPZUO7Al2/72zFGJNtv3hHDwqNbA/QP7Ll6ARDUOLMEvV3RuPHfme/vCm7ufFf41odv7Ez7xRUeZS6rVQxJLz4D1UKcgnKtXpCb2zuku1BD1tHhWXPPPtW9vvzly933/74o+nCXR9vfPiwgCz3akd+6BrBElt52Lbus1YJR9wDnX4hhxd9QffGGcNzxaMxKpC+cdAWwJa6nyjd2RRvlDk2nVlGUUePdWWPJJ9/n8HdcvyKo2Kk73pqJWfIUfrhqDic4I+P/0YrUEZXGupOg92Ufvq//k2GlA521rHrxg+lCOc4gOyj0l5AKutykjdU6aGuRFuPhHLXuFI33m9f1GA+V44KvUBci44ZNc9RaidBkmpuBMGsNWHUzarQj+aTDMieqtyYvoVIguat3JMNpznqtTsqrCDHTEJgosYmIkdG+9gGWDJTDRzKCwCXchiNOMRYr9uP9ZhmRwWU12wCSs3PkQvDUt3gqEhdKY1wPaE9qL+/xjTuyQwy+9s5Yg7GVlMoQriwHIeEaPa1UP1NeaoBwoWRgAjsUuVoHzaFVWcEkS4A0kfiYTPLiaAcJXJB9L/sqGgRBmUYNECj0dDO+z9ENc6Oigpx1Mi5hiOcUqxjNPT7GjRlwU6kBjZMO50OJNeKtzKYjoq8wdHsMkTvWSecrEwRHrLbO/0MhnWLbOzGyG6roLppL23ATEdUTLOngM/MpZc/0Vtmg7ztA3eyAezTmZsjfDz3md/EU3xWnDJv0ICG5sHcPWn2tzPw3I+FyxpUwRKt61Tp0HXnPN/uGO0xUfX5taOCJ70bR96T/QR3TgqveXENWxSx1876MyDF7xLwSyOk6HYUSDO1juPab09fy826OqNCzPktR0VkX9g46M4G86zkCI1uX1BaisgfwUXuTvKOQejaqTHvwxvzWLborevJEyyvy7U1Pchq1iEB50T6DoQY6EGlKcJgjp80bDML53zAcq2z1M8JeVBNZARFtIwvHatVv5Gq15QE8jOqa27oWToKI+gdPTvP/+xzOMwNNtf7GMvKzziK5OttEN1RsZxv0OCi8G2ykoon8frNOWryIJ1JLQJxXqcgJ0cFMuCH7+hnKt+CTSMYPRr2beXmJUw1PgD+kZ+k3NKgUtbtiGOSc30ejLil/pxAGQVj1qzmI1nXP/odjOOvpxmAX3ZDTtHcXz2fThbRt0r/gG6ROdKzLgkuxHN3wE2tKc+TI+NJS7Wona5dyio+I2jdez6t9GRHwsIrpEvHHVw/7fPuOIg+ODeu6SANwhHw+IgI+ajXH6B5rtH2fI3zK49L1Mr+iXdE5kNl5bZgGG5GD43fskGAlcp4NHDLuvnUnQLsdlYzMjYyWMK2JJ1pAPv6mbZY5sLJSUhnWICQcSmyptGse7T/nqMcciv7G3wsaICN4ovJZyaIgVU53bpzh2WYmIET9ILeGRH5/5ajQnTrRes2QudH6HmI/gqvAO1sp8LWfqejIu5BxPtPgtGg9YcAhJ8zYt6OCoKjc4iVeGyUB0WPEGbrEVh2NhGvGWVAJ+Zy7OFd3seJehyhb70auirom8GE4agJ24z1hKoHXTk9dXTlqMgR2PZqznsHqLkyBE5Fc0oAmGyBgtbVkraVzYBxodIEs77BP9p7sC6970jT8yMYoHjNqGiwP8XPLNsddBDZQg4sWRiqy+ycFJPd5wo04VmnTRI6W/yLc/DChujGU+Ldzqy0sw9ZSVmpgGCunRZxX/SHNA9PfVdyAutmQD6DW+Wc3NnLWyWjAOquCwDfiQyUcB7JwYqeHepvc1om7BWUuOK0XQfL+xQo7DlxjdxvQDLqPXuhfnF9Di6HlY4K818dNjvLeD4i+4O9DpKfTSXITjE3caYjU+7rb1/vvn/7Bt5GjcMyp2Xl2NG+CS5AhqX7R0BXVHUDZzkk45PjRRlJwLvkDI9LqDP07PNaSGd2D5ha4pCUpN0u5/mqwAn8ZUfFkr3IPcc5UOZy4mwKaK3gpmYvzzYCX1k4wUQHW1M39a2Rb2KrEazSMro+HBXvOVkf1/5rVsAWtMCV9CTue1T8n//GuoY2Khxx0tNUR6OtFO7RfuHnLpkDYD3SrSGcWZ+X/LObVfzcSnY6LVadPoXZuqZ2tOwdFUTT8Wb+g0NNRcZCxJ5a9ClAVDbf4ihKOi3mQdkwNTBABtbNBPvmbShzGGTCPYLf95wcFcW/i0kNoKo3QkN0CnLc5wjyXgO7bAmO3UbjVleR9JodFVg7pHzS+YF5MXxmNNffcFR0vxf3pwnxtuTjU/cAxslRwQaRpAG8QhkVqGuqsfPVDwx6CmEqmkGkUksxJ4hga58rxlruMsIdtfJK0BdKgQzI3Efoqh1MaIbvBdP4M46KjLTMSB7Tr17oKe3OXlcA89A34FA1sfmka0fFOL3+sqJFnksbBluqRMTaH9++3335zFq1MEYjPVVnbH5PB3qcmYS9BSI8ZlLkqBxRKbrkZu9pj5c046hlUwxjyfXzgpt/9Kus+JkRtXVqnp5xq9q6v3HmOI2RD/Pt/Ymk3zTONkpb8aUD0Q6Iic7KRap5d4TkWR6EzEycpsF6f3dK+Kznt7Q2OdPa5Cyzwv1dMypynhOwswMzfe3Ii/gyAwH4fXgWjbVaTyqe1bSvas7z3v6zWZPNdiDCdPkxqLQ+A5GK6oVhEHak1PEeRtmVEUBDn43qaBjUuuKcyPHlqLMCk3MFRZKNiED7k6I+LMb1WhAk6E7m9XpwBDvgsWZzw4nxnuhP9K4fLCLTxAHsK0K36KP4SGY3XbxgcFTIi7BnUeWoYBRqOzOSdfNrcM3gqHAkXzT0jKg2ln9wlDyiOhuoN9L0u1aJTooLXrt/2mEvGvhTZ7kiOP2aXVDGMIcjsGu9bys8y8nQ+eHuUhIBM2Uj4jTAVawDo7d5y1RyTnXmE+AzDfSJbtiF+TrkQGvqKSU59VQ7Enfr3R3y/XufeYLBBOspSwiaO9KTtfDVBPrQoHJZ8iYSc7fB1ydaVWkF76kbBWeUa/ae2m8EVbbKZHBPgwKtm86mXxPc7FHWFzR8dFSYybfnGExZ9kG6ZUUNu5eRSpuhIS/1IzTIzn6B+xO0+BncQyEBaOr7yL5RuQuOjfp/lJ2x3pDyqwRbbqf7HdgBFJkeMT70CWy6FJ3YLA1l0Bd8XHX/sz54e0fodGjY/ekTSzkhq3ksd9ez/dwQHgCYGpJ7L6lX0nGSIOzzMwBOl9SyXGeQB2U36qojgp5Nj4NHPr2MPUJcSrBIZKTFZL1dL7tnM2UHqTnKm/0gDo6KA+sF2P3MdXfmd6xLPJvlXipjGU6KOMMneaeoZWeqVJmnosdVHlCjcJR72jeDbKo16WV2GMn/evf1ty+gl59PP4ZAGjg/c2Gnde06VDufOI8te8QOBY8rZJuj7+Ozn7FGisb3kF0Cm2AAqx7ET/ZfEI8n2C29cM4SyEO4ZqRKKdIMCOT7fANLkc2Z+n1fS/GVrnvaZtmSCMoHhWPATeiZtQN9MMrsPAVfD2yEfN6OhdTv5PizM81RKGknqewOtKzEMEpX5vNa2cOQjc1KWaT9gdfeIyDNDhVl/cpBEvvlkrY+U5VlNa7KLClifKnftt4tPajLDlevGZx5HeO4US2K/jZzFoZLkyfdSmbhkcps7rRXQWiVHd1tLmAYE6+J+8OJGfdGWXSXc4TDl34GaiVYnOaEI9Q2/ODP6A8jWY9g5sBmBPqnQ3FyoCSmiLJvlfWfD5+UWa6/id2DsJIwYpEcdzlG4q8s0btRDYJOiWvSrulOjV52te/Vrio3TVHZohMNeCln0hj2qp0ZcP10ft7d3X84Km48VR+X/QtXQAdTHl1HGLM+29pM+//+ZzRKrSY5GSXQDukKyMzR9/zboGzVq5bHXd/Bg75xVFB5pjDMRl6bFVxrL+si1CC0o8Jc02Zdsw5tkCPaYgRVwKBeWG8RThuBFNA3EBXAmpPjD6N25Kedemu8DiWtZ55nwTwzn/78DnbNIN6sYMwgfYJKqplJ4VUChc/jVSvAXxKmfCCNCuR4ggBRg8H4Fo1F3ejaE7nBUeEoEDLoWqnBGbMRoJxTH+vB6CwkIu1wu0NK4Q+nglI6VcPUgDlLA/AOZghJmUqzy2U8iq5iaEjzVOYOx6r70lFRadpzTOSOgbzLUeEG3zZMG4jlaL8BmNbS3Z5RMUc497XvESPt8yErXefT702FpyIWmGK9C1lmhOPPnz/uPn/+MpR/AuiyLF59kudemVxQSnoywnRvRldvwK75NYPTS9GazqDCtZ22Ncq9qlIV4Md7RpB6mGc2eNc53ZR06Xx8jMPNw5pTSmeRU+jBB/fn6yzs2jmxWFIk5faertjqVWPvjfn9aR5yeScescgtaIc9ItDPa/JsclTw2DRQqjk7T47RdW4j/fn7ei4jkPnTUqFRZ92RMuI/Q6hc55VmhYv5Jtaz27u/zlFB8VLljLqjwlHBNmYGR4Waeg5OBPDrw17/oqOiHCE3OCpUirKCCbgvu59zoYDTqagAiZBdLGXBYA02rL+7+/L5C+pgM2uyWYObRy6OCm7E9MOxO9KVTqN+0bk8zezRIEgYWZ3KLlTkLLQJ1ZA/84Pbv/nLHRXSAQYWo1IT3c41kL2VvxeOCp/d3co7CplGrpzw22fd3UW/XQMlbILJcz2Abt3pODsqzEOSYtdzRB2cZTDm37u8wTsboDbP7eSoAPgoWWFnZdzrzFU66Rh9G//SebHnW8Nx75iDak4n3xcri3JA2aMiAQthKK23EADxK6e5Jgu61nVrtjcHNONjBhq4fO71MK4en7vpv664KuIs0g6w3ywJtwRMSe6jL0CTgcVj3c9AUdA4p/u1xlr2BHdnUClYxyVvDBKzZBB5lINFItsiy5uk3q110hKwD8RTOiRcXsiRv4zMZplbztelliKKnA5xLI/mkbPR++yoCN3eke/uTcG+A3a4EuBhI24HXbFUk8+z7SyDfM7EoKOiAmr8ufec/dNIi8yoeLh7uRsDEt7tqNC8DZDG3NKZCXJ5n6OC4CnXwCW73M8BwVxqegx7OMruAJzcy0H2Kolsm3JUGcjb2Rmx+dSte3kz1ZCfpZcBfYFxcBYESIw+dY93P37+gAMl1jwwBPdNKCDQyqT00Q6EbsBtlyUjBCAtsjkN473Bu1j/333ERsfDfaurD+eznME9e4KZMDzmmfWfwRF9EUbbit+EHco+FcCHBfYyWIDZQpld4wCSpoP76VeOCuAeKP3FMk4hkyOjgnJBZxD2/6dch3DexHjivIWDwv0D7ejic6qnhvXxWfWPv5n9ROPMvf9ynTbOphOWYsd4nEXopcouwN6iV2k4kh4JyIdT8RBskc5gB95q81K+K4ggGzTLSeySiuZFzEY58+Cd7gFHhded4kDlxQosp+gnQXm98VHPCHOflPTtt41savcQ8JX8sjWlR2+pBrYnvlDz2qnqeEXKM1ancMnYs6NCDrlWXo22dlJ5EmOU2It1Yp8cVkixthufO4sUJwjf12p3TO5KN7BNlg432bS9/4X3F/sw63qW8e90VGzpQs+HE9m26YejYrdUH5/9vVbAjOe2jIr/+c8x6pGeZ9YDhae5GweuvToUroE0H9IiwRzldWejJSrY9qQOAHQaHKpJDY8rGZCVxR4JPwX9wj9BQeFmQgZ6VgCeUaIwERpA799Z/gPMrIGMZYyJF2pu2W8iN7+EXirSMvK6mkGF2FEk9kAzfSvXjb/kzyCg9CmZbvWssBc/1jYVRCiBjLSpNe8PHiN1OYARwOiOihyWBKXXxhECwSq7gWol1CCGU5RtpMbzHOFF5UCRxCq5RUPNY9Tbd3rypGxiDWxEbCLICnPmXjsKlCCMajS7MZVq43Zjlb9XrUUAN1pjG4tUxio7p2eK+FnxfV9tgxgLhiHjcXBWLYUxuDBenswIkTBv3yz9DPqN1+pTd0D4ZRV1L8vTqEBjizIQBkY5bmRXGDjWim5KXpDlTSrqmL0UetmZnaOC/AicKA2OOs/lnOkRJSLy8VRes3pbHc6mMMjxFoDevk+TPpvJ7g3DiUW0dOpNv5uW6ZX0kXEkogwrmj6DSl1HKruzhIzAGPDBakwg57CRBjUnsOYwJe7RSIFWmGdDxjTS2O9A/1tgGVs6PX9xHq2DC/MMlN/KGdrA2RHEfIY8h6qtSy5R8E3JpMb18xztwFNLixNBjuvWRtQcbuZV2EWvi4xa/11R5gSLDGzOTiADYyx3wfRyGwzgxyl17bCbS4mZR0RJwR2/qPvGOW+IadBZpt0YPLGDZJa60QytwZlYbx0cfj4TU7QfT8b6UwaQ+PVQy5478vnTZ5w5RpuH3jQBXO2xO7D4yMNbveE6P+K1W0IK5ao76uTQA+DO8iAwil3mxrJ2N+/OeA5Ee+Z012y3OPm86vXSDR6VPVQGcpm4iJ99JRfz2S1Iw/pvghZT+UDs2xzUoWvYxLR6LYA75ACmVQL9rBxnUtwHasz5Wl4JPBhqf5MpiMOf1z+zfhofpb4q4E4qXO/Dxqxl6lDQTQWkxN8ICsGtoV+xP4d/LB/ctwNlSHBi2KjYeq914C4jwLcykKYCphZntl4WFoWBVMhalUEpAIjjr9PjIJZo/hnnl2fW+7xbQQCdKDlKXRFP035C3qjEBN/PJ/SIYjEsglaK8ET2gRyRAEDl5DJoCWBV6/8QdeXxDuqhnov9mA5MYMCNSlAJFI13B0iMJrnK/sMY9HxmXYhvNX0Ie493MmsIWQkKlnKUKvezsjQwdkUsU6a0YIMh+EUrEhORrKb+wobis80G8hb/yvVDSR/SUoLRqklv/Rzla3Bf3E5asjM+dFGUkEIZmTEinHPyWjMyF3vae4+0M0dy7YELtO3YJ6DLBzqNT72MXPLMALYDBjjuCKgKcTjwbQAAIABJREFUDIDlpGKpUapHDqKX6GmifaJz70U0O+2Rqg7AYaVsh3AcxFYw+HHKqCym2Xo8MLqa5ZbKSUAThuCrG7GzNFeM9efdl69f734+/ZSNq3MYFcNQeip4TQsOwGEqnln2QGU/kCwK1LS9Cjp/fLiL3gZoLhwldZ5MC6QXOgxJlAV63yfozjXkWbOdaj6BMzjwUbFg39BkU9xPHlO9FRi81Z1sdoCEThGlp7pNVc6Rot/RifmArKAImHDAWDVDtjM64+A0NjpvqMNEVg6cj62EU5bG6aCxHUepg5Ir/4jMITl8elnMQdqlnPHYRk4LttlxHeFNzFDk2bIDluswZl5tJasyNJjpRX5KPl/vNmZjmYqgAzU1d1PtEmy80Q6NbkK1Y5LAPG0HZ10XjwcGJl5r3m355p4u6RnTy3N+PGTcxbQRqPtZdw/HESuvqGze6xhgRfNqLAPVhHf+6rUCNqgzxXM6S0lJpbbHV5pOjb1KIdn2yIBBzQ3nJyul1FMtW/o5XEaVDgbZq0MgySrpd2NO3WCE+nZqwuYzS2t+5aBDf/qRUXHjMn5c9q9cAR2LWzMq/u1ncwkI5EItz2c2X1NzMxpVkSUATVUT7EZTdwzU54AHs0mNFEDVqdsa8nYKmzs2Bgq4sRm8Zib2aCP6OpR+KFeh9kvxf6YQ6d59OyuoVFTqV7yuly+AoqXIDzMXRptICWqcmPPkOwu03dPCQyuXk4bmKWK517MDkN6kTHNGhJLHBj+sJ4uyDKGgKAqpBBDNu/qvDCHajDZQobJJBWl7msYURIO+55gccYMoqVjLUBbVkA3pr67vp2gtR3n2+r4oyRSGoYwarunGpJShbUUW4JiWJqOdtgKwyDfWPtbJkfsZ/SunVjaIVZ3NeH7Mx9dHCQx48dPU6/vtmv+Vvs6mdxHFNfavoDJcqb4DGJbCaKYlejDGWLqyamfQ13efAKF+HvsJrreaZvhJ0EoJ9p5dZIxjfdN45sfvd84KbrEiOexIalVBRoViYBpFm44S1MtHLF2GYA5lcsZM9P0rnN3RH90o8imr18pp2TdJX56y7fvqOdrT0UAn5Wg0hCqytkeHGFyBMWhgQJHA4x5JUbLi1r/EdAhYh+Fb49pxffGOBIaFPrQJDqd/+Hw8b8sJmZ5RwLsXd6XR/gnOuwwtllcYiG9PDtnkezY893M/rcgAQHq43ZnTbqSS6pGXA9qAD42Yljo0WEDxbcn0BOPcMNBp8+H0TlCrvQurMNWutnPChotKdZiP2+HxvvM0NfSebu5i0WhAw2Ipy1rmkVfM8gPy68AcZ8Ax35WNfJUyLrB5AX2PzLdeWL6i1kcCDvDzmTkQ4PuW9TBp7NEp0r3xA/OUvo59ANAiDuvap3aSS7dM5iTrwGcV8LA+nzpcjK9H2uVW9ejDi+h773V/Rq5JlD1y1pDOZy+L0u/Z6xCgyubAnWaR8l/UPDMvTeZqfTzfW/hQlx+WGamHu1TghglbMvdaEdAmHCWpfgwBtEEnU4koZymmLq9ISaxJAsTOXJgzhWogPFunGe71FJbUqMzrAo35ucFSZ9wGGBUgZmQVRDTxFdgRowEAiGyEAnPjHme1EzQrvnyVvRWZJGUbVfRtwEwGxAFyR2R8AMmtRAzkGzK7wtYJ54lAM/SGoMMh/kW5N+n0sf4x9lDNwCNabz5cpGySdMg1wy0yr5k10cpUqQRIPDMe5tJSPr9xu6OqMX68xOUJx/2j1TJR/ASC0nGlE+fMka7HdPBJdh3lYn/6TE/MjIufcOR2J142ODZArRImcU2VD6Lek3L/lb3z0tmiwLTQpyJi3c8H8L5rlCzyx7gdINdoimWZwf24r5L3EUVPWp8COxTHZccHHIqiETsYsSvqKcJ5vEL/i5JgcYYxZjmiCBTX+fJez03vWZKZILLPcfwbjrKf6ouBjJCwfaEIMSDRJX2GQJGMNi+nGgLowkGFEmFq9A67UAEXoudwwESpWTjnFPHvknI908Z8jf0JxeNkmw86XeOTC72ab0/BbH62DOksCeielbEOUaInHDp2thmkZfADnWe2a62Xm7clv6FQZJUJrQXXlSUr6zjxDJsXxvu9bi5RRjpTsIpAZ+uY1kiHkyT+j2cha+uJzbXVxDttTjsJ0slaC5raKWhW3EIlN+kQddWM0dE/i4k+rqAPZIRIZsU7HMl+cngTP2PpL1fsgKMiMKmWJQe+r70hzXAu13JLznRlMGaD72Z/eEVMA6NNMY067WP3jKksPuAWyiBKm+6QXTWLf/9teQ18TjhWOnN7T9xSFo4im/wsGdwAie3efzx3r+yZ4jLg7tELXtWy72cNwXQBGrjQk09rYV539f3b99YoAuejrf78UfrpVxf1477/zhUQ8d7qqPj3iGBKDiUvMxlw1Ph8RqMbRThJyPT+FZzZrjwL2C2YcTcfLBjnhjjJzFRqqXHp/NXMG3JnAMUkiKRoMZJHZXycHdIiPL/AAUNmibgtMXYrQymIVI8OHnk5XLrHlS0ZzOy1BsU9t5uexk4oLir5EBfCiXI0pFqKnaKPoNhIOe21gO3tpvGkjAoD/jm2UOig8gz+XDZ1VVIBxWjOoYs0LP3ULMn7wbrbzjaQN170ZScKayJT6YSAUCpoOi0cPdUit9PoM/K0CTuwoyJrqzuy9xDpScW5IoBjfDAaWhqts0CiPBp+ZGCYjq0gE4hZQQQrzlDUsuax+14wSjuucVOyEj3jsyqxr5NVOSpGIJcbdLtZzmf26+vtfRxFL6VIkUacgp5lsQQOzYeg3sHndoVs76hgwjGX18puZ1nz+KgAarOO7xjAtWFJvZItM8vfa4AnpecETNDFK62zGecDxbSFwLXNHzmv4ThjZS0IeHAkO1jkdOM8PhvqBgw8LypeNKDjZ4jG2XK18UPzT0SgqTEjzouizE5KvZ/SKXd7bZ9YZdwPe95pi8vZbmqE5k9HivGj+C14RBgDyDAsCj6dLzi+Z2DkYt3OSrTlsqmZ4xlOdg5CMwF/tPHveqtr9Hbe5milXHyVLHRTSgO9lrmDg6Ov6Xyy+cC+rglaJXh8AzHpEj5nr2fs9m5UEXgFhy6+g08k7DQnnpn9ru55o7UbAWPieYwafPs5NfuySoN/0ogzUGQwafe8+YTXCbp9Zc/emRNdemNNOr/qqPirnBTLmZgnP58R09QUAFLOhXWth0jBGxeX8n51VGR0+1SeDz7Q7bNvc1SsfK4O4J9xVJymyxr8BG6KfYyZUh1MMF80XSGYSMqkmxa7bFDvZYG1bwFA1sENfLhXwsnJWGf/xo3TstFHR67Q9bccYwQrqf9GAF9hL0UUsYOY3nJUxBnntc9DCSWW0bFj2WU8Imqe4Gr/SS1e2SkB8Ndm3N89KKq9xBYbRAfIa+Ayxkmw/IWOigdF1Wt8iJ6GoyJ04ArSoq4R71NQWPJqUrFC2xTVzlr2D5/YL4OZ25Kv6MvikitVix2AHvh2y9qVPQdd0DXOJ00HLQgbT2/Mf4j4TQemFjHpUjI0ndPud9Kcld3nXwvufoth2zHqOH4A7KphLCOSuYdBRz5D5gmkVa3f/SNA36QxR4BHA+xPtmG5B1WyeZUJ8b4okxr7DaBdfaOYyRN7QTvYtqP7b4AfdecN5kJgD/urwDoAferJkWdS2Q+P8Q7ZhHZUIMs/Mw/Gs+XAQRGQ1s9ZFnWtnTXx7KBdNEVW827Y9Q+Pd//1X/+F79x3BHNR4E28x/00OBc2x4azRoC8o+WdGc8zwiyOtDVt205l9LDmQeex77Bx7UDZNyM/OSoGXVJOj+S1bkovLkXblWfl+/fv4FlofI8+Az/vfv/9HwwabFLG5YgYQMczGE4wZA25HLYcFWSHrFwR/2J+chabpjNAI3okCEOK8SR9Nkcds8j4M8i9KcMCjhA5LLxPpjOCsyw5vQs2CD5jrRnOgKdwvKiR86SHlk7cWGhjtsiGEe2H4wGO6XCsu1TdwJk9L8nDpqTCOhc/IOZR5Zlcpqp4B5WCU7ZUVqRAJh1tVgSGoa9OyQrbeskLJSwHbmFzozlukYUjW9CluNxXaMUBNwvQPkpeJz4KmrPDnBGX+ZM60uGRs8Pl+s2Tw7Vd7HJ5KEup/kTdQXF6btcHsbZzQ/DhHQdboNmSb45/R1tpY5J+7ET8yKj4ldX8uOe/eQV0KG52VPxMBkGvd3gSqaBknc0GsiLsZklANhA3T5XwEKBG14trzoSdIo9Eg0ONQINEM2huRwOYubzmVFak6D4z08CK4W+//TbUSA1lKn5YcYpi3A0G4zt+TiFuzzScDBmJ12Fdi8V12z1uGByIGgjFh/uFuq03lniwAUDFizU+rbQzTZdzlY2V/5Yhx6wL784olu2BaFHsE9BHZ3ifcz0hFEeD+yYsGmNY1RJEAhjprKEwhPEhYUusxqCSQbgR+epjyEhp5mPLsfSQGR27Q1jNavktaUbp6GpAyGZljiojnTvCOq53jeVolAcFhE/K30NFdaQkMyZouPz4ySZ9NrIB6raMihlmxnsXGMMAV5tdBw2OsMeeJe3BuK7KUPHpTgorGuGowPjMfvDvajR5ffpzdOymaGauJmlAtCgHFisX2Jjr7/AONK1wg8MtfGdBOHSGe3MxWhqY/1/uqFjev1dsdiva52IwxWP0WTJt73Z9B8BZ+c/oIRsaM0hygQzxnETUG/ka6EMG+1sCcch68PaOW5r8p+jATxXPaGQxOykGqpwcRAOwJp5gYKwr/ld0kN85eizhrv3MT9H3bzps9DjlxQwPB3dHSTou3GzEpeHSxmh+xvKPyq7M9dHRTuW6l3Lwq1e6nQ1QG7kZDfoWMeQcMYvt1QNpDJ7P3eXmmQgHXSOxhh4mdf9EfskEGStQzcEJ6v1Vjorgp46U3vGElb9yxAfD6LDWBlGWr4lMHNZcNaumMndbHnPDHi8zuTLitnxnLiU2vnTn8LQc6Xwz7trR5i2Oir2jQ7pIywZ2dDOnMTK4fQJL6RC7PZqdEDnXmXdehi+cN2nQC9raW/Z7zbJhtXS50xNp2FumF4iH5yhqE7wIfQDcP6A89y7fyj0hIEMefZabVyR4IjXYQdIfnI1GeaPsV4HN8WyXKLGsYABOAdfb97esYgJvskMEXhlINwCLLI1JBo+FseotRYsExUI3i/FEMBIDCFguy06ImFPU9g8WG9m+GZEN3TdswSj1RrkQJBDXYo8QLc2skPxJ21PkrewK7NUn6tBR9x50kFumZs2waZhJ4Od3fgptEDJLwVDIrhi5B4KGWh+CThVJX5MTHVkJXaeUDYwAtbaP4YCgH2O0Zzh3jokgm/UQlwNiJLuj7O2wiDnGvna2neO4c0S/M3sUwR1Ny9Ne5GknWLun8hipAwMB1oY+9hhBKGGXK/Mny61Fj5ynu08PAXDX/pinRLk1OMOUye8zywC1R51XrgL5Kpt/gx5FF4+Pn+nAbWWZPHKfrz4TQOvhDEGvDGbbh+MF9pLEUDhcEBRjJ0z8DsCWGTrm33TkubIDr4kfBApq/5lBxMAUgOxR3in6b4RDBKXOCqzvkd3kFcwucB8Xg+xxXc86WXaq9YZZefzK1+J55o/O5oi/nb1gfc/zdj+Zvs52FlmvNQgfa4x9sP6o+Zoufb0bsDsTB7yglULqMtMy1WsUpBpjxb2zU1Fsg7RaDcMjW+1RPXDgIFHgUGaBdCaUIK7q30k2WGZFhk88L9ejL3pb7r7ycBq2BtrOhDpmz+a8GpCtJuQxf/O4jn2Uo5lvzmkcznbp09Qz2AdK2RvKOqAat4YqrDqXFiHxHepUMaYI7oV8CNxK2S1/xlEBXiCcxj2q+giTNvce4bMNfiXoNw4xBopWWUjwM+smAz1NAWJeKjsoFdy6e/0pK/mEI7wxhZU9xCeWebHnHz0q3ruEH9f/96+AWOuNjor/+e+Ras1RpsBSdQt6Tgt4ZvS5basRIDzZtIhEDeYc9ZZV069Hpc7rg+fgHfX8BauaomiDwcEzHSBzpuVJ6RfYiFTZiDx5er778uULIkl6fwRWxDVY7LqmVIrgSVezbyrXrkl6yiTxJDi7BBNza17vovQTgETVYqVbfU8tAEK6Eg2mVF5Up9pS8SM4aOdNx21odsV/joCCuFTGjBj2veotGnLXmGbn0MlREbq6sC9FzZCuXNpJK9ImWuUlQui6Xm9c0EtwzXpEOkugAFuoq7+IJ+3IAKRZrj8z+OD9CLoPYDXqnua5sLKmJm52hMXyfP7yicr4AEjSIMto+ubsgfKrdE07z+w4KuE1GV9bM3y9pmb5fqN9ACTyQf0dpBXvYRibVkAZjVWlEtZ95ieo6bs4D2xI9D3iarphF15rR9afcFSMTook7ok42pynwXqPd/R0OL7iZZqj+YFxPs+rHf69ETyuaHfiwVANw1FRp3snzp63zGcgDTqBTS7/5MaBAz+bXFGdfsCTgxc9VnNN7v8xdmzFmeysnMubDFPhKUuqbJtQgN0qS3D9zrBpn5vmshkfDDjMwv+/XVTsBwCXJqhs3G7uSENr+o4gCcc+gprjhQa0/Ck4vAS113vrqGgIXTr2IyJLpT5AhwMQ3d4b8gsD62MpCjhxH9b5ZnSwIzj3lLn7dF/6qdK1xSN0a52jtobiPwY5+/C5tfuIxx2Bxb2sKsmn2NAaHc7TXmFN54Ur+Q7kpZdJAOAjmrtxod7P+Q8PPil15MxtSfT7xhi+deRbMjoy1N143++ocH15ni/t4YRaz58vTm47rtVg0/ph8aMG9uEdBTqOh0d1lY8cJZ+4XDFAEN78FkyS31v/PK3rAbHPR04OIjt4gn91p8UOeEIkLpQ2lyVS6R33jJJDokBaygo7KqjvMrjG0ZbVV4CA4g7krMU6TvpojlhbdkYFaBmALEuYsmkvewMAJI3SIMogdJnZKzAiQbvkB7RjHFlUTg9G5zsSvhOAZ0V+NgYQxcSelDnuyHKWH6GDInvXZT39AOHhxRgioJ9+uleOsiL0PQBN6WKzI7AChzhClEiJ/6Lp8Wdmb4BuVPLUjZtRsicyL7IpKoFKZxWQRaMbXpYYmg9E7Ru/8R7E5+j706KPcUGeS1J6guo6D9xL7r17lQCkm0lKNh3G+lz14q1T2UngALKxR8V68KMEvG0S2NEGSuVoCOAbcjsAe9lrO95Pu/CVpZxFs25ofv/A1Uo6fSU4HPYyfXIOs7KuTEeHz6adSTh/LcPf59bZQtFk2/OH40flgNw/wvvkM7wrl8e5suRYZC5xs1SeFA2fqxwW+sfI2elM/aQFsGE6GxAljmd+YrZFnJmw5ZBZ8Nj4FdU59PJQ/5FaJzldpnKX5kngk3amHnnsCiQnRbR7Oj/hNHhf6OnIcOg4TgNceQ0zgtEbcSibV3zWtIr3yHlnDbuJFgLY6jPhhuIMjtRVyoKw08dzSceOKxNc6eDm6XL+wMY2bxJW4Pmvelyn6XCgVOlv9qBJNd5Moh3Aetp8nnqPDeIy0hd3wRO2dbSALmftig3VL5VYDjKDlKUycAOVMtupBub7sexZAt0BurpBU3Wk0VjGYMc8Ux+qXg92xI/0sdc0TzIP5QZVehBHV+/OAOA2FjgqLspt7s5G8fLdSumzKVuHoI36MMphCZ6rPiRdfvQ4CIytlbjznm7ffFDIj+t0EaST+tFEb64kD1L7cFRcEMDHV3+TFbA14sgOAiZIcXp5unt9frp7ef559/L0/e7557e7/9UcFY6AIMaidLvnJyhCiAaR0js2XDbLiRO/GgNQYJXjT0dIq3u3OcCOhinUVyADOIZ0k/YaPl99JKC32EPfhI1KYVjRA/iWgHOVrUETNNXGdV1GR9M/38n774h6zGU/ZyuiqfQOIrBKiFhJggKHxnqVLtyJ6eSocLqtlTLusftUdJzMAtWKuEo/AeTX+hrvv6cQLweH7tmAgb0El1c70lyphFLJDsU4fjhWlQkS4Dc6UVb5uU3ltBlno2xyaKXxpwWEMnXwALn5Hy7NKDPOFw1NlXJu4eA6nGl0S1GMaIMXZ1RIK4i1YT+XUiZNyQwaYzRQKCbM0CAIWsJrPUvrcamz4e8MpHodtsrNKfKwvyBfb0Cy00qax3LiERjF7S5dQq1hfL01puFj/mGFq26wYVQKPO15r6l5QX+YX9BV6qKrrZPCm9/GW+BUczL+Ce7ewS6DO10BSqeDwbJmXM+vxZlozfj8fTgqaldkiE1lpnxtH09XBq30+9wNEbPdUaoHLcbBNO7YBWZ32dnNG88KWj3RwPzIh+bvR18AKW49N1OqzkqZdnZOvIQXsi5v/Avju6Xb757rNe5GKteVUbjb83ihmM57dibDOkcE1nz+yqCcx+Yx0ShVnWE5Ee4jAwaAUGsaS6aiTWz9olJY66x2wzqBH77Da4jyKQd5d57j244Kg6HOqivvl3mlGukqGttOAdAl/ufCUTEDtTxmo+DCmQs6WRtg4/kb8rQMLq7lklRqyLm7pzlG5vU62EXXHGx7U494breL1xjAaMrCnr5NMpvpv7v9xmEWMZYTXylxNy4koulabXcb+85GqnNkvrV/eTqo3NNlkz1KVkL5VP7L4tjmvXsCmWVcjWPWoTrctcs4vSKCE92kcVzMCL8ZfOa5jjHqX4AmtkP4b6eVlMNZcvUFILwzceNJwRt6ZHJ3VJiBOxq685G5dMY10Rd2c7pu1CQ4L0f5WnY6otlBUNHLYQzM2T+dmQG0s7iearSbsTeV/RAj7bXe5ydir52h0MDCqEAEUFLAbZStiX37BP2WJQ3ttADQK4dHNUCOTAtGy4d98fCgcpDoO6UGsZNuYLDZtEzgJ8bxzBJPn0oO2hkTzwI9ofcHy4kZzA7bgd/ZUcD8EPcu2PG/gZabPCpwlSWm6rru6CxZGnMhSMdSTZk1pKj88d28j447Zsz3eRC8p3wxv2Lj6B2DVxCbS/w66l/gs8uv+P29tM6yHlGmJxoTowwS1562cID0ZMpc394nr5Ur9YG7u8dzEHimzIag2dDvEPz3HPsL7wqoCnur5sTdUcE0CJWOavaC95i8gxyDfUn4p2kz5uFeNqDdOBvPz2wGrp94BHpY/GBpKwD56GPBjBhnIzgLIObk8r7ODInzFjyGegGBbmcBxL8x53gOouyVHRCyP85Yd+JiXRX9f+axF4WfWynRvF9OAjgdosSSMg2wxwKDszTfnbNaquQYbU4HjVVJLWatPHJeKlsI2dUyDTu9Ws910CeaRmu86NWjrBaW43YvHjndesR/3zjJ8nC8RBZLzDmehYwRNWo3HWeG0rS+oxzg2QafBSZBm3vITnvDSY9z3Uodeh88r90ZtmMueJ7L6BLgJiIR8iJLOkk3Br3p4cZQwsvi98xnO5yP3bkd/MUl+ujYl7NTD7Uc7nTUn4nxCVPDsYtzp71Dhr0uDhp5eq6MlPkZO4mHc2Ant8o+msd3OzSdnxF8fBLMk+KT87lSKCcnhQPBaJNUeTL3b0k0AcJr1S9pa3CAV6WfTlP4NUfF2EsQ70bJxgpU+HBUnFb84/O/0QrYQLjdUcHBU1hlpIMiOOh97t/t8Ee0zNYajFCR7XhELTxENIbqTbYUZhtwUDpCyUMkdfxuZcZgiXOxc8TUYeSowCwMOmk+oQBbqWFNSvZHgHqjhnhMg2akDgSSmkWF0LWj4uWeqaf2tDK2C3Wqau+7FqLlGASYvkfDOEVuwCALxQINr5U6rGgGR49lFFmL/ONcme0R77ATpgsaW4e1r651aNDZRoqZMCPYYwm9PSk0N46KCg4tcYIIeDlL6NxyfVk26KNh5shkjUcR04OAdi+OAfRSVJ6kLRw008kzKOhMBkTAheGzEXn2itN7H0aYDEbUgP2UAFRGtqF+KdRnRnyhxuIznDCiIKvJIErKtzn6msrhD+x31eNl07zevFT01QCpVcnlrGj00FmQSv7W+LmI2tlyMIN7/nKqj6xG11YyqNBXg8RuqFKgLo1N2ltnSIB8huvH73iWis80+CN5j1aj/S1e0UqJmXv45RlZKD5Y4/YVR3XpyPcdlVHjrkt3joLZgbFhJebSNcq2x4ujwm7UGVxtf+8UpTTko28MSgCVops71Brb93HOzyPvV9k0KKaUMwUe9+Wb15hAuHkfn934TLt8ONsn72dtdp7r4Y0bEFpEN2Szgb+4TN1u9+1smgyfrojPt/V1M92M2RTj2nT6GafF60Yg9OCo0IVJp5OjIgApGqpBA5ITTf7UmntszdCejT6tCZ5iZ89sKB5PUn3h/jfDpa3hMc5QHtnROV9nvprWU37XPeRfB0fFgT52plSu6cb43TeV7nUfepQAwjrOxlqTDV1HOIEhO2M6aW970+lJXM08kY3mT5zy1Ew7kcL2qmQTOxl2yNogOR/GW1bsTDopHOKdqNkfeoDkDP9pMxpK1TS6lPZrJ9ma6t9lW3dUdNqmrDuClpdzIE/t+gb1lBr7LZL/uNu7dc3sxirZmWDKtGbJo5pMwhkRD+pyxSBXjNyAGfa1ZVRYpkZ0M3md+7qoqfAlL6lZnsglb09bwgES5KXxU5nbvJqA4Z16ADBK2/YFMyHMgVT6SFHs8TSDbg7wKRnJmwxwRwYHnRpFQ54/nBTSY+loiyhujhvrpElRt6fTwQc49PQYo6PMux3IDALNUZl28XzXs49vhtInWjM7Kzy+ytZHruUC5OY8CE/jhbEeLMnDHh6cE8HrSpJWGaiM/HdpKPEoT9wlfTMK3M6TclDYiWA9k70xXNaL/MXlXiIjv8vhuseZQnRAxXI4QAsAufeo8ZiRDhuvUJN106OB8uenaDLMssEj7Vj+d32ZNnTYXnBQRTaLasOjBJJUetv95hnMCKUuYV2E54w2sBuaB9Aa9hUAadlHDk4DOBulrQD2a0xBmy7nBtlbNi/PPrNsrC/F8w2cYoy4P2iadmX8X6wFMzSbA0y2Jhxj6qMTjgjsSdyvxsimX5zXVn44eBkEjAh/AAAgAElEQVT6XijSPeS8HRmfv3y5+xkZHZZ7snHD+Rd2XFyHs/qJwG6SYNd5JuYTuvYQANc1ZV3bz1k8F2dDjpL43SW2Eq/xOoqA4hVsVq8QS+liXoNOT+y1Q1wh+bcVy7Y/lrvVb4jAts9uOBuGsy+MZQ1SEbZD5o65xRrDKaVnZLlAZajE30FbwD/sqJjGqMepL849s2Skh+JeTc5ru9NfZlvMf1dw3higU4EL3J+gI+AJ0teAiyD7RZk8d3QkxrkM51pNQVlZrZyWZQP1aOJkKE0WvOkzHZFPP3nezJ+6TtF1pEHei8Z2jopy7MkJZb4MOVQlwnlmyxk7i+GeSeKyV8S9KiDQtMu9qWoZ3LQLO9zjPzkq/D0JtjLQ4kyIb5G/lKznfkmv1GIRw+A4Uk99w1HhNXc/0sJLVgdIxw3m9ePQmQ3pn9xb9HwVtvqRUbFbuo/P/l4r4BN1u6OiM7RgmFSwnDEwzo4HlSZqvw8KDbyxapDXGgcDcMq/zdiqNq2VBAj5pyd4B+FJlyIG58LUeNAKFQzMZDtkMrQvFTly/3D3I2oR3jNKHk24IAwMwIyOF2eOxHygJKnnQbhPFuZwbCJeVvwgJNRwB46SySrEn3YIZQ3QAPnoWFnfrVrKUvxoH1yly+mFqTkRfHJTberNqVItMqEbvbh2BhZygKNAsWyxwhhjZGbCqVSDjDOtBft2lKMs6MIpjgaa3jp/Oa1mLPZ7BiM+0ZcygBnVQ6FpIJc1XvkT/g1Xp6UwqZRJ+SnqdZBN93dPelZXDOjcsMJW5wvzrbK3beirYeJ3o56mJ95K51DAXgj8zWISUEjR3K5Y017j/JfyUo02B9ocXt9pe3x5jDMymcY3k25tvJfcLqKcseru0EjAoIFr1j2YmbSb57heM7DcR70HmvYU6jVxJOlIk00d6QCseUhOUsdYDlvyvvP+duN6x1NMv7sRd5DGJHEEB0Ey+3HU8Ma9t3NxplHyiiTCgWGfsq58Xud5pAPAa9r+5dlzuaPicVBWJ+dEYxPDK45g31tMato3l0rc3bYCJOnLw+VFzwXG7DHf4sEJ9jXgaZzLvJfTmegC4Za56pp8RzMkTvT70tDuLWW1SZIb7HajGRkTfdIoaY6BbpAc5nQEO49nsCCbhTbxsLdM5bprKDEl9oeo06YvDLypGV5e4zTO3jyrgwiTsdd4TQJao/xP/rCZFrION1uULHhPtO+ktJnQ6p3IKFJkHwJkVG6An+m+eQy7ATeMZd7TwrprogZlabB2eUPutP600mDT913WVVCEAI5dcAY5xA0n9O1LTk8Z5GMJmaSZ05MzOtVNtsXI4PhxiSiVS6U+KVujgamXDhnbKIstcpKXDaSzY+GiHMX9wRsHm0oAYYC6AHoVSR+lkI7roV4VLGnzrKj4iBon32ZwEuuSvwqYBTWJpsIlEv0GHhQYlQCJdE9nrDjoJkYSJX+Y3dLLzUZGAfXwHX+aZ2B5eWSBudzkd2k74rCMPCH4VMwh9jWi8tEI/PHT3U/1dWDJXzWSjTUQKM9eigal+Ktf6/HG3wTFy7ZDeRxdyH4ELKXrElcBdMbehfPEYKuzIljW1Pb3SlPkufy+sxGfF5bDKp7gTIGI3Dcg2xtYc68rQ9C8jBkdzoIpm3DR1UB7yvDwgHRGXJILz0+WMfZeOsq+gaDpSPihZt5hezMgUXLqNfY3ynFJLuN9XAfa30WHmFM4RVDyitUZkl/Oy60MDPYV6E17BfUiwp5Olx657x4mBsXd26HWlmUr44fZAw5sNM8VuClAfgA1dTjd8JpESbvS1SpcEcJnlbRimuG/qR/pHMfUHajYMwVAbbqGWUHjc7qTy/uRVQNsx6aDiWO1zZJnqxFBjCszc5qDozucQXHuTdElUSvz5PKgO77o+8niCpylPVh8MXV2yTuvp51cOMfO4lO2Tcw95uDskIWkDgRvvZE8hsGCsa3nEqAqVa4G9uzdVw7/eE7MB86ie/bZjHe42XtmMKm5d+kYeVDJ7Q5i7WSzXfVSKHWoHhrnk4GoY3BP3wvzXa4Ry/ox66p4V6x5zxCLM/7Htz+QsYSM183PMIdB0FTGWme0JymLHqLZkN3OhwpmWl49YSn9+9P6+Ro7KpDN5D4wLVPDc9rZP286MNpef2RUbEnm48O/1wpYUbrNUfGf/4NKKVM66aDggZHR3E44lAIoN/yujKyuUFCZBfN8Ud28e6UlKeUthZnKLIG9RqosygOxcVUcTDorCB4wVZNK5BxHjzZ6HVQID7u4dAh+R+NYyUG6XQiT1Fg789X8y61N5XMx/j3n690vAKjKKAD3njgnBTAbLFEG01h2NH8yu8aUwxuN2pr6geFhBWnDYVF/NuMgZYTZuEol2ory+ICTo2KQhX5GB4xsL8igAJPWWtpgr7mt70Sava6HkQKjS9fp2Tm2g2X0Zx0V2EO90krIY6TAS9hGppDUeV6Vjgo5LbqJJEdFOOPGvXWzOSsbcpIJPNs37OKo+J0cKVLwGWFSCsRJUL+Pd40ZFeWQyB1U9JMVWinQiuaKsmB9i7YCeSKGpVUiGEtzVGBicxN2b0PNetYxPQ5wK/zRM0H4zONPX8zpMkd/kQ7SLL2EHzt94TaQwuhO6q8hbxOP1db7vr6ms3Izr/dJMToqstOq7Gnydooaxqo5pUILJjkqjB5XNgp8wylzOZLmoCC/bZH2Df2D8WN24xrEUrpPFGIuO7//BNxkpCAiw+TyPCjo8zMdxQiDOc4ZHMGMGiQfmp084xMYOVn1tIufzHDmPNvx71sitrf70Q5mX+fdtZlR0eWLDfnpMx6/HdcTIIIXrDu4dSOMluAwtNNZOTlb9nzYQrIdZo3val2H8y0M7FZHRZZ30/pfddua9wJSxRHMRAwSPOW1G9Qoz1Q9rV/Vf8812h2wC6fAct70QT7PqnESGukeZ0QO4AJtqwRCf+52vy+Ea6eDLoNIUl2PrujlcR7X587jBwgFcITXW32d1+TEm/Km29n30d/heMVFNzxkw5CExj5sdhp3Gk/ZGrwuMolRp5xZrs5unZtN53Ry790rw9kXb2lGWk8h6Kd1pdDeSwRm6bCxth0VCD4JZ8CGR3HOCvxqTpV0QFPxhF4Mhw0AQmWdtCEEKQAARXY655nyxXy/9waBk1MAnuSvx4LSNgjaGucYwTCcg3lXfO8+d/v1cKYCt928o4LLmsDFmAPIjnuizInrnP/4yV4BLp365ctXOVO448hiwKOdfULZGuuVeo9YVZl6XKP43mVi0K8AmeucI3o3KDguGjrHdVH6FeVWXgNU5PrtZMvIC4ruXLaJToHiCXBiyVHy/ft3An2ZUSNG6CVuvZK4ArQvaH8K1B8YoQSG1oh3FHPlmkRzbGUAIdvM87Jz4w1moWwSlhlTHwfxJoPkKM10d5elo5hZXj0wMC4D7CIM2r3KkgeNz5na3FhQIuice0pg+vHu8ZMxDoOnKonkHg8qXxS0gxI3P+kYcSlg063LqblXCOmOmT/42ekkqZON2XOuMR+3wXlmR+YE4HfHB+bnDIWpKoR7OWAOchoEDpKOeel8vt84hUHbyoJgVhG/70F4DJ4Lm849UobyROqhadvdVS28Nujl0zK2nUVTPGFPW9Bxw/n6+MhySq8sa8XBoJxD6iPxN+mX6+l5hKMr3m/7hbhJZM+4bFVlB6e8v3BQ20GSDtOsInGyELSO6ayrsqjoIfMazliWu/Mz3WQ7eHnwPFZ8aNkL6czyur1fI591m2Qt4hvxd5/R8+sz+KExJ/ZJIY5oZ7r3s2xNZpPEOadDg5zHJaHozKCT5svnz9tAFvKE5hxZHBVt7l6XU3CGgkPdX6cHpW41g19wVADXVAl06zPYR8gW9rfqDuhlH1KnO+sqXSx/OCrekEsfX/8dVsAa+W2Oiv/1b9/BfnoEBpmLTdeJ2Q4y2N8VyGdjDAcSMkMKuWtxKsXSNR3xLvWVCMHjSCOkacbfyIBQySYoz3d36P/VmFM4Kcq45ZgCzIPwIx8kQ5CyAeHdtyqNbQnkxo4d+Q8ZOABjZtte73GdEvBQunK+zoqzPig9k88jw5pqjDemPAIg9wDuWRtUdSpbnduVGqliU9y85ahgxokjVnaOisUQlYI8KGjtImSrhCJ3yBBZIv2lGLkkE7JhrERujtrJSP0VR0Vm7LT9s+JrYYqdUjSAsgdFbzQC4EDrjbwbyOJax57G4OoASY1NVVnPeJ70GPVm4wT0r6wVbsko4N4yzde3zCoKr7CBOjqKOEiUG3iJaLSoocmcp1CuormjlRfN0lSzmZ7r9Pqw8NkubUDjsfMeRmGNP2V8zkCRxzGU+sDEBrfThtLOH9VayHafANP5zOxHS8dr/65xWs1fYzBNLfxpHOMOOH2vo6I/EWb7IcIoafqAzO/ea67t59p502k1o6LyuQZHbtiiaSy5tvq8OypMQwR/rKVXHV8289wjph7v7owdHRUCVVAIYWAk+3nZMILRqdIIjgan4juWMowzMkc9+cl0xHAdHcm2n8NMqTsjbM9ZjvzmQD9bWsWAOa/5DHU6HL8jlxp+BqDtYg7zZr1B6zdQYPK59VqNww7nvGAPZPbzlXOnyGE03yGjou95d1S8x0nhFaVeRDWsgFWDAZ2z847TSfVeQ6drPypjvl3WW7eidKtcsSlcW0BPxKHIcI4rHUhj+fDm3h6N19n53WRxLJwBtuYYXZ2/1+eug9qeA8Z/CFgBfz1N6NaFTUI68Kf5Df0sbd4BrTRB1ToL8XmPrk2+kPXiqfcmyHaeGQdq8F+R2v77xBvn2ZXTdz/v+9fTSWIkqbPkANRTzdiOGKSh7J6Ips3So2oWbAc0wJ1e53zD7ggu86ccPWokHCVJorZ9PEPZKQFmIgvjgaA7AUuCY5SRk50DMvY7KmCEsvpAHzLKykHAY1kBTCr5AR0IkWl0uITTQiA1Iv4FaIWN4gx8gv2UEenEC+cEdGI6dPBd8EhlosSzw45y6TfXlKf9GSWxnHnBbHCc0QcCpLE/EfnL0i2MDOZ+rZM/OSoYvKWskEFJvQPwF2MNQHAE+8tR4XnCvpWTJMYVaxU/VWrXunCZzwOcOag7BEHZx0N8LHSFDHYrLnJkG/exRk+w4x08EXNFhYPISICjib0f4/dwxjibjThA6ZjxOfSal8gS8n4xMIPEPWrL3VazjQARifJdj3ffvn3D81zGyX0D7AyyozSuiTngvIpHJbCofgOBVTiKnIF15QhZ9Pse+OJxN9vOul2n4Z45YB2Y53l0VOD4O+gkxv3jB8Ztmg1HI/pg2vnRHCtdhzI9+nmjHGxl5xxMYyeGSj4HPaIckbgbHCSqkIDvmhMmaNPv8dxdWWLHPQLXQTN3g/xph/SVfmWZaZUPpCO7sv+NI8T37jfkSglwMrZofwfx9HVf5IKB85ZFgZKp5l/zDQ54AkBW54wO5RdmjbkElJzMnbwz26jR2V5WvdPSny4v/UkoEIiy1vnHz+8C2h+qr5B78CjAuNMOS39TDsd5j/UJh0R85qxB+puIR8Ip3J7X57h1VGSK7i84KlqwFrAYyeiFBn/BUZFN0i13pIfMNiToxZmMu607BHrg/DTy/3BU7PWOj0//VisgCveBUuTMqZn2f/zzp5REKwvfVP9Sk+oHptCyNmOofa1e52Yx4OhWCZfW/ADMvyloAUJDIQ5lUI2LLDRtkMyOCvC9iCjyawuBYlrmM1Ng0yBWU/CHjYIjHpqGDyWomQBT8+qH885IooWxGFiW06EZo9ZL8LQGlIU4GNLHUE+2DJVRYaCqYi92rOWXz1+gHDjFk4/mmKH0xSqlVtkcFTkGmrH8U5Eovr8p3hkwwifnknA1qoZfm16ONY01KTEE6Kf4cS0rjY5qQotIiBBeoqU5ZsAOjUUv8N5oqLNDZFbWoajkuuVNQz3Y3ogMKaMJDtV6sGbwOJoEAZVR0RUg0oXAKSgFjJ2HIb+tnV6OCjY5rAhqCPgaeiPbXkbiNsbFtVgNL949Gwq8DplRcFRUqS5EXwyGc71/C2Rp/50tlfRvFod/3cizRZF60dr4OshQAU+cF7fOzkE7KrYjenPBrhwVxZp0VeMJbSW55xtg3Q6aYSfM5xX5tnP29UEbrBjA3eldVw4IcIgbAa0d4Ix56v7+PeckgN1K4wSqdUdFOvaOZFl02fnscCAPSIrHlYaTx6uMwAKH9y9/bywTFWOOt7/7tH7DforvvDwzQq/S+V3SoiLhTsRLZ0Wd8ORRww3zXHdz3xtGR3Np5zk8cBo+Y3JUTOenBJHHRnk2/LzlqNhO650G3wWXKNqYdQmD2OsATm83QEXCuc1RMTv78PeN59nT4qqWUCWg5GjLKl1yhU97lqbxYTWkc53bmt+6H3qqHEB5l+YbIAlBKNaejx/UWleUfj+Pl4z/ylGxFcLarnbmMTaV6RjftaGTdoHXPV4T8jX+ZWaVe22sI79oF7+d5rHs84VjYLtDBzqDzooSpyrlpFGkGO+8cco0wB41x8NeT9IDZ0eFZNG5ZENXHPk7h7Knv/tX1j/f/QSdo3ySDotUl1ZQtu4yQEsgn6BN/CDKXyCjy+Ag+hZOkKmXjUENZZtwjRitnkFpAvtYDleNnxX5XhHVlAwJXl44KhDcpk17y/nT19E0XO8kzef/hlMAfRnoBAjd+wnNqhmRG0A4MyXYbBu1+uP+cL4ARFRvEXlGTCNxzuGwRZTyT5x7Z1TF++EsStukdDY4AiOTBJNwVpaCklIGr3x8J652cp9lYKTzC7hiSS7WbTeY5ShgO+rijaxXz0bS8WyXkrJDc6bd8Uj6xDFTx/RnEB8ZBUGxyvToz9oebQC+lNmo2BD2TO89ib0punfwonvGJXArx0821sZZCCfHzwpGlO7UnZnOoPD5CafEj+8/dARfshoBI7zrbMXv3VER54OBfZV5Gs9ks+ooR8asEADsrQzTjg90/bnGSjrbAfUOKEC5MYDvypCgNzNfMegCWguX1MJ8BID361zmCXQiEBl9OXWOEQBp3CaFufVUroevycw2ZSMlPai0lvtdxBnvMhaBFWbPLXtEJtm6hOLhWnA6j1IHLhni8lro5aCMCp8T7JtKi7ucEhxUMTbYrewFlHw3zlL2ddkMSdk64NHBRwf5vMqKeBcCNgO/saMGTnmOldhXgfTOrCCewMoj3fEyjyje3zNUjkJp+uJkSi3iTlN6+HSP84QenXCMsVm9e2VW78fiK+DdcITzOjhizdMUuMF9Im9myUHJXRGVdaVG/CIHe1rf56iYg9EYwHBobv8LjgpnNMa/Di7oerhlwNEm7/M+bOaHo+JWKv+47m+yAuIiNzoqIqPChyaiayLawdEL5BClMvJPR1Xo88SDoBo2wKU1tnpVI7QQdtlDQin3LTIgmBybDEkpRxZEKeqhH6WB2wzA7qgosVB9DT6pTI+9tAC8vVvNmrYnlYpZA3QF8qfZgntqJLdufDfcCwjXOkrvsMBkJAsjsbrSv0blOPqITfKovxig6ZkZMeT4XNE+ydlkDmg6iEfC7zRQ0p8zOSo6IDoI5oOjAgaFosNgkGwY/g5kxXoouweRNKF0WXJOz/j/wlHRnRaI+FIqftbGdwQzFK7eCJUmTnq66ljqWDEVenFUKJ3TTgs7st5yVHifnE5Jo1jye4rOvxXmySNyoHXugxTXfFk5V7qCg/koDXdQiHQosA6LxsVPolE096F4TtIlSqSRzrvSy0cZXLByPZ7Z2eFmwK3duodNU7P2W+r5J0cFFe8ydodHdKC4vCjePBxbK+7zuTOfiGdjnaaf/tEJ+J4/PzkiHL3WaXY2kPrrf8VRUZzH3lXtoUAlRmYJELmF8U4lnlyyZr61AwYY9wwaCuSwys3tPKr2W7/eaV0dKdifeeUMSqeogCycEZWuKaCIK3kFrHkNBgO5wXAjn5jn+gaxvbU3k3PkGH7bnsMa4DoWp+cPe7LjdL1B3zoHOvT1M0c/vjWnG75fnVjDCd0+4cSvZx3Fkb9XGRWLs0/9j3aUXCdvHFZxfeoI0NEABnS9ozl+E+Ct5xQnPmQm9SzZZVVulWB6ixwVJRGStQ4ADXio6rv7laszdd2i42hkNydJOiDEZ6yEGB96jJgrPWxmLHQyUvfg4wcOdaCn/YiPdHb44tIh2wF5zQ2D2fHMLCPG/UpdwOWgnLmjII4EaKUUYA2kS7k87Dxxn5Wdo+7Ma9kctP8YnN4u7Ms+owKAjQKOWLecHe+wRBcihAB+K9+JCrRllwBo7HW/x4GCj7nnXrzfpWGdvYIM9ucnyA7X6w8ZH7pjAHXMHHS0q5pvL44KdBTQ1iorYOAFm/OS5QhPpZ/aokj3C5st7FNnC0XpJ5a9dQPXAlsD1GVfCWaXOaio96EJ2mWEufRHBddYJ2fTctUvl27PCOkKHKJOThsN6/fMCO03JNQx0CPlsI5xjNFzRvTxzx9sBtx6ASA4QXY19qtFuaPsjcBN84XuUCh9d07tqb4UdgIGkB2g4qfPQeN0YohpmXWtG21Ri4buoimA4gG2slqCbe3oExGZKVHWhwFpLO3jM+DsGc6XDg8HNbrMl4For38PcjSN1/7GM5jhHy9xo3KyqPGM0VFRn8GKVtYaM2AZCR/3ufSXs1pzUQw2TjoFllE83L97HpCmXmiB+MMcWzkiXBu012xiXKtqFQTHOUbyV5ZCsz3hvhtBS2v5aJepYqR5OS96Kd/Gu+2gEi+hXlKOr5gys5sm+/ctOSGnozGS/oy4FXzNWRSNGnspLey5HLNBcwD+xZtNA2Hm22kRvNB9FeywmwkdwaQkVAaWet4Mf9uICupK2AdlCYGPwVEfWUN0pLiUlvmCr41ePSx3NepYGfQqHrUV2y2bZhnYdMMy8sY8IBc+sURTOFGDlmJMLI3nYFnqh+YTdgRz7HXOejCu6ZOOolhT8ZoE6zf6YtrM73dURF8pnzva5xfZFKDPHqQzruBVjw/MN7PfeQ5Zbp+ln8hHtFKt7O+VHTiI+y4yP5ppb9Wzjw//VisgbnOjo+J//x+MwIjohFCKIjIb0dDJlGZ2FYpp9XcoVkSNEvcpdQ6NddXqmjX9g4ExjAKMLuoEZhmN17tPoYjK6AhGFUwQyuiLFDYpFQP7D4AyIn5a3wePyUIjIo7ijTGvz4+f756ef0I4+We0ndygTz0Eem3G3p9ItaAWkK9Dm4mJFLyCVbLBqsh9MGd5walAMLqDjeLu716Uwhs2wkMwVinvoWjHvEK5oKda3ufmmTbCCwW796iYG5Nqmwm2l8TSdo4it2UcSKcufWxyVBhgdjPtjAhxmYqGG0HfxuZRvLsuKNYLym6UfooIfY/PWR/8+1cdFZQ/dW66c4IStSjO1yFLR2NkqqL6sEjaTHo8HsPP9L8AQkdFzVZrZmLoHEEJSwVjPI9uem+DM85wrFco+/3HRlaN4FeYVjfEoRqP72hzR48Vgw4W0DM4SW2Fq6I9HWbn73IPfD3LZiBxFmsUxttICx5YB6A7yFNnPmPzi4ZzWnsUwUB2rqXHLgenaUYaEJ+bgDlpyQpZGSrkC8SadMZlFveePLPii/kJRJ/aiOV7k8/pl5ln3eKosHFmMM0G05Wj4i0KW0BAg0Ji4Am5cZFQKYX7TePwzZ/uGBKIVynDdiTyKZnxpxR1G37Bi8v529Xui7cfhnZSOncZFVdzY/+JSvO3F8tNZ2PsNkLDOA3j0tGqu+faYDSNNu7aLp8ntZnkYd57U62h1w3AveJPrsOfLsu0gbqWzt9JOztTTVS1PeMtG3CKYrqB2t4kR85tHlN/8v4tW4NTEjlpStNyCYMTADo4KgCwnDMquryaJ9eXL0FgRYUmb2hGep/3MMtTs8RWwsU0kdu9geNLw3KIhc71hqDst3jUO+J8AOySbkZdqTnGUzfab/Fpf3hGOxseG1zasO3nee2FRmouI3iS/834NS347BtQWvduP+IjnR0neFiP3Kg1svGKb1uW9CheP6rLzOz10KKQg7+hyXKU4Nmc+3JUMFCnO3uPfHmMZEiCOoIHWCeNWDKMUceR1c3M6If7CLRhyRrMF3qLCYy/O5ozxgygDLom9V8D6ADFpPPHMBmNq58G6hAQiSyhe0bi6rsf33/e/fb7b6y/r7I6BI6jZC6z0B0tHeU7LW/W0k90VFC8KkNBsroyn0f3msv6kE+45FHP1Ix1CBnP0iih2yGjIoK25JiIMX7+/AWBdbGuALnlWGF7pldmSwmINLgPOnpkqZKYVIDQBMk/Z7kY6yVhT0WddPd+8vICLH9kP0A7fRxhDzBOte5HvWrOrrYdUHZLApLSQZ5f2cw79v33r7+jgTiD7bgObqQePCN0ROxz8INochs0JxuX50kScTrLJIcVTo3PqRcwwCzmQocUNMFBtXVABB0fI3/ClQbHTa+vd8Aa/vjjj7uvX34DrcW5/fr1K8o/BRAb9gt1F54TlCibbJqg3Uc0WGem0gDi5znk+5EdEyW+ZB99/xaVI6JfBUtOocxZXOfeDbKlDRjXvKq3RLwvMAqOjcGY8Zx4njP0KPFL5zA+IqlAvbaVxabjjYApAW+VMJIN7Iwq6/0uGYZSws3pYidNvCfoO+4L/jj32vD6xnU8Xy9Dc/PVfiIBJYahcQZ+BEeInGPOFIhrhzI/cnzGdL7/+CEbWvZQd1IftCnyJZY2dKnncG5Fb514ZmQUVWZeCd+u37N0WDjBKKBpL7M8VXwWPPfTZ2ZpYfzRK+HlBbxi9+OzH8/BtbEXKpW31btjf9VnqTsX3A8FPEuOCp6paLZOfhfYWWRbfPtO+gVltUC2t+wi85jtRGRnJd+a5X7TieksUmlmqc12KppPk3aKH9gBbnrHWF6Yzeo+TuRrtFdA+2mMKONIAx+4zGALkkeJSlMBG3XZuFuyRTTQR2p8abaLS7we9Kc3Gn/jrVgT7m/8OPuVdMjydlBZu1PI+MKFzcVMZWsAACAASURBVPuRUXFgGB8f/11XQIfoRkfF//Pv37olBUXZAp+18NiQyN54nqJeBqmUnFXdoWEWyjhTC1mqCLVALZyzbJRLJBF9RLSKDq+hROPnFOP1A8U3U/zo1CBzZ4Mk1jRUOixAfIHKLVvDdSWDJyA9Sw2AQ3nKZlmqdfj4qMgeNS4NRYSed86tFKaWmgkwm1KFzGgDSpg5wfhMtTgjBTBHe+57+t+BFAdGi/qiVo/2wM7yGAEZiGIOGnhiFBPSgpWCCmOrRfFI88iUdSvMjHJiHguFnA0UGm2fw3DQ/B11NgBmMWQpkvGMqElrQyqBkSY/FlrsU/bqugeGInSsmFiv3C6rnRZuXDkYsw0ks1DPf9UVJBShePA2+G4q/aUBULTxx0pJCWJ8utCTvzeobgXcEXa7uTlzZf5uVFbjWwEuMZdNXQiYTViXMsY8Sk+kFF2+bVYOOihVJ8HTrMg2Gsgej1QULUc3XBCp8hrKJuvb8m+u7AT95PSbrqD5KHMD6ajthHIQ02fjU+kkbBEwN4KztRd8HqLnEhApgj+UJMc9PcLa2Uy9BBeXsACWU6RszGE8V7yHUZ81/x2+02lqBnpmWkjDWSTE8fdsPa53gbSSWQdgdHuOpw9rJSdq2Oukg/NymBsz4svAVKTMLtrG817P1148pC+1OfV20fNJt6kK1CRq7b13K+/AnvZzfQz71TN00k2WppGNhCvAK8CtxiPKwMowTC2rhZZ5Sclu08BsEPncHwHFLUH09VgvMIjazwpBh+0sC6HWo2CUDTMq0Lrzunyao7tstDQ6LDNsfTd2001ZW8bNCJCM88NTpC8yUKH+Tt7rTCZHf4J1UqcIkIx/tjIOjYSTXbXX5sgP54tsrvi8OexocNYDoRa1MpF977lFnBQNdd4X4ANKNbgZsyLBO4g9ZDlk0EpuakXj2cnR+oNQVetyojkq+rwn3aQD9cnSDusEMCv0J/SCelbNbcq2k6FNASINQeCM64bvjkb1dis50ekpz7vmkYk1tzBeXYOa3qa9CTqNeTjil01Q5ZJPPrin2f761TZptEPiT56O83Xi++08i4qW6HIDDmELPL+wlFiK136OdX7Mas2JkSOza0nmd5N6hzGaPwVAaKdbZbyWLqYwiSozA7o1OELw5sDRDkuiwDXJ/2SHLbgH5V5D4X0gMBPAaYDRBrZiNujhIUcMgSqW6w0AEc90eTmfYenC5Metzr2A3ghOC7DbtgbfNTUwbnthexQrJb7OTEeC5Z0cAGaqXBwbZ7O0UZbPAqgZ/T8EDKvfwrGE2o5BNrhtI41kP5OvgV8gs5slssgLOG6WJnKD50knnWjZPNPytPcxIkGSKL0a0ZOjiFB9NGLualod19q5gSn6f9zAFuMjCBz/odeHbMxoVB50/I9//H73PcrLKMPHmRekFWbUBEgetGIbvs/X5cAAIsspEWuDjI4ArIUVsN8I7dPMWlKgS/YveHoCr8U4I4hSJaK6/uaAMmAIwgSIKTDrNd4TdBELSbyAgaIONowxoWSVSjA5UyOcgAhYVLQ/eZScnVhb7kruSIucr32VqSSeb7qO+fyQs2akAcDGad9DnnReAW9+k9EXNfQt02adrPdFo5juNFo8Ls/fNOfMZrAcES0BxFcPG/Y4VW9ElW8FlqDP5vOFwB7xUYDr4kXp+J9sN/TPUWBerJHPXuxhvCN5izJcYoanIAJnVIS98PkLHWDOIOTyjH2AjiK24TIxF/CJGItKQlpfcgAAgrGQLfOMvi1wjP/cO2ZuEes8ByzFR2eL73LJvFHu7HR1jq36NXXaPus2yWj6aRgMKuqAHBt/b9Zfo7+t/SD+57JWcEpHWbVwkGmizHSkHEF5UQcQtz4YPLKjkjHbg2+tM++3HtcCrz8yKt5auo/v//UrYCvMoB0F2qlHxeyooJjonr2m0E8N0poJdkhx472obJmpkTxQboRLVUuKvJjE0ytBfx9ce1YtDKxK24EBhUBRH6WYMpLJDdSCYYQDI7zijjYPm9JKCJkWxxsKULw/lCUqwdWkl9FRrh9YtVvjOjbNUQ3Y0EweXA5BzY0HZflkDnAMO/zDYGsILjo7ztYUWFimPnM/HcGfO9pecj0amTcphKd6wjbyFPWRYIkiQno6LPe+mschoiSUv1A6JTTYCF3NvBsua7YcY13SBb0mPbqgZKMW1f8Y/HK6KCOkEgi8MlRnR4U2q0dgprGT75cwaYCe3BWNXQgoS6987UiJo5G7AARJBXW3g1WqaohSPIBrV8b8+Gav37n4Qwf2qDqQSOKs+2dSSbef94NwpFErjnI8mf64NW0d7QhTNJ15UpbxGibpknMT0JTAvM+pv++jm++xk3B1VDQNblri/X6a5+HirugcwGQaZTT6u8ECYu8A2Z9yVJgPjanIR8CjAQbbWU702RW4WUFV0RPusx9mi21cUW3YjmeeI5Z3jyj6XUfvbDc7JlgCoORA3ruhy2FuU9ZaH0evT9tB2OGaEVlZgJato7w9YKnQugVTxLPE19Jd1elKm5LGfJKtHBXHa+MLfsk5JjxCQFEOu1HXf0uKXe0mv5tsh+JJ7fwMBsXJUTG/ykb85NzY8cBhFphnlwXNqDpAipQXNPJzrBe6gpY3SwhxwSew1plMclRwsTTJfu4OS7w/dW/vx61XLPP1RmoqJCSxAAHiiMhtwROmKb+zSzc8Dvf3B4pe8l1r82zI6B2Nn/YDQYQqC6EAEWJSe10vPg39iaVuKgI5S8FNCygVLRsHm0YGp+Fm0U22pZNP4+ns922cf3xDd5IVc81rXCYjdLQAAQBeH/r63EovI6+s9U4n3YWjZ9yLWodGBg0EsUO23thBm914DSId55ImXn93BREwcpVALEoSidYciJLZuSgv6wxFZxX+gqPCDqME8Jr+ox4Lphs3q401pH1G2wTOKJUHcuNu224DOC4bIV2iOpPpgMTxXIEnfK9mvz6Qg/rkZu6ud48IfEVt9wvTscdSRm6ebHDctg1BcwdxiO8czDV8vJGvx4ARZFm0csoqlexo+Mi4YLZHlMoNsJONqWeZ7+GM4DTHGuOPfYD+qB6PCEiZzM5is1GKiQB7nNEfAP4/ITHm5Y4NyZPl6cUMmmHZJEcSu+yQI4+/fvmKyPvM6gj7+1NkToVtTp22O+ckxeEchPNB5cECSPz9H78jAwJjjvmpCXbcg/4YqmSADBDtPcmpnALxHQL2Wg+D+ZzifImHu49KB1yDrl22yjYv+HfL6ovv6eBg9jCzq2R3a0yIaG+9Dr1vIKdGs3ZIuOTRDKBXEBvPLcfGoFLOo7INy+ZUJlgrK1xZ/yvnStLXuPx3ZDUC2DcIn/4sXrG7r2cKWSyDvCa7IujDDqi0f1sljaEhcxtynJu0l1xabedcEL9zJg77sNAh1vfAWAZoxtkWLaAhTybKIxOH6NkHuQ4SwqlunZTVNpe8xA6uBpbHWYhzAjAdGSCRPUKnDpx4D58wF/SR2PCuQxeH5E3g7XIGoL9Oc7JgzsLWZmdBqQDlqOjci/zywEwPQrPzS7+vB7bs5fDuHXRSw8mFDCqViY+gBOglzCBCQKgcQ84o45zPjqaTo2KHYcxnvF/z0Uz7qDl9fPH3WYHUYmWsvuGo+Of3HLpgASg0IawYscCfAPnjx+mXZpY07i4AAuENZeg4+kXsV175Pgg4EvRIg/IYixVioUF+K0pRQTFkCj/SwCUsnIoYz7fzwQo8GYeNedYBNkP7/OXr3fOTG41Xk1JHcmA+TdhE3U1EnmXTcDPZqmOqcJRm8I5Uc8I8nNZtj60F8rFhnRQbRiHRSQQF+pGCAz83OClSCVDETmSXhHKXjLfzcQRbRAQSlbTK/mAZEo8ZSokMBioDMbaICFQzM6yj6mhqfd1Y2GSWgsr1SlVfFgq1x7RDgLq0a/V7meUSERi86QQK9N2C6tgyX15iLIs03cCBouHnbbOm8zmi8Tr9qL4i1nYCrahbq+6llAKDuY4Cmx93dlQcxhUNBd/F+MQMuskkOuxAZvGCaUT9gMyAn/nFNJ5Z+DPasfrebB1+IjSe5XHuplkeof7d6XceNT5yclTslK1L4HOMNh8iQfYpOojqQjkwlI54zqir+fKcizPxNvt6zqggFczr0YpRnKnkBj40OyrGPZVDezrvpzr9e4qlYSrGuB/rVJ4Dw4YVOzlIHsw1R6XUUVazo6Xzm0tHRZufSzzBgM31W0/iAMRMtPaWnr81QgY5P9K72mwyrjYtqbaUeGHRP2TEAOAW8+zATV1zm6PCBmbyk1sdCV0BOVBrN4Rz3954/iyGxjM7vmgnuuiVael3E2i2GyqNdoEL9OoMte5Xvt+dDo6QbPQkkoZhKRCGDlOdezujrgInNoKiY2ezIfw+udIcM12G11FUtofOi5yAjPxVr7QoceK0+4pYGJYq9Y9VECfvGEQUFLBJdvqCBGymhzWnhGsa7xydXUYiW1W1oR2ckpG4OwIh+pbOiogYdTDJ7vIxIlTBES0zhbzfd1bvuXepBrPcFk0huEbBGwa0Cdi1uvrazyu97aipaL2TX8xl9XZy8JJ57ih3ZYjX/FfNn99awPYqA/5hO8X6MOo7wOKySRxxHoAy5RdC3rOECmXghQ66HQ/HupNrvhxgd9Thlh3gErVxat2HIOyqWBPSYYBabGzt7O3k/nZUyMbBFFRizXMCEBV24GOBQhbvHbAfWSkOhfQY2ZIqI4MPG0jojJdYP/RtQANdBjs5KxtZ/Cq3E79HBP6XKN2yoyc8v+SfLzk6KnweolwRsv/ZZyTYsx0lduaHVWL7b+eomM+M/3Y5JjoCGOgCfRj6TfvBnyz5FQ6FKE8T6/Ht2zeW4n24u3u+e2ZlVt1qrR4Nwl2eS+WfmBnCHhTkK1FeiX0z2fSaZbucAYZSV/cBrkfEfPQbYFZEb2Abem+UY/r69be07ZzBnWcCsmAs+8ySay1TUEwuQErfR9IQ3agfBNZbnpmstT8EOLGMm7OGHBSA+QW4q0wNZpgxEp7qE1cunk+cgufFYzlF6Xt8dgbBSSjHXDi1wqkUFQqYvcT3ESuITDZG1WdkPApd0Man7iuZqnNZZZlHMkngXx+bitDxRI4gz8/2/UBpSTx0oMSPy4T7+LAJNXu42PmFeTYnA23gkmF7FltR9sxGYNCnnWgl6kSjcu7EixDkqj4foYMFjcdeBZ4GAFt9UVy2Kt/vybqfUe4FcZtkES1Ugna/VAzFnWFLRCseN6uTtODO+zuVyos9JKWirNU9Mazs6/PC0ngDrtIW7OSoiK1iplDZhQTo6eXsn/v3k+wm32DmMp9BPnJyMu33c3Xsmrec+N9Rl1BGRQV+inerRB4yKyQLQKPgmRUIZwyGzqiquOLxDPxkY1vchE19ZFScyODj87/PCojjGXCSEDhmVMhRUeopEZg4UI4KcVQFD1al9xe4dVZuwWBkDA76jco68bNi+NJ7yJhdd1Fpko58XqKyJXwogJni5/4XaICc3nYySo67Ra1NjayDOYfCRaZgZsuRhiPEyrW9o/j8SfUZu1ffEd5Z6sjlZmrOXhNMoRkJSzTfUC7JTZg41/nH9rkblfl7CJYG8A67tgNcJGgMsn398iXrUA5Rfnb2oIQCM2i6UjRnx1RkUzlS4KhQSbDovUGQXXtHLl7NgqUUuUFgNlIUoLOWIhgBFS8zHUAV7Twbv9uF1dZ1R4WppBpsZ8uE3NE0g7Q5c+mdXZTXeF7e56jgkim1cVJu9hkEK00WbRalDAb2Ox0VVFYblTeas9KVc9Z3s1IoUiijZyRinms9ZDaeCTQye8sGnVPK11NUzozZoHXaZ90z878ysnjNIaNCYE+CBh53jyQaBlaOillh6TxxnotT1F3LF+BF421cU83hFx0Vtda1FkdHxQHc3UmRvocGinuDUx6ntaTKux0VW0+gzsQGROjA3BBa3sojDGsKvrvf2C2orsXI09L+hizPqkMzCDb+bdrdK7jOsllXnqeoIb0iqjoL4z1I7toIonQqCQSDzMR1L60UYR5Y7GauR+eewWtMsz24QKBNnW3qLiejfSsw5zO2uagb2v33HSzZb8dcbV1JDxlWdUC29yBnljbxg5vRvptPGfrVDPgY1DBBk70MjMsCuNROnrsGshtMsQPjtL47YJZrwzv+rKNCXHbhY6Y2gysVVR79AtjAkPoNG3wORDwdC7OImX2dtoPgEoGz/Jkv7hkqub9cl74Xp0aNYQQzy7dKZ6Jxc0ZRz6+vGtAmS+ieume3f8hYVi8B3lPls0Y+uE7z7fO2vyKluMFN6wOIDGX/hORpf5GjYu5bcQLfOy+d5RNno9JN2sOR977FMQTE7A7MtFSjjeCmsOx9FqB4gOi0+9RUWtG6KC3jfg90LXPU+c6NJL4o63IC1NMGUPAS7DNE3RuMrd4J8X4GkLF2PAFYRunDWaWDmcCWnN4xZNfGh3NDZe+qHKXLvfVsT893OhsOMmv2pBZmjfjG0VYDWZQRom1cc2B2k3vGxbxP4Br5dWOGGtZVRgXK/gCkZ+ZD2kvBz2IdP4XzkWV6Wb1gI8uHPR/XIoBG4wCmDZz9JbQ66u279F9kbpRTA3wCNsJE8yr9hCbF6r/o5tokxYYZqJehHco9kyF7dET5JwG71WCZYGa8OwLsiCUEwB9ZdKysEA4BN1r3Pse/BsDtqAj5gMbzT9E34xm9Xb5/Yx8KB30lAA5Qm5knbuBNJ4o3mfoJzyDxCJdGc1Nng8PhecozGQ5FRG+L/yJ4sDkZkTE0Ap8zZ/Uau4qE99X4DvogaE6Wl9HXAzobouOj0kFlmGR4nIH/q5JGcuKkiDOI3RwVxlMoX4pm8jfxIMzTDi1nugor6nuWpblM51aap0ynVQLR+YqS1700Yr+wKQFx3R/fvt0FPhI0EU3v/ROOivjBGQUuMukDuSCiEGTDsZeQ3x3nGA5oY1YtMMQmRdf6wdHVB8PPSRYjp0t8bsdqTCX41M+nKLcWgW3EvpxxdCoJbb1wXj/r38ww4FnueNBsi+xtE7KssgXKRj1ev27k8kmnre5snOny+A4srii/ObwYUB1OPvJ9rxn4zZcob7dmbX44Km7YsI9L/v+6Au9zVPzHkFHRlFYtT8GKBIN4RVN6wCl3EFNb3/Y1GYCAPKfh4f4STGjO5pRgAxeDrqP7B8FRYV2oGadGPKwHqRI/NnYQUU1DBxEYroOHxj5WYpiCR6brZl18TjZiimbhqnUX77ASRRkr40CNvOxRLkY5rhl1Y32WQICFF40PptK11T8Cfm5yRObIHhOrVz6Xr6VvzqeiM/Zu9FuYOnKHYQvsvUCjnyndcxQCoq+U3WJlCKULUMSTjpRovP7yynThJK3YI80XNNSa5OE+kVBScAfBB1KsdQ/FwY2fMmpQRL7LLlgM1LZniBDOfitrXJp6PSedL70dZKicBOTL9owp9TfWdIncjEkrM4WaiwJ31uyLtzhhB4ZFkckdrszukTy5QSTtsUQQTosBCX49/bTz7u9k0PjCVNSI+q+podTwMzKDvzJ1c6/gV6Ttuj7zrOeSHxqvziqdJ4LUc/wGxTSm7ixoPTvGd49A2kCPh4yKuB8KlDKrnFVVDTu9lYqkLqt5eDVnPNbk7/xAIZrD1h3Y04rXywCZHWh7RxONc4Ns3oke4Q0SOr583TtPzbQ5ipWTbFtpmHRM4zwnWR6FIfuh41AwJjjoenUXiQLiJvEwkeUKRFim9i0tmuG7ujyuB3qN+lrp+kVA6HM3gNfLmpTnUmSmIaqV60S05+fcr3pUlKPdctDnGEo/yLMypt6GBHecb7/fs6Mi9/rEPM1rNru087Lm/k+yn7c7o8JpdclN9m8/lam6yHjwgzqQTyOTdbStCw1OlxaB7BIWK+/mkw+nLsf/LkfFbotcPmhyuCaPSvnszFtFXzawDo2EG9gzOwnpqGiUPaprw/HNc2V5BGWmHW+BxoxMNXcNcKIcDm9HfpJnBEjnKFODPVWnfSSRGJcbV2YQj8CLMym771o5KVbZzruTL//a4StQU8scQA9BUwLSzqZg2Rjuxy1OdoxtQ5xcfz3HBk4DSHZrkuCJF8F0gCjl3u+hnE3Fa8fTcIM/YsdBxLvrK+9lzNKlkwB4fuJ4Yo064GT7yN8lPzu03WFQ7m5TS/cZdVc3EWeTW0Y5B6DsqHFGyBtICxA1gDGA62rmDUA3yg+Jg/S3u0Ex+oA8MzsPwJOuhTmiwLoAfEv9SwthOI+2czJLTBHADAoo3Y16RpQKekL5oJBrAfI5kyIaXiN7RHzTGf4IDlFpn5mmSj6PjO3sAHqk/Qq7h/dw7rQRo4wLMw3u755+svzxTs7He4c9awpGRlKn05/nLBun67Dr7Zn15OwaXAsng7J4c2qIN2aGH8DYCFArex/ZAjrvlrkGORFc9Bglm55QosYZQA6EtMoE58Ere1Ki54XtUJ1zNiNmA+0Cg6vRvO1L28wAbwXgx+9ff/uNPR3U+8A0nDY2gHTaOjF2n0fsh7JCerAeiZZ2Gfgz5hnZHJRHzDhQGSgTDzIfeH76GYq5Rgmi3Q/PPPcxHFk4j2r6DJzgIcoABW2Rz5L+XPZJOnfrb2x2gDVMZ8DmzSkn2wnujojWX2MfBFKyE+dK9r8BcdvuDj6jzsKzYN066dz9OS6dOj2IlU4lZ3v02VnuxL+RsRNZbF47Av/RO4XlCr334G3hJD4wfjpbKwOAzcHv7+5RNoq0YF3x+AzJc5ghLh9JBp/ZJvFr9GcJPoKzHhUlwoeiayIbL4ju999+x3k70tNJaZAukGFJOd/JCXUlAHvmxJS5c7LvTmqH6Sp4Bh0sKm3WaC/1rQsHbqwJSoOJv0rcpFPlETpkYSzhqPj0JdZ5zSSZ989z2u1rPxcLDU5BBB+lny6I8uOrv8sK6KjemFFhR8XokAgPaCiJVLwdpQCmN00Tuo0iKi5XYLixK7erFfvwmUqdG/+4f0Qxp3kcVIqhsKlXBRRVgfQExJna71RApu+y3wQ9oaNaiGgPpSy/vj7Dm21mYUcFVxrmfApGR+dB8RAQiogWgE1vZFR0668xH9e7Y0oelTyozicwLiPH5VlyevuEg8mC0Sz2u+c1cB1DpGZHVJSVAIyJioqN/Pg9UkpDYXDkG4dqVZJCgk6MiCh5vfsUgHEYHKrxl03srORkr4oq0xIN87iPjFR4zaZxI9adwsuOKlExM2c+s1G4vP9Winer4Xc5gtugQBo3NoWnc0InRVfS5NBZXtKBksloGXEO3WkwvXt08iv8kinOmnuPplnnuAfpKhrCd3gu++s7Qc3R7hDCjW79hK5ImlKgW43T4V9KAa3xd8IuQ3QW+FTomZ5bYMOJa/GZ1qM6ODFHJ/Mc9rUYHRd0U5Sx28+d5+pneGns4BtH194x6Pzn0gtW4v2coQFgo9O3wB4DAOPeeY38fv7dbNLT4tbnA5+r+e14mw0y0KOAj+b31n5xpOdzfIBMi0lMYz7R+N5RIU9+c8p531vzb8Mpfmd66fr8GZFno8T800CgjkGj0aKv0v1z1/IgzY6K0watEfgXZ/31/u4lrCux937uch+VUZFRauhN1CIAG28eQRXRlLO34p5eNzgMLpQLid5QBlTHusdvE2G/Yj/Pbih0g+JkGHV+0Z+4A4Zyj1ukXIHXOlHdsN/xxDYF6EtiXuNYT6MVW22OdtRVVoSyMyrxLO0TgSazY5WBunj81o/eGfx7Nmm3RZKxBmMX3q9G2wY6ABhhPgTrmPVJpwwjkDnV7qxgDW4vgely9YlzKl6csWyXl8gBEjlOG8zdUSGD2QDdDmiPQQYg4obNBCZCfya4cjzfOCvUIWMMqLV/uL70nOZwbM6wDDyyrla+l/fs6uCksL4U62Rwm00quYK9Hrp1jBNwwxN0sRZ2Ijkzw+UpDvTcz7YfG893lLQBNNoAbf8XAKQyU961UI2+zBYIOEZkLMGy1It9XpE5LLsBPQF9ZmdHw37SxAbXiG07M8VumtNNARJwJLA+OWmeID+ixyewkvbSI4DWpDkcuDAxu+6jsCCA4ZGloehy/c2yLwwwi+cE6Bs2aupCh8A6nwXXlLfj0hHcDkTC/gdQ9RBliX6kLRS2BErEKNvHdiKb7e5SDhunwLJPOv+FY9lZMghGUoR5rGs0wkWpIABqsedBE478n5/fIpans5+gb8tODFJ+eiYIXnyR9m984uwCBv/xs6cXNqAeeKkatqNxb/TQUCmjLwB3oz9C8WSPg6VzPuM5BIW/pgOdZYxiS9xTgfw8MQGBh1/cnPiO+/bla5TiUlNlOcVcsjhGT2cTyyw5Uj9e5NJPlouUFes5gq2lklXIEHp8ZJS6miybj/neeK6rBMSc7OhgEABpJe3UTxVgFV+51F/qKdN+xnywtm2srLjAAMtw3IBvKdMDzrdwMtlRIgY14MoEISrw6AJ07rx51g/Jr9hQnHyk7Blfm6qyxuMqDVgzrT16RDw+wkHlyHbI9pZt6OcDEzo6C0R/aq7uklKnksmWReGo+PbtDzgs4gz88V9/3N0/0kFrp1bMFWt7dJSEzk+Mx2XDsC/3KuF9o2c7MAc7SNBzAlhWlHUKJ8kLSz0Ja/G+o/STmtZjD8B4z5Jpb6OOcmLI0G3766diD2i6rD9TRoUdCVcYxmm4Dtzwa6wn0W5oPVOdtXNaZ+hMPI+kH64T7RoGTzyFg+qOvUpCRjyFTrlxUs/013X1W/SBbiMPZ+qj9NMty/dxzb92BXRUb3RU/Oc/f2QEBvtQOJU8jB0qXQECk7mqUbRqjeKAq5wLBEIzZAdFJupUpkCZFPdJ92U0jQ0ScTAxgTjsEUnx8webIAbTQcRKCAM1S3N9vR75l/uRwrsixGCwhmJlDpf9HQy6segflMBQpH5S6Q5hSEUoWd/gONiCNVAq7cAY0/tYt1VR+a0B3edP9sx7RZUtoXTuRb3dIVlWLKmlLOQZuZsdxAAAIABJREFUY/VeQgGwQShhRdCCRkRwaES2vbZIIpfSCUURYJUMfZRuclT/QRI5Q8SZFk1iIcKkycoXPWIok+qajOo5kQ4BjYH6v5VpTd1DyT3n53ME5fBZX+g8W9z+fh8EoJVBOGw+QSmmYGyle4KmIktGJRXs4LIx7mApOMGUiUCZXmAcg5J83qf11Z9WUDLS6gK8mLWFWXCWYKx3ZURjpOCjREQ4Oc8RI+tZ7MHnBGbzvROlDjM0sJkf6heXu2pNw6y8u2RONywWHwM02TY/1ZKsLCpcsGHxfXSjo0L6C5XwfufBaXN6A43SVYnvCgsJeTTq3y2P2v19eZf3LM6z+YxfA6MD7xLfstFxVMJUQ9UR3FWIsDluEcnXavQPLxJvUvQs39OdCP13OpeXeV8sKPnN2H8B+zktxbhF53UyiazjFM/qW30kHIIW48+OHw/Emc6WLssydT33XsCh8yx3tDNNHo7bY2srjWsGbrLIdTk6B+AIazzOCTrB5qzO+1n8YXT+zzQ4AJReKvMh92ywAXwCfefzecPhPNlMNCb102TckZqaQ6zfR2Px7bM6UscYIQZZLf1lN6UEGrwf+KAiz8j3WYrJIAIMaEV3wugDEEkHCeaOHlHlrD+Ve7sytjmKNved0Sy5m5zDoqY5lrbLh+sk82eefJLDKouSYA30Ka7oDJAnWLl71gmIMbAkxtJVIZaXKqWILHmMjI/bHInsvgK7/Wbk51hX2s8enT3XYP2V84GyTnxQv3gprCtx4bQNKM8QADllA8u5sLTQ/GOdDuA2GsuyZEf8HY4h/+21cAPafF/bLwdEETiXk0D0C4cSAqwYAOTgLLIJXktQi5M4rYd5nde86LrsQS8F/lX2B/T90DFlA7inBUqHuWY/QO+o9U7Q36UvSRthH1Yvw76OVd6G4FU6NVTGL4DFAPV83qGjykkRn7m0ToB8EcH++nAP0D16FoQACRuQQFMFqBk8ijONnoHZ46TZIRtHxZa3t+ArB3jYabbUmNfEPZfKWqK96yyBkc5IvOi5kI527jv5G7NO4JgXaB704GyHXk4FgPoL6+B7rOSVjPB15v8AqKNUVdF+yUED/QUCe12jR4UdXmP2Xe89KX7l8zkBlJH9bYvs2/cfCDQIuvr5/cfd19++3kVZXIK7EfX/wrJOqvvOLJJmI9gZIOdQ6kugadpXdNrRcRb/wkHWg8lcUaGX+/H57XakSpLFWrO/Ec9n0GzMYejzgzLI0kFV9ijuMegNW1r0tRM55mrZ/6WJqDibKNujrJTuLIh3OiuiZ3OgaoHeGY9yNlNc6zJY8b0dM9R94O6aWCOdGyhxFo4jNyLX2e0OHfJCDtzvYYARMwMM2FvEVVDjlBHf5FuWeXbFBu07aLeNNHUanR2sdfSKeH6++/2337BnCcZT+cDdFtnuKeEG2XHuI8BtpzVTRqjahebrrA9nebG/CkuNwXEpxx6avctWpaMqMJZqXs4lhNchs2uMMZg2IB+QQaTG1wGS2znTaB3S3Y6BWeDFAy7SWnfNtK80xs7vrKfYUWy92jxtDqbLoV294KCvXslHyz87xOwo77wfY7soc8gzMQ4sdShUtlh9Ls/v1a1ne2nS71I31H66zGHO48NRsVD3xwd/uxUoxZRpzfzv1KPiP/8ZnnQK3IoE+ZwNzQjUUDEIpSa8hcEQA6gvpYEKRT9APq4Zba5aumTKNEjBxCUHk0FAQZNJY0yiOSqCsSOdE2mbIXzcWI8MpCvqy9Z0q0wBoMgYgPJd0WUcuyNmiYRHdIFr+q0R5vEmrpMVjM4wtwAv6raGAGeDa2cXeK1peFCJhREEKcoxwYiy/dsn2a20ibn5nm2UXU+9hPIl/ULKMowpl3NSxgoEOSJZuf7pMcZAZdK73NRFsz1Ewzw83H2O1EMZULWKf95RQe2D+5k/nQ5SO/kFR0V3bug1KYS1/mF8xk9EA4UTws0OIyU/HBVUOhQBrDUu2uFAafw4CZdqLfdIhisE2+gAxB4I2DEIxPq5bzkRap06OeUyljrHNOVU7hkF4iiidN6c+OOUdUJepdPTFdNdsEUvk9adcAIrwQkM6EsLxjpPdVJ9nhYwU4as+Vksbzkmyw8w71MnsAEM3YGyDTQseq8n7HU0ZxNJqSaz4E0Jtrhfgz9/HwDJ4+Bn1KkB1ZH5LIOsN8xq/NvvLpZZhoLXzv924JJ0qNIB+EPCojkMOy3NQFZkx6XjMu+pbACet5loN+ZJLsU6Z9ZxrhNQj2sg4LCMF+skK/Zf5ajYhjphuNVMOf5Cy8Im/+Kz5Egno2IJ2OprOfcLMCg/gvMWhBiSz60YydvUV/zGPLbL6hn/dRTc4rjq/Er61tG5dQKoT3wS89p/WXyrghguLidhz1mxrcbz1RDm7xyxfalvraxiiJqfdnvsySB+47PsDM4OKrPHBBuFj7rnNNobCGE1Pmt0HoPIPh/uVTcQtnANkHBX1BpPvtFRQQCmdHqLXztopKquW3dVvigVPOm8jemlWHJ/MJUscPCQAVSKnPPCJmBoGSXHiR0IpBuJrkv29/bm7XSNec1gv0yR7Y6Y3+oqkg09uh76TvQDiX5q6I3g+u1qlrmTjbK9Qv9jRC7nk0C0HBUsB9KiqHmV6JoNTh0lvDunO/2Ja9DWrwUWWO9Mh0yWOBppwkFLyFIQ0BlR4TH+Kp2zkY+mP5C/GqIr6h3lg6TDIYsJEb/PCOoJ/TGBVmQL0dZzA25nCwXpudcWQWhmaJhH0/RQFoX0BNurGYgyLI3rjo86D2SbgMUEM6UH9YyQvifQg6V/sq6/9lFnqq7tB4A2SjoE8F7ya0Tjay3s/LETJ+YbtfHDrkBQkhvvxlqEs0ZSmPzRTjLtifR3LE/jRwYO4x7buix/EwuWBjtIi2tQNdl7sEAub4LeJEf2tGDZ3bAfXT4LjbX1fx6OHdSOAOf6dN7BbDA0Kg47OiOk2d8kzmpWIXAAS5Zn07NaH8vMZKRC0baKfNxZFAgwky1sENrBM3RYPBU+oswFV4mQ1kGHi9bewPZ4tkk7DAYN5wIzZeKeKCfTI/xl5mQTaThPYk1MOz9/ZonAIWrejtCWGRHPQuN7OBSmPpipYzWMwP1M5QzoOkapfi2wwSW/dX3X802Lxj9qPYp5ufzRUAZKwZXOsOiN0DN74DPXDMGActb4+bRtzMcii4ZnCTTUcIyTjlT6iQJ2daGbujMglvqKx0hnT2T3h/Yc633hqJCDnXZYyc341XzI2YfxGRzpysoh/CEA/ihO/zpHBXi5S6U9PTPLy/1tG85o+dEzk4b1vRL9B5vixJMtczuv6xgdZSWloWXpTodfZGrDJyBfNo6KU9PxEy3NzpbZDvYcyrHM7Oe0Tz4cFael/fj877MCZdTc4qj4j3//jsMJz66b/kTkEQScPQY9goHefAt/Ks8C0fGEBqLp0LvfhAUGFNEo8xOPt8Ne3JeHlNE3YBxSOOmJV6QHooGU4h5RE4NSv1GaLTSGd/BDp31xPKrj2iPwIcAUWaAIM46fYyh+2aOoT2Mo8MVCK0UjDAWmMHNtx2bfhWvKWQEFPxdviCzrRvdghM1Ao9elE6+cIdn8R1FxZayTvrD+ELqkh7iefTRq7gY2exT4HJJAp1U0ZJO3v5UkgDH+RkaF34Z/9Zw+nQIX2p74VwtC/Z1rNVw67uWytu1ZaXw1xZ/CS6UlsicLUTynpkPIOFKUEnWA5+kQoNo8etOpS1vILjxIY7PhEf+ytuteA5hl/06BHEmlhCMjra2MXp3B4Qntj7GsBvWqcR06ttMVy6QBgBE1t6t60UnDwQOWSBI+0cZd/O5oKRr48/rx+ox+Mg/U7KCozEtisKhNql+y36Eqe0ZjrZViyUaQbUkbILXQRm9qPn05O1ny62EO04TqoOXla+PFZRQN2x7hoq2SODk8QR+sEyAnbu1b1uPuZxkypBteklWQM8VJxnOwuLFqOch0mkHb6aZejHGOpHxzloaV1h492Wmjn4nZtq7VPkUtn5pphzEskAtR6/5pDun2Ka4Wn+5nsZe8m8nfcxjpvF+13qFK49NZEkhIqZSgbrKODSC8CyLojoqR9kQjyho03/CK2Gj239yDcym2baDAeizGTw5G2e5Z4E6nnpobtkxudqbx49BaxH7yodM4t76WtvP6Nde9UO6B9VR0tPQPAUDWlbbhjm+u7XBKREXdUVtlrfo6DbrCXNpxkGqS50tpkNPAGPSjgTBjxCWElCEUoAbZjka0E7eXUYHOzCvUw80gyVNHJ2v/rjvvTzOwXmyAhE4V2gkEoBxQpDgqAJ17neEKeOCJr/NpGbxz7MWYDBZZz49XOlp7mYuGk7qS2DzsBeu7Li3UGlMPJ0l0jRr3qFM9HswYu20iR3tTpKvJezT/BYAfupUj6eeAFI6cQCfFUXegbb2cryztK1YlG4aDtQMifu8ZEW6ozpJKrTFo7O3zSZ9svZq0nlBJBP4jAlgZFPE+18uPrAk0So6yGYpcp+6LEdIB0WgJxVLkEIBNBBtK66LMEThcnDGUgSgrBZMMR5lOmue+BA8KQD1Kumyd0WljyoZtjtSVX3OQyGmRzRfrnKXnFNwX7+k9SPg3s0/gqPj6FcB4rBUi4KEWsWTzwz0Dk7ieQTvl2PVZ9yoU8OVMGfYZdFYb9u5eJeJa6TdnrrRYIz7STbZb1js/p5MTgUMvtMHDoUDAUr+7XA0cL/d3P3/8QAT+ZLLhb5RpVmQ9cAuVHAb9ii7itThHot8nNb3NQ4CYFwfpzSX++FaUbNIZjrWL9Q8nkfV+B2tG5P3z80820HVJo1ZiEOXBeuP2UySCy2mpv4wd4siaCIA7+pR0oFSBftYVYz/Rr0TgMNbAmYl6fzlC5IRRiWzyAvbaGH4iQwd2Pp21xgFQAi3Wt/VNyWdAzFBPrxJE6qWRcVXWxUenWTospFsAc0D1DJbrYaBCjRFnVVwCvDUcn8paiLmbln0O+tzqPPN5lhk+bzOAPN+Lcl3CpsiTx55F6AMBG5V0bqe38ZG0NzcZFXDQuuQ3B5cRVdY5Y0+YrUEZUBmSDmxc+V198tc5KqKZOHnSM5xrv//jNzh+Oq/3+gI/7H2m+hD3YkW8Zf/lpaNC56zjGjPGQZqducw8qL3VcnJUvO5F9gUOMz2/4ZYuv7j2DdV5jb3/cFRcEfrHd3+PFRCR31r66d+/42AGk3PGgNMEA/RDCmYoPYqmCc3i1Z3tVSYITF8ZFYujIo0pRrf0CAlEd9smaxFcBgKhOOmQdqdAfAamDsWLQHAHD61wzfuxVSwlkJAZ0Mo+lSFqLUt1X1XOBynAUC5TzRsV153h9UIhH89GKZmsOcm0VGdVZFooUlerlM4IsKxOntFAKYNliHTdghVN8DV3PemCyqoZuAULlWFGB9jJZYXe47xyVHisUOpeX9j3wrXlXWvcNKFg2RQfjY8XvNgcFaYZlxhZUELt2SSPbnJUwJDX2nYQtGf/NEdFOfTKEQbF8Y5l1Jgyqgjx5hW3EgiFJyJbZKitjgqbxuvGAnxV1pGp1LUyd7zqvY4KPovNpYJ/dJJfS83wjXXNCDAYxLCzh/RWoxyOk0CfAdbUBeBZ2ousse5IO33hlG3bpEvEgwxZ8gvyLddUXppvN/5Ucx5Bd7k5ldizB2SwNm1T9mrYGBUzKlndZOnrfJBKv+CoyOOSA20jxpfj3P4KR0Wn9+S0zTjpPoB0TDnCr59PK3ub2rCI7m2OikEthfzqJf64zjMdj6s8rcPkqDjJoSv9oacrd9o44HvDowjyzBQloArgzUyTwTgjgpIGZomEntEz73VBYp7fLl3cVIIxHZOoV1qKqxnZ1msL9znwHnNDmZrr1Mz6m+HrxeqOSXGrXMcC6KgnWB4OIkTGI1b0lo35kwrjHAleUeR7HnMVeX5lE26HuXNUzEz7DX5G/kvgLH25WkOUQPBeTzqJDds01rSXv+BuqRGm2lyR1aQo7bXKh+QNE7M+vXs8q47Y251HUxybZqb893q4CaicFgZj1tIcSeBH+AuHotG/gY4s+Wn6db1mlRk1aO/mvEf/mUp+Zva0z7oA7nJUcBaXNadvIMyj3jHtEWpHo+ce/4v7rPfvaNzBOfjOz+p0knoIv0wQs688alazbGxFlarBdcuS2LELO09741vbBut4uY7x4wjsXfQnKbrAPetKXaYxOljlbdSj0CBcXO8+gOncdU3WaVAuh+XyUgDMlZke9tOXz18AXqHx88PD3Y/vPyCnHEzjjIlcfJFtfB7+CEfPR1PrzFxwSVzVvY95cK/ZswDr/KajghMhwF/NhCOrNn5iXtvgE/MLg4h2+OnsriXGLL9iXNXYGTbf4+Pdf/3xh0ruBr3K4YDyMD1AruguSiAbAIe+qohqb0vPqHB4U9+y7qhwAB/3mIBrYM0v0URc++AAqN4ceD6uczlGLmyVsiK+QAcA6rxHGec7NnmOfXbfIALLY7lBygf2nIusBmRWoEcBHWBx5gK4jXLN8eNgIzhfNHFXMwDALDt3zpyM7WRptieMC9nxn1QyacAitBeuYDGU3+P4UV7JmVMwdpQ5s+XWBOWhS9j5JIerKLQsW9GcgfhYgyB2NqhXmWnxvbDZM3it9fGsyHxmplD/mzkNZRh7yTxx39RzI9Y7MhD6j2U7HVHaV+BJ4ahg0/eiz9KrUsfqcld4RDnOmG0U40aJNAXcxlMyi0kOqCAUl7iKfYjrT7zUGQFiAhf9JDhy0EuzSXCOhIc508L6t2kYzm7hbrCfM+CqoncHQF08mfxaG9OCWY3VWHfAMctSjt1RsdP3cfVfVvoJTu3EjNgrI8509rCRMzHWzVlUW335SvYflI+jo0IKUzyybCmWhiM/q5dZrq0yVus0ndVUDQ4ZFX+Vo8IyyTZxXzPz6bjmw1Gx37mPT/9WK/A+R8X//h/B4CnwnRr99ctvKPHE1OZHMhqVn3n8xKhKOB3QMDmOKdMEedh5bEvQ0NOHlF73P0CkAUFwOCqmaLN7RbBYShZARuUrFIqniLxQ3dg7RDZxE3Ye0p0gNGMyaIlUP9fW32VUvD5DiWIGARVWTHcAU8t1apCTrE0XvSgyRoqHhWkI60h7jqgY9+iwYsbnOCJWTXz0vIiWybmdwgkHRWMq3aKbJxtMilHF6edaqT58XO/USP/rtY/6opkRIEA/DT79PYN8T7HfaKgdtFZpsyHMLRqg0Jm6+pp3mG3qReF5uYVgWyz+OqBMO8dO+0w328gegq5ahKCjEVOIQBFk0+8kg1DuPqmBtzKDLHwsL51RBEM+zpZqcA7ZEC79RMofuBDGqaivofn5FIHSb3qvo4IN58uQibGa7ldgdDyfpJd6e0XLlSLmuc5Oin7O/QivtyPt9DZlPfmgMgrOvXR0smh0DgsxKs9O44ehocivXPHmqHAE1eDkTEC2IlV3QOe8g3sdjSBDGlI2rMCn+wTMg8dpzXNcbBDzg/6wdpHXCaPA530DNzR4QqrbQPIJU0ma2dnc/4ZDOYG7qgFvgw6yxU1M2xDNS8faTk4FSEoa6XKp0bsbfH1W57aMLrCa1lPIV78FZvcz9GccFXj/QlDj+GZKeX1hc1Yb73YkpnzPvadMie+DPkgWoj8/dOLXZr37nqbaB9zTN89R181R0a4ZpmcVaCktNR3z1sfGBmRFKo1nKPaqeF2tXWo8Q4+IG9DVi6N561fd8TBGcu9P9kBvDXD1ftz63tzWjPzLXJcdoeHyYUXaWc9zLWO/n43ck1ayz3K0AxlYBzs8NpPYOWiKNNvIOgjNaITbHBWHBaTUqefbeGcmxOHnVbq2+3c00NMZFAANBaTiSbvtPryD51M18NtZhf6xqkQcp9FsO/oVWHEMRtg4KgzSd73WU1vSzdrSnPSIopP8Db90MLhnWwS9oJ+dQF7vAAHSNeSR0cvVQ2WlBckYZ1oZQNJw5h12HwKSqst/0CHQnQVd149HBQibQApisvbpUsWfK9h2dlT8v+y9ecyu7XYXdO/h3fs7bSE9HUiJWP4waAXiUCsoSml7igYrdYA2isXYOGEE0tQBG+IQY0oaCVGKiBrQxCGYokAYFK2a2LRSlMTGAtGgpRjaChU7cM639373YNZvWGtd131d9/vu75zTnp7up+n53v0893AN61rDb011DtTrJR1xVVI27LmwA7Osr85B2G5oeqyefji3hkmn6jCdsu1UJBkxqIV2T/S4ewwAPgBEymwC7Y7QB4DdM41Fr0E3wS7iN5dHMn8GqKxm8j5j2POITnf5lQtHRY299zUgyAbdUc1md46K0mNLfnjdzyVAmgweGST1Gw3GJZkJrKoMbGsA60wUOhJYyhjAOsoP0ebkWe16rWT2FL3tfeJSl0MLtnroQtGjQqW88MxsGaW5nNhafD8r+nQsMZso+r+wxA4zHrivzhpI4L0B/HCAtnJN0bPyvQ99CG82YA3ZYaed5hK0QacF+/4FH0XAoBs0t2j3rmMm+KngSPNxjC3Lv5EnO9o/VegMGB1lAXXossfpVJqlAuVaPBcOgFjr6FWAhuMsB5fZxJYHBvOVdRDvCAcC+iTKoYfzBofgDf6b5ZD0fjt04qyeZcvYzw3rZLkx9UUiT6oMH5doRNks8WHKAM3bi3Z6TnFTU5JLZfW9MM16LV32yjhLOG3cE6dnwuaqaxzhRHVpc5QwinW4KKXoseCEoVSbKky0oKjBZnEZRGBgzAYaIuRXGRWt3C3phivB5udhh7MRu3UL0KKqC+BSCdtdcMEn0lHRSyrGWGM94+PsLO5TK9+7DKSalcaJsewcFRfhGf6p298px8Qe7cQHr14qacYSajymSTiLFrrgxo//1hkVnTeb1vt3PkfvHBUnIfTui0+9FUhrS+DodY+Kr/g8RgmQwbJXQzGVUoqcDfEISg8qUjMDI5WVsYxEGsUSRCFq3LwuUlSRxokzP5btwAGcYFeDjw+jeZrqTkbqJiMuwgBhDwcLgwSxJmY2A0P2Qsf3ocBAEaS0qQrjchS8fvOSjbyRSvmwSsG4iShWrQRINhbvjRhfMxIhXuGmWlCalEIOIyGbjquUTAMFS447atyAkFYsOaa4ZQMcMzJwjWFg9DZWTwCasifssEIDtgduRshmbzEpRkAx8wQ0pPf3bTDAmUBnM3qdUWHVx34vywv+dxQgg4nZ9i2n6QacA+ilU+sH6+L7ZFR4mz0UKwaIBpJCYFr0NY6qwJqoydujG9XdFf3TMGyGRApzRXUhu2jEgdxMuxug5kcGMOK/bkJvB2MCJhPzovLWjZlmSDUnYL4jeQUdljYSVmmJvse0dXI+pHLaotvPnpMccd9f8wzyLZ2vLAFVZW8QuSfDm2Skc1QV7vh8GbI2+pw2zyizUtStpNvRWk6ks0MwykvBlMmsLRnuDSAy3zurQrl6IAAroK7x2Wtf88rRIJ22WXMsyDm/0H2DE6LxC4AGGv8n21GxGnN3LhedT44KsYgOLPUlmctEE4hrB0ugVdHnItJouaC17qR/Zb80Jbzz1Qs2nE/v0UGWJwZvk3WdHrR+8hka1dne1ZnPjApSJQMRyoloyZMGUzgsZbHitzaMYURWT+xEGPGTutHf+6E4282oneqtc9FUBkw2zn1rw5a+QAOqeFVtNIGwFZhQ+gKN79K/ljR8ZUht6OoKaCe5U8cz6bsu+fw4GId+fw5zaY1tKbzOXUs1F3CO918YkHYodPJgsEqtK86IeDODUtjI2OBmf8YAfKScPw/9XuvXJuY1YoklUa8zgwfaTk1lY9TSeWc8FwCN6H5Yp34GwlGh8i3y+omay7DPNQhda8dIyNgWixF3O4Oz9FzT0Ao0SmdlL7mKMhdr2iGIWHwZI2mgSQLzd4Ine3rCNgxzn3WVPMXGaBgEpF4Q1nUYDbsh92FfdI1Ks7oUUnzrZyR/X5wt2CmI4o1mxwRm3QQTc1HZWa+/eQ0aRuNaZhpUudd5zD3TjOygOyrKacPJev6zs5MlhV7gGkSkR1Caeqmx3C2dJ+XYVYmRIETW+pMdxMUD2AmAlxkDBMSYlRDPiBIhvSRILzdVUevq5yZwN5wZjgi3ey3IKyP8ww6RjQKpoOyCFxFl//gmx0j7Qnyz+ft4dCg9quwZ19tlv9ABYiRAPMpBUZyp9EsT64bOnJlP+5VnE84iyVtm4QeNEJDs+qntdkTJ4310VNCmZQYRwHjpjTN/zhPsoDLzOb3bQR/U729R+skBSRHESH20Mk7TeZXHRTy0swr9HXuNcjyvWMon6O3Zi2c4Cy7T43dx3KIfPNuLyaoP6AGjslkG2v382CbYrA1ruFVvGPRZVLlh04mDxijzbX8VvuBG1AH0I2NBpYVMfyjTA2cC9xOUoOBMy4L4L0sAscTZ+tMyKpQJFdNm02XxcM/J9KYSX2jEHs2jX74kOK8zE+C9SyLF+F0yy+vNPidR6cIZ/9PImm3Ecr/lHKMdMkbve94u/QRHX9C3Srr5ftC+e3kgG8pOsHFtaIPR0e5sE1BFc8ybNyWViPfGfXbaeM+SLPv9yggIrCfWzvt9wkW0NHTiRZYGS3G5pwWym6QPVcDPKDPdt5LOcvecPDfT7sB+z3LmOspRkXgLAwbJxypADvyMgmHxebuMiiut0bqaM+kcPNB16LlXpoPvhoFdvWShZ251oa6XRiWBrN5SWJV1Ejgq5uzZ06DGgZlCV3YOzuu21PZ6gjOP7nRH2ia/LX2De/zOUbFho+++/lRcgTKU04B1KuLrl8ebiNp/dXu8fvn8eHX77Pjyz72FYhoH9cnNDRSxUKIJZlr55zwH8GYCteqgk2mimZEih169EbgfDbhDwLwU4IWIAIqTfhiRtaCIAfIjKZORJooai6HokskAIE57kofVQtB1Py3cWOuVdWk5P4J+fncqGuGIkGJtg4FKRymeUFIFcMGAkOGGUcGR8wCGBVNFHyu1+bnGXw1gMXspuK8irfYcSgfaAAAgAElEQVQIxVJr9/oVFCwrmvFKRyDhb7t0EhmSMnfyDMT3LFMVc43nM+0ylBlGZ/hTQMC5rjquUWRBCJ+gFxsNaNyFqCs3XWtnI8EmGbBWYoXndqOHwi0cYFSUHj2+oXqatY1HOduFg0GmGSjL5WgXp7Gs40JFSSXFDGZ7vhF9o6VNg89akO9vHpMB7DeNY65qOB30F2dhcsh1YZNZKTDsHGXJhbN4w5q8VukM/KBI80nJ6+9BhNvCMo8tovFqxUZQpOrkejyDsqYeNlZEKlKGZyAjq9OBZKOQCjocg5GSryg9C2EbwnjXBvD0GthZ4HGlwjpOOqNjcRJaRD752tgYeMLyxvUSuOJQshyeEahJJJC9hcFBJd4gXDWijHW44b6qdikVSvX+0Y6zKWtljIFnzkdsoYFW5FA50vZSy+BSETffoVIVk6PMtHiuL25jhbu0UvBLGetllGpkNNrHdP/kUQNAQC5YDEx0u9qHaSz9MV1BpUyx7OsgKtel0xpfc1dq9ajKFtBIpVOQyGmthkacbT3i/izzMZUrWO7tlNrsMY/XzsZy63/U6cyNS10qoaefJ1Z1ZWHoYYWt5xmf15WgdRW4xtk+2fSuxduCC3TmBBXRAS9HMuy0DZi+Xpf9adHWby/wa8wychzVZjzvxXnvZHwmaX3T6a8c15R58b/zc2rB0hhszlI8FKLeYFNy1lNQwDDRzDagfDI3oizQO5vzJGqDe91dcsEAAMqOtqbeGbUsgK4ydHaADnc6M838fl2+c1SEHujms5H1CN33Nvi051D6Ctk73nLeby1ZlTvglVhaOaIr+CXqdO97MvSeXP1Fo0rnjArXTR0DV+LVBM/DyUOQkmOhc4G94cSbDZLpjCQNGriBwFwXWd7tBjOPdJpaAMf+JO35RfbrWPDzPMfNmUTAp8CYNN4VpPAy9MpXBEWDJzjaczU26Igt8hm2CwKkKpN52CPpVm6k69K0p8ANKLR5nJf0VJkTtcqUh0V/RRP79UuHhDI5SAdXO1EOjx6tbL1qt+csocNMjLAFwikAOSoANcgxgtwcbMYRKDinnR9nXFiXtHMEoDtKOJXsG7MUW4YHTqkVwKYIZq8GZhvEOXSpIGYtTDqXwHHyCAaR2esI8FslQWMmVes//ZLjFkuXZV+JaNB7czx9L0DQyDDhWlCXNQj7mtHzApgDiI/7DNiHfepywbSVeL/HGDo0AXDtgOaC5tVq3stWN97RWicGN71ixH2UZ4m/I+P/9Uv0WrGTKfmby9asBOKDh8ezZ8+PG/VGsKMrs2hga4m/BHj/xj1ZDgQFIsv+0SPQk0UccQVWabCOhHJggW28ZgBdArKzMZi2pMC+lJvcWmbwSPfTMSHXX2UyMUgyzgmBfvatwIq/fnM8ib406DPD6hMYE7CLwh/EJZdyZQ5AMy34HrA9ZYhbVzbf9wk3q4n9NI3lb+KbCEK9ucHYMxtAFTDsTLHsIC4TjkA6meK96E8xN5xW2VDaqFw7V9VAKbzo7aGgTKh4qd9SToVO8OzZ+3AUxLOfP3/Osn1pf2HjaFLp+TEe0yYdrrd4D7SiNobe30KCMRkiMTPTYw8eJO/v5DI4yxa2V2x3rCfo98UL2cTxbDrHcdrFz4J3Bi9gyS7vcIFuLo/m7A5kTcXaq7RXBhsHdiQeP2QXXlRS8OQJqAdPfHw8f/EcGBj63Kh0XlQ6QZmtbFj/cBkokbogAnBj/iy7R75ju2oUQoNOrp+IB3CbE1twL9RFFiTm8bAF8oXuI/5lFYHvbzZiADuLzP9yCCzE80Z+Zpkz97KJvX3JNXD2k0tPxn7BkargA/NqYpAX8vlU/s56RA3qXUbFfv3e/fIpswI+5YqooWUuI+XsqPiKz7tN5acM6u6UWJ2aUmp4qFgzE7VLDwKPpSbWwXMpHwI7BKNHwI0Cwo6FjEbQlEIpMMBnxSzeDw/uwTp/EKKIOmEzMXupg/FYmJYjQ4YkIt0YMZkOGgMaEUHkElOLPUaa4CM6KuIZXANlnaCZ1S1+R03Hl6wXuQOKLczNtGMsqO2oRmExF0ZYMX01zcfG2SCUbRyXRqK/6KywgwIRFXKqpCPAZbgUkTWP1deF4hnbkuAAwF4Z+MvmxKaIbnh1HLo7jKi4IAVc0RXDODp+PUc1LZDtAcAwwNL1cwOY0upmgFyhCblvqxNBpbEIpEew2TnA5/KX6MshVUtaySTAJ2dTD4ToUUswnrM2ojJ6MppuzZT2jgqmt1MZ02TQPG0d3YId1dkJxdyRdwZ9/ZzxfQX82plZpakYfUDhbUdVL29W8xlAvals0EqP6HtWtXqpmA2aQbu5sIS+sdCMc8/yl0GBntYdpQdqTWF8Q1Ml8v8wyjt05wS+5jvOoILfODsq1trT2zkq0g7PCbTTOhB4f9uuEepMfd1hkQDSRit7G0dFsrnG76bjfZ5P0rm20uC/ygoY8GJ0DWc7nw0aw92q8Po1cGR+MwmBz5Jh3MHP2anT322jk7KqxtSv2YHw54yKgfvMLtOGpPVdJNjsyMMh1Xyi//X7RopQgk5jmuY5jboafZwdFb5ej6DF257HvfvJdFQYTMBZVvmNJf/NUjMa/iDTx7Pdgc/Wd1lzN0hu+tA+qwkm/6VmzNK+GMG/5h8bm2xxngpsGu4R4I0ITzhrj+ORSlZCLoueyinJ0i89S+S+joqh8XEjtZ2jIsEdgVPW/eoMNV6L4xrw595RUVGTLHfhEwb5L+cQdqcFx/QTAWkUwTAz40ywUbsnIx0yAkO0o8J7XRHzrm2vR7AR6oKndY41718Ciadxrb8YejVBL2pncoeSb4zz+zgqSldpr+pyXAAhdV++CP0KkMVQvHSejUESOyuga6Fv3NpxAz5jh5yj4a8yNnbrmSWeJl1MOoJvu/S36iL3xLOdVq/cn/dB5rh5rezI5ZCVcW1bIgKhApiLD3uXsdRUldjZdBdt9kQHbgjICxhVGZzQa/C+hRMNdsnpFGnfldViPZy0QL3XsqLWl7KjZyDbTozAkzjH4fCqZ0RGucofTsFAMSaU+BUwBVvwYYD/to9pQJQNXj0RASRHCRr1UTSgaIPDYGKMg3Yx2TkcZrnNLDPjT9rCi55dxbcYvR9rEA4KNMcNJ0uWPiZfQxPfAMJ9YBqRxFfVyDtATtk9OofpCJQDgXtK/cg2dcwzxhGgtQM0qhwWHWTI5lfWJ/pAqEl3ceFG+S3rP2VD6mPihM3Jbgd11+H7OrrXguVy7Mft81uWiVVGErMUuBm2k0Bb4iWWjf18DQEtArWxbwQ9YEP6TOGstTLCCHqSzmq98bVK8Pgd5psIprwhfcGhIhlFeqoMHQPU7iETjgDzisiMCpKP70g/Zd9Y/6IcjEBYBm+6hw2uVzYRg0eJpaAcmIJbYzuwnnDsSbfRRGgDE7txlkVkKvCMMSCQWV3lgIhrwwHX9Z6UvJumApFlUh/z5gqinHkjaFT2LNdDVSbkXEEGkINoMluM7xjsSpQ0I413+4BngJlvXS7BmaHz1Pd6ZxvwYuKFma0CJy6dpnQ6y0kkmz/GcjvRU/LNzLDiPqGPCPrdjv3d+nqtHBUaFtdDOgR4tLKG5vUGvaL3J9/LDFbbWSNfLp0wdKizTtftvvk9O7kLXqn5uq8PdNyomKdyYDjzKmlux1RVUTHPW82svquA6pbB3TC3d46K6/V79+unxApIM8naiNeOii/98DP2msgazMWsOJ2VBVFmzaAAKyKkM0caUVR2EqhFxkIIklcTaF9gLRRVMRkCveVU8PNdhoVR/Uy1DKcAGJZ4z+zptwLE8fBJ9hj3jAozbjP8K2dF1nRsHmMzVjtFLACsEJ9IRcGj2Ug7GyF5D8z0Q6GgYh0ebnHxfFxMqZcM6bv38BFTuWMx4xlIa4zo/lYSwgIVD+zWq7Ud0ZUblrEMFhUEGs4VAZuDusioYOkkZcYI7Xetfwov1jA1KOY06Jp3jwkq46uDE9307xFy2GNnaiQwL6HY8S4oiZyNbN7z9hWmsdhapROqTj2Vp9XeKVW+H7sMDuzt4uWE7A3megNoRSvvwMIrRwVencCCMwDMCUZewIgmRqLGnllBMijjqJFkI6IRP5+9XiKlXMqZjMVIzw8lkkJ9hMq9uKnYdCfFBvSeudjWUVGsc9jD0UkmR4WBbi5YGoenzbcBpmbAdKSGgVFXzs8n2+Ngcp7Rj2Q/KgBcu3dnBEnS6AYVms/8xP3RGHFa4/6kGWRfDkj0NYL/Zi7jHV059Xk/jTwdBTIc5pdejLfPBWuO9Hw7STmmgXekc6MyY8gPnBrGO9ZkaAYieskU4/U7vPc8S01RFw9KeYoygg102wLOK/oYdm9aufX1NGbc/JKAco1lPEBriswTXFHFOkP5S6+t6y9bze6JSto/RybMvdvVgF9T5xZH3fCWK4cMaEORhcQWmmNrfv0qMCCPxWhIdUeFSkALCM8cknQ0pX6GfkbOcoMUTNUOZ3FT+35JzIv+Bz1Sre2weBhL2wDcE4CL61P20wiegcKUG3rgzuFgtpU8pd+4Zi0cF2hDAF6CHZWBMPJNBmIs93tyZJZsSj+C2JfLCmyyGu9wVFAAMMgn6SmdDtSVCFJ2gHvMxKP+1NKZdjKzAZw28Xf8/ETKeS9pzPs2OJ9OfHpzHjdAarwC65wRxSbhtRBnMBOj/eNzq5rtLP2yjpYuFY3rSh13vXd99O6rQFBxn8G1BY5a1tfOcW3meZezYnRUcJSX92RJvkXJkNUWpVNFYKDK4qImPoLlGbjV937//mqs3suNxToxcl0Z+cjYj0CpytwZ1t8OnS7eWskav58ZvWPD4S5XvT98P3VU0w/A0WgMrmCq2Gc7HlaAPehg6OHGqPFoJotm6Xm2ORPacARXPSZnwbtsSl/Hnu1RJZGrhAzLCxO4I59lUNmV/BK3wTVsnnwLHf/J06dVSiicH0NPgVFDi6wV935kgENVCehBbhyXe444glplAdVzzA3dScMNBD0iQ4XlAWPNuCcut8RZ9A+zF2ftpOkOU3Ucco6qDTbTL6oSqHR2jk3OaEfhh40Eu72Fy7NaAmnatlMfZ4L97cyWU7aCMCRc0m5zCV4MWY3qgXvMwLJVUgG/xj+Ip3BNvUopn+UQoYOt9WNQg2r37/Sq435jP9JK3LgcwG6rEOi5lYOKem/QffCSdPY0eWt6zkwS9xFBtpwC76SvVClqnitmmWCARQ0Y8MaRmsrWSFOg2wVTQybWG1bwMH3jTtC6HC69T5pGMzspwA/sMEpeWv2YHgcfUfnwfja6fNniTnonHJwqbWdHUpatQnPwKl/m7IZ45+rjiigOjsj/tjVayb6Vs6KfUsgRBQvs8DjawZQLxA0jLIclyVN/ykEH/3OW3Nla2fHGnfwCX0VzefJs91h6+aKyj4g38UzE3+mwG6o8jGUcPdzZHs5/Y6alw7xzVCzJ8t2Xn1orUIp6KocXGRXhqDAYYiPSqfec1wrUolFEpstrrFhGWSen6Lr2cICNADiiqbCU8FEBBxSTz7NiRqPLDMTeQ0WkKSUNQDuAcnqvq6RKRX8yg6DAUPKJKlHg2vVlsNCQpyIbRk1ER9DAmT+RUYF+G46SE+C1EwxdER6epSgSsBw9y6m9rGHKdWBkjVJHM5xyBHOXjgowQvZFsGMi5hdCCUxfj8DMW1QYAyPq+bPyHo4hN2uLfca73yKjwmAFA9vVbFzN2WGERkSWBHWWGJpLVWkhC4gx5YqmVH6J56G0AQu+MiAS3xnWA0ZIevTXJ2JIq52ODKJmRBc8M2NJow4GuWTSYGNJkeLQbUlyHjbWiEE1wNRpkwuavXJUnMDmBpD7Pl/Dmuda616qR/VY5/dw/UPBJdBinvHqpfvNKDIr1AfV3tw6KqZ5rZS7fskIqJfBNnrjygE03tvuBh3kTqSTgjxlySKwZY50K0PRUfVUp7SzPHvJn2ptTdFDtGp73d5RURcNmNQVQNWn29/RHBVp1vXamBeOIj8GsqaBkv43aXlcxK6YbZ0gizENu9AdSsOmNp7ZDDZLNu7DCNEV3Z8dFZgTFOQ5dXc2kgVeM675ZOCseG1mrDgbyxFDAoFQvkSA3Rb8Ojmy2rgWxV3X9GSZOjoqRkN0DRTOJyP3utGMRzQ0ASTDzNvPR6wBDINOYif0T46jgryA1FTBEqFz7IzgHUOLx6wdFQAflE3nCOEEVcyjpJ+NOfqT/BGIu+JeS1nRgW7dlDyMXtZhv7AK7iEhcFmukowE7ADMhotefn1FTzu2bOAmyqrEJ3QhgqFnvsvdjB/W0XckUzWzxBwJ0ENarBwZC7VaJvYJQiuNg46uLMkjYI7PJ61hHTV+Rpjy/Y4uJAhU5Tg2XtVhrbeOio3AK3l2nmQvXTTy6fX27vpgCDqkE9e9pzpgOu2hI1fjLRWQpMCTlYkDsNhSt0e676hJ9NGyWaHPBmi6cwLekfmKt0+vG/n7fixeTesdnYZ0BJcLbkqSRzExJurp50/StwWnyp28eHGbjcvNwg2U2xabn5ZsXjpCnB4CTG8QHQ0Zq7r+N0+eYh9XTqY4oZVtZAZl+7L1HYjoV/UXIHg/zrDbaniX7C4GtpFfGGxnZgUbRJOXTUQl/cClgoLPhO3kgBxsdSvtGauNaxVEaBvW2Qsca/GC7sjheo+OX+oltGlZmk2Oit0ZRpBQlF1iBHzsHSoaPI5yMPyOQBtLQeGd7X+9t/H4GHM4OVwqyKCrMz5KJwzAt4ie5cTIbwHoRQS/MlP4NgY/IppczZnTPn1VGfrzXqCMU6op3nNz65qJnxXNcNNRofXysrFMUQukA528Pm5U6qlHP6ejQqThTJngcQSaTyeiyY5qlIzAPVRriDLexAKM2aCvgrJ8cJZVOgwyoAV99Tc5UMxyxbI4nhnPx3mVfulrsoF7q0Rh50XKu6bTmx6N11hWIkdxCkxxSa+4lr1MmYkDp45Kflnn7DaCQWCqPA6EkO6h7E2fczhUOnA+KC07HW3Nb3eOitDbs6TTzWOWrQKmwT5A8U9iMSGT6MCL87X6UIYTX+mlq8yjWJWgeFzQ/NuUfsJz3IBbDqhwNsf6s/E9G4rHHsQn/u3yuPN4E7+LM4keL3PllL3zfpAzLZ4icaglflgjiIwKh0YwOIFwVGIXCXSRf5APrnS6hfC1KNmIXTtiY2Njj+yoUCLx0IfKdGgMDjxQ68VxLSydxKD4W9L+O0fF8sy8+/JTegVSAlcUy4Wj4iOfT2Wr0unGfhH3dlQo4jEaY7G8kSMIQ1OR0SbAnZ5slkni881gU71pil6ltfe0VoLajNBgU2+WisnUyKjXbyMGSlbL6pCyY+Fp4D4EBTMfGKUa84CCFArjJt07mHlkJsQnDUilr/oZZkoEFir97URGEjSo5ai1CYF2c/Mk66dS0bSjIq2xfFQ3jIeIYRlet7eRSUGlGul7qHHI6CQ7C1LHLh3u7KyQYULjgRc+gqNi0eDxIqMCPgTXBpWISaGiPimsHUtjO4WBlZEUS3Y+jcCWoAKtjzMb3CPBzqfqy2BwMvVlOWquHRUlVBJwkdIJ5UP9VgYQsm1+109t79nYsbMRyozACNxax5wRUq5GZKcMPIIbC3zDv16fUiBH0CmBEK8molKoiIQxwsiwqhV+eg2WWVFiSlGHQtWAV54P1pmGU65FbdxrNhuwvN97yqgQwdsUn4GqU0ZFgoCdb1HxWX0i+s+lD6zEoJ9INvXiXfVv11gujNb08JPqqHCviqYkrebbjYeuUPnabkTbSO3PKUc11/dKaRto3KAsb6ITCQPg/8h24Vo3gnDEJ/m0o+DlGG+Y7uCo8LjgKJHSCBYKmGSxLFaMR8dv60OpcdXA+ry9Johs0/QImFST585fxgEY1uvftgW4l6Oi9gJgbvaoIN/1mSVrasxpw2saC+O823WY9+TA8Iou1PeJk9aZtOPIAJDpbndOSTZrLrNbW0byLSYpnzh+EpBKJ/SYvu87Mec+uWFB7nZU8Bxx7R1ZWnSudM0c5jhg7tead11nMbR7hhJoEup6n0NCcmmtO0yv9KhwHrtjrb9m12PJZ74dbj9vY1cyExS1k1nSJ5agl0fpuqlCArbrlEzFGZrNaWBwvhuWawdQyPhVC/g+E5dgEBBpfoM1nTIqVJI19pcRiAwAoK/9rDvujurbOirGdRs4+4bKdju09/6TB8pg3zgqZn0rgBwAw64fjyjgKnc5z3/QAa0jbKMRmKUcPBk95gzmhm6zU1w24P9pH6blKblwsW56SGelOfQrT8WQOSLAO5n1Wq7BzhK/RhkeBIYxap1R4bT/4oyx58SOx64dR3F+up2CiHHZY7vST2eJJ/mFwDY3lx7H0uWtZYXBOstZlhdyeSWW+mJWeQTZvEbJKwa1TTz2TYDRLF0cNEJHTpxlgtxVtq7pKUDY1DcPYCEdBrSBytkQfMyOyAAQkT3Regb0XldBm2iQrgyLHW06mj9mAQeu3gH+1PpAhqMHZ2gjW5h9+SbL/Djowv0ju4M1z7Pm7P4IVN+YWW8QO/5NALRaXFgE4DmDyDzLu8HtBrIeLAQ8N50ekqs0Yymny1aoUpgEeyn7XEFhdNpXHxFgBTb2VA7qzH+ly9AlU5krWgs4K9J5Q0dGVltQY2qD900sJu/vehr7kCgARY6X0FeAm6hBtHGMeBbLV/GdMY4AtI2xnLILGs8MR0qUjba8hF3U9O54WXCOx3FGoscEegmFY4yOykctaJN7r3MdNIaMleJFxG5Y3qlnXEAlEy3lmnenxaXd3PU0reAm0KPLeARx4hxEuazoBxs2YWUjk9ZG/tr/FZhZ4DSkyyLuxLyAv0QQ68uhd4vnV7rvTsrz+57lg14iKvEdPDdyE+yoCLrr2TP9qcHeXYaNfNNN1mtFVjadnzH+JgwC/VnpQCLesZJFb46Xb2KczjrVmVamPOhlqAqwd1RQ5K3l604FcGUVO6jM1588fgK54L0ydslS9twzSMh0VKTAXW5W55PJp96Vfrom7He/fqqtQIEEBjmZZhTlRs49Kr7MGRVDs53eoHRjhQ+RqhIWEBIFnsS3wcwYQUPHBIFM1/3spqnWEV8VI56Vx5nhAsBW9Cv/lgKgNDEKaAqJNOYNYun1qWRLiY4okVC+4nl0DLh3xXmvTxkVYqRQItSfwp7tcDhUuuH4LMxTWSLMcmCUhCMmLNSgrLVGphb4KZAytq49Pz2xVHafPgnHB7EgKCjRCMyGhRttJqOm8sUgoRGAYPokDZIYF0Xt2piRb3so9QW9z2m1SikNOkkbmptHmuJEM2qZ/zLN6K8uQXoUbgDprgsvBxr2tmdm9BT1hec6HBWYn1Ikz5RQ854NsQQZBSwSQGvXdyVZoKcdY1YOC/6s+wCq6TylzquIyrtN2KsZeB9HR0XripJAYlea+tmcweraKjaW8jkog6VAwqdPn6Qh1ulp4ESzsXsH8DKYIS0F3tZCf89djooswuRGoaLNLQCaYDJrVVLbalFvQPJUXiJ7ffQT3aIncmNHqGuXUdF3+XQ8VoBBM56GM4YHuan22AB7xD36So8P66/jWBz1ptPd2AuvlVyZNMNx2BX9ND/fPKsbL7OSN66PzmU2AZ3MV8u8zltaKRtHXJ+jOT0XN4fLWGtFEDYzvwP0jQ85chNlGsP4jx4uU/1s0tX65K/gz5VxXuux4eOnHhVyVEDu8p6dgj9znIHPN15Og3/i7TZQRiZAmZAlF0uf4JFU2csEzKrc0Jn76ZsIn1x9NuDaLlq6G1XmhTSW946KpM2M+rLteuWo4GBN43RUlLTIczQY3zXH2qv7SwyDj+ZjYmdt1UZ5nDiQ+WUrbWN9xr0IKkgBM8oAik5XuyyPHd1snS0CUO0MDzA//h7kXAbRuEzKep28omRrcpI6qllRwaCDSYca+A80300ZoryQwChfY42LYyLLpFMqgTQ9zuViUKakNTYfdJXkHWPGzds7KjjYNQdZH68t9W34GWZuR4XPZr+2Raf7jeahVV7VoPP5zKcu64ENG7ybQ/U0ADBvJ+Zmcjs+2ek1bbjpleOyXJ1dnqO+I9ZHV7MADuvsAtdUT3x28R5d78CqAOLcl4K2nsq92VkblLkEmTroyMC5WAf3X6hMBZc8kYN+w8h3K0JbjuC5PywFVJ+uu85rVYEBdU5dKsWZA7x/oimVe4m3OIq261PGKckjeHYIboZTgUFz7AOhLAoaTzoDtK3RuFnOMuvicVn8FnZe/M6mzwzqi2bdu3Pqklbu+QgHLviagzk4DpSEsaMXDxvnHTZsgNNuBsy5WGfTJIQbkKc545qNwV0hwf0GGN2vSHQ5jGCBJi8gJ+T5mw+v9hh9gApw5r1l6/hs+W7KL+k2Q+ZNlR5zlHsvKZRy0lHgsu+jMbSzS3rp5Zkf0O5mFL37+IEOgiZaloM8z8lw4axo/Rgcxe9otpRR0tUCLI1sldgr/LdlaCCjJWzlCEKL8r56b+pcdpo8fHC8eE4nHUtctvOltQYWFOD3TTVkt0On28PGXex4wL+jPwXGIjzH++0tVaknZ5v4zLyIzAVGEhGjaE4LnLXUWev87/oi9cPS6YdH/cxxwEddiky9jeJSZwl5v73PI0DfqCGe84q9G+M10FdaSUWQrkqsBR4FKCmqmDijIPWCvWaOk4iA0epxE06JKE0Hm3UqlIGxblVlOtAQ+IGMMEkf2Xw85/fTNy2Lus5JPW/zcjTTZhY1+8UeR2Q0FCdotpZshzeLHhXM7FiP8WrolhfmY/Hf6MlmXcD80k4JO46zL496+GzEWsrmQW9DdYomv37h13zL/VZ395Z3379bgU/6CohE7fWX0LjLUTEOqxvTE0OwRmXmJ7Uglb6e7j7UXaOwKADKmpaen0BAjH9lrI2RqAOjs13VmffgqHDppGgQxOjmEBbuccFoW44jngtHhTIwXF+TCgMFZSqNmrTTcuN7RBZEGh+aPlXEjrMBtgy6lQyXSNwAACAASURBVFhyQzZnh1BAyxgVYG5ggvMQkC8ng6MUEO2gqB2LUjiJzNWsJ2LuPQS0UYME0iwY4h0EGTguKJ9KdYx/o5yW3tONAiqRqV2grAXURFrZsuOpQHSF3xEQsS8B1sXHkUMujZWgeQf7QAfq6dFo1ntt4x5OrF6ztUUyWU8NwWWIkY8qQ2JMu6z1o2FAYwMNyyKFUtEB/X0zSBWCK2gvFVU13spzpmOeZcKUJh1Tdzopjv4Y0pMKgtOO43mZup0GhN5CDb0pFdy5gRaW+sJGiUhfV69rT8eUU7dBO0qbZtR2Vywm5jmBhz4TNJx0XlqmU929Hl85kHgeGIVKQ8E1WkmTU8R3EXSWQTMIjxRZO7nci0XO1FJ42nikXGZj+nY2SLN5eKiE6cuhVYMBdYO7U7/wSXOcFlVOk/YtFXpFdU3j6bhbdy7wexmA7bgvXjZkNxhIwL7bfhz69cxPsPNkHHe8m3zxQTaud8TYeQz1zdmR0VTcts/9HI7AklKJO4npHA0hdD5imGOV9utjM9gNZ2Q23Qu+Q/43l7pbOSmKXGbVteRdN9Lz/ZtzDR6o8U6ushZB62erxMKOHWy0acuNDtINoMGwga3O9huW5OCHp4ONosmr8xxmvVpe5nnwfeu0/42fIveF+1GASdURL7mNa3JsIxWC7orUGkHGn1VrHDMTEEbgtUskAip8jFPsDMD0TRAfT52nSmHMZ+PeYKql+mZPiz8V3eGvBNtIV+ZplYVgMK0evDNSV/J/ns9wVqWfkc0IINSa5ncO0uCJK1nYnJlDdoIZdLPOOfLJuD4zTgELd5mYos9k/hPIqjeVnin+aPpE3fsx4CTXCLpek7dJH3t53kHeHNIFg92yAr+7rd8clNQf67MWq5Wl8frw2zIa/PX5SrDKOpze6edkUBACq8RN2pLtAYwGmEqXHEBvZZGGTk7QjJGndqDwWNd5zvcYTBN/YRQm9QoD1PslFx+EjsUSpACfVL7odN6pUChwfKTFdCJqE1O/bE6h6olRpYdmOUVQl7ot91HAkgJ5WIKNZV9REgVnUsFQyr4OlSDAWu4tM3CL79Phh/WxrHKwiHWo5izVjHMpOgjkc+TIcusQ8Vo3Ew4dn3vlfQ1AV43VlfkAsC8ijdVPypklCHySHeW663YiRPNe803qAqoVP9lGpVcwCNA9KrCODhxMQFYZAfEMBQ6e6FlrbDvRkdOxFq9e3aLsS2Tlh50cGf/xTvaGdJBZ7UWnIDpRuK+sUlDcwH2vDPTZtkpHBQB0HJBmf6ts0MNyGKQO+obAdDhJ/OwuW85laxT0pez01FxVsstnx7jAJKC1BU2nagEd0D+iIbyaHzszhFgDQUwDxHTCyKHdYJDIwInslaA/R7PTySGHkcsjy0mBAMtwTgkfwN6pIf0bNEUPe5QlD+ODiHmdR2fqdn3mzCdENa3HQpZhW8pAyr/UH5WZBPxCZ9MZEDHHGD+bONPGdunt5y+eH++99yE4VOLeiPhHyanUi8hT4xPzSAdnK43q312GCpkKWp9Vo+aUpZNoHvlzExRerIZo99KDfl7wNpedjO/iTGTAZ1YcYJaDHTDgVQ0LqlcRL8mxyv7qdLxyythZs9I6vPbmq4j7aVly4FPSmwbsRPyDZ1kZoMqycGAR+V6VAc55eRn1m51T9DWVTLlyVJBuC1NioLZ03mRNzUZZ9Xe8cFTsZG1/b1dncJ713tlB2u1crMHGid/3efl+Zd/Fb+96VFwooB/0JzJl3S2P3gd91rv7qHLhc09HxZd/zvNp2agMlLI2mRZ2VDQwrLtWbY711FMwT6fq5uMEzsyRT/h9jiDcG0o5Wc8iaamUhh7dGAoVUkrRFLSusUxBNEFE1rVSUWBAoYy1PhVIi+uCXj0wHC1gJ4W95WAgO7QDPyYCOAL5YF5ugmmRwf9a4UOE2GToWcmwo4IgbDHMAm42DoqkijVA4HI/jiiFcixFJFbX0VA0xsZ6oYUljaZt+aoUsy6gk3vFOUaUxSM1CCsDj8oMMiSSLjvNCOjhJqRw7fcPxkk7Efm9wGr0X2kRMohwUJOy1f6ifqrqFEeJsDBQbp70uq4t+tEGiBWCyWhlAkWtWemDAdCxhixJ6QHSZyMytCsuBoUQ0aVIiW4QnJtjCaBOhWt/Dmd+cUXqBaJYUXGgqZSJ/pr29/LtAx/qmQelSENZk6I6nqBzgCvPic+XjMOWWYUxaCDjHJmtxNRYXmAlGrWM7eSSAoa92ER8xeu7o6LzDrNf0jG5PflrGYcFePDsiewHEIoyYgOKdbBKZ4FK4phJ0fl+B4gbRlfvzjPlUddu9nvhiAw+qyihTKFvZ/Ls7K2Mr2T/dlSkM9Hl9CZxd+c/G/8TQOxbZkdMyaKpHBAesTs7cf67HPJ+Bcii76cxOkJs+LqVEelvIi2tGnz7nX7KPL4VbfTmm4vredBy3HaYb42Kzdqz9431GIJ/PsON/Z3jnU6OCkZMiymm45yGi5yldqjbMNk4Ki7JZFoKR/MZEE2H04Wjgsdxcx5bwEPxAgIfBPc7k9TKDcaX5H5ZramLxJ1zBGSf6z4Gb16RDdPWZfNz8pwqSpIAjeS390dOpPO9ezm02qd+/0iLLko1Pg+7IOO2dEQ6gZJvrhwVd/KSdoGax/azPEd2rx83OtJ6E8W6vgcXlPOHOuJZDIz8bHyr+f5yLAZDpJ92be5tdgirGnLKQQnSZS8dFQqsARjSSj/lONtRcgkZnx1n1xokcM+EXkqP2WrrWawap16eXzvCxItdNz4Asg6YAkyMQBZFwddcajKhB6OEFXoEEIwz0L/aIzuV3aMg9FeXu1rpaJ0Fke+WPUmbod5iR8XoqK+xDvwMOnM5JAKUA9DVythwLwkuMnPQY2VwGALMMtCHzZPdt6CXRbFD2nwfkfnIlpJd2aL+PUbPc9bh7RDyddZHYg9czsN19C3HCfo+zJLAdHLw/wzsxbIahKP+Rh7t0k5BFygTI3ikmovvmQxLjTCrIuYRQDRkECoFUAc2WM7Ar1amdxI9BrgBbrs0sEvmuOQSiCHs5dIlWJWmdGj2j2C5K8tDB0Y9fS+acjMCmuWsRrvf34M9BCj9pCodxDxsf0dJrdMnsspUCikqGbjkHW37KB3WeXEMWXNARjN/Mz9Dn4Y3r+AoiGdanns924nIP2n/Rilc0jib5rIslzNqYkxPnjyFvvTiJUvD4OzHesbavua8kakT512APSouqCy19RiL9ngXMlgyA4fjtZNIu0M79OYm38kodFedsNN+o49sdJW0RZqjIvuUtuoFXR7TwcWyeTdPnmRGR/wbfU2iRBKcGSyR9uz9948PfehDlWmE0mMsdxQMse+N6YaOZ4Lq4XTrTbXR5Fw818El6MewECRLEBkZRi3Qo9mj1iP8KK+PHczBu9zHoIJHqwSQ+W3YcLtKHDtuYN5tvTllczosDTm5lOx5r1NHs+ozXcKeJBOuJeyCr0mFE9cFvb3//vv4+r0PvYcm6bF3rjIAPuiz17A5O/owVzkhlvOOvWh2sK+Jr9IOPpX1mlJFdBP3ah0wfbXmq9+cneblAE620/Wv7ICr35AVwh1756jYy8i3/iUIN5jKz/2CDx9f/EU/57i5eXR875/9wePPfN//A6LaKYNv/aKfdjeUYknvncofbEo/fcXnvJhWSMRukGQ62FFj/vyJezoApfrrdpbgHl+T7GPpGeavZB6pAHeOudnPs0lBENSplV2A3aaiwmgE1/AsxbmafpM3Vi1SZhKwREBGnEjJshLjUgJLJ0W35uaV71bAjDb1a/UbS4AEOEphbkHYI1VsWWAOUbrF29ciDEqcrBYXTyUDnCwbp6+l8jZ5vSVXGGuUikoza/C8Ulu6oyKF+wTa2wFk5ZnzsqLcaHPAblopDEUAeF89r4qqDZ2VK4L5eq2hi/gsUaC6Pi2dEa1WvYVdU/xsjITCAQU7I6RnkKQiTwbjCE4ggVmpbNS9SCn0Hr05jpdTNkKtZ6uTqibfcWM4miIKbPzM2vw81n3phBUlcT2rHi+N9B7d2TftfOiHty/A9Hhnj6ahcVQKx8r5Kvsw2U6uU4l9yCIo9XZeAtw8H8jYLyq7bKhHmo9IJioRo2O0m/fzutpRUbySf+k6bnTaWmwa1sHodam2adCnLRqU2Y2zom4ax8zLLTv898hZZgcGz157YvDraAqXvYvooFyBpXaKZm8WP2iKkGdEYXfYnCXFRqT4FLefe0agf56e96CB43lnp+V2PY5blXqYlddLx/aU/NxP7lJ0bJppl748r8tazm8VbBOP119AbOfP1+vcl9l0fnY2Dn0OWhztmFnguYSl77PBDL/UiSAAtPyKyOVavB196Cjm4OlIVDSt/nYmaZOky6XYrW2WmksZzDH2jIoEdZ1RsXNUTIeuwODVfg8LfI/tsyPrvIbcydflT/XxEQES2KmSRtyr+5cIkMt2va76Nke1YkTJX3UeZTT7DArjx1Uz4Hi1MFtHj84HKU76y72Kpk0ZP8hIXcttPrd5JuzMXOrwcpwvyX/TXNSOil6qTSt0D2KpM6OzmGvt/RrK0Z6f2MFlsB+dN++VI8E7yEN+VNGZfmpaKKKNXk5mfvMVyLCatzMKKujFoL0iP9XnwCZUOqwamGEsG2A0AqcsZ1RSdxuJyVKbvt7ZamUITCOeSKnP1UBmrpn10KXAWeyX9JRwQrARNZ1BMSZGlbPEUYCoKNuhvgyMGg9bLvQqOgEeKKs67DvXVWfQjSdQE7HjeMjsbvOkdbDmf+yNUdkfnV/2QCeQsLNWVOvdK0DAUf37lEHDgDbaAgyyegzHByLdQ4dMUeQycvzCNM5jdj6sAF7VAPnm8c3xIMpHvWSPD2d1BF94+uTp8f6LZ9kRZw4moD7JJrrIltfyBG3aqeCgEtK1n9DqyCv70liO7xsc93ImmPaRnSIHlkH4otkQ53Q60VaPklbR4LtLSC1cqz4U1wPod2Z0Z4k5sQrK4lkrGQu9/iYC5ZhFg74c3e4eSIf/cDYLA/noqICDUusX16CPi0rtEPGVXZllYBmkyEbZxMSiUbYdML1PRK/CkLamshWMg0QQ1XP1UEGzX51DZrBHaXAFFDZ1dcfrtrqKo951IHCu410tyLMHSNlBEmczsnTsvGOQC5uoo8eB9gROmMcMzvAe2dGc+I0z8pVt57E6ewOVH9Dnhn0dbl+8ABUgsCycmo97GdPiY1u+nzrmmufxWyrIeRYOOgp7jwLQhHr8mPZVYoJY00ZF28laaL4zBpEYglUDZSlcqb3NgdDflWWwZ4+3qwI0+QUHWvQceXID/nH74hZLsnJQli4rxcDnUUL+AuMfe5tZj5DTEud6WEOducXC4rLNi3ayYq+/V7Z16ZM9eHfcQfL49a7u7a93jordOfjA3wdd/1U/67OP3/gP/dLjl/9tf10BOK/fHP/Ln/6/j3/rP/sfjz/9f/3QO2fFB1phaxQFrNILue5R8YlxVHRDhk4Kew1xqJGW5Mk0IaChWtEpxU4MKpW164WY7a7+PCs0vR8BHRVs8hOCIsv2RJmQqbtpPAsleEJRfhlK8avj6dOnEACow/fgYNprA2qIZxenuQac2ty0RlsHzfR7rC1AVDsq5nf2iHxEFKhkiN1GTalYy6lVJK7ErpVv119WI6BMJ7bwTsDfb7ino8KlmFpUlxVWqMUZfado+RYZkXoBtfnjgUvHDKXBHIkuiMuOOZssdjyo9EM56gmsM8LDJXFYi7fvs/ffQtfKuY0blnVySZI6P6EAM7KPkXL08hhwsN+xlaBQFlo0tYbRp7qxoGPVot7RnxvzWsE7GT4n4G6kklU9bcwXB+B8ZleOiu4g6k60ph7mn8PbW+QK2MSsLDXF0MpaOfDqSXBUGKUYhmywlBHH7OPCvgBMre8XC2hqTfRclgD7QS1b6cXBh8PIYmQPl2k+fS2Ssf1GWrLaW2mzUGpnYNJKGngxPyvdJ09lOqarT8M8stnRc1ryLJPCp67WCOOwcTbtrHlsj9CD46eVTalnSvEv/aw9rYCNGHM5qcth8YFEa86p7dcMFsBR0Ve7X3umGVxpUpv4906GJA1MG+B1wuOG3zo9eQzzHEYavDtSe1pByz+9mzZFiyJdLfiZgESoI6Xmv8xb/Kwlf2q0J72nHBIVyWS+XLpC1d5eDXVnHIF1cMFPpyxBpWxyLL/sWzlDCnGZzx/pg7qWzxV5TXzd19DRup7/StrvLKO3OSlrLYKn4Wx9mUa8ei79RACGYF0vJUOf9lq2EMnYjLUOzHSB59xv7Lpr29W5rFDP9ljKjz3PTfKVl9VNSXPv5mm0nhOua5+X3OWoyP5eNZ712b5yCm0cFdrXAv+dCbW1srfEhPCMJoPeiurUH4cAvuSXZLFBuFxjBXAYHK9yGIoCt0eAJ2opM3dAxQz2JqfFvARSNZKL69kvgGfDgHaXHjm+tqQAXLPXFZ35BuvmdQs10JngjrQn77uIFl1sXwJnk5NnYMFpelqradUSNClIBIHMthNRKtcZ6Y8DrIwSQbRVMku4Nc2N70MPg96qYBQ3JiUoS1CadgKzDNDvb3DmlJwAn2kNV7umxEh06uPYQ9k7BhRnOVIyu/FkZYiFXhP3B/gffdgiojgi6uFEUImmAK/h6A6wtAGbdTYagDbpHpiz+iCEsydA/LBNHz5+mP0DgqBj7OEg+ej77xOAb26GQYxFmTA7KvIa7m2VZIpshiq1wv4+TRZGfXaB847sL9qzDkudKWgDpZnVmyKeQyCbTgmW8mFT5figpFMUoLcA6cT/hrb8KJut658JHKaWS2yKF3lvMf7oARLNkHuUPzIm/Cz+t+tmDJCRA0BBS9kLUiVlY9bIyAFtkRf0vbYuNzjKW4lJVkzgehj0t61BelDPUGTZ0NESmQu2T8BL3F/S8qiXQG7MqOujW8C04j84JjlV4TS2Y7PtE5pji37sLDF/dRaOnTS2C3AGFWjpHhp5rYLFnEXnINTASKIaA+arvh+xaghUlfM3q2h0cTc4i9dybRuMkPtU54E6MRepnDPcezr+bmBfIlhbTahB3jvQfCNqU1fSWif4r38P+ETwviwZWpszqFOr9wQ/XTgp4jvqadPKZDlgZo4Zkwt+FOcC82wln0i/XCtiBzxgH9RRwQM6K4kbvbGdsVmm7h0V85VmTcrgxnpVkMQOl3nnqFiv40/ot8EkvvBnf/j41n/xHzy+8As+LOWshhAH9Ec/+uz4Tf/2Hzq++3/7/nfOirfendQWK3rwwlHxkc+9XbyhDrNru/miOaOCDLAb6QRLy1ERjZ16KR+o5PVOlBOZmIeM7EHx39vAg03uZ/le1pensDZgGdHmaBQkUNiMD6AYIgBkVssbHcpTNPOKCBVnUvhZBnm7ILjLMbH9vc1xN/f+vaO+HAlA0ITRUzB6WoNTCHYpkY6+8Jj3dvbZUTEbk14HGgiOhub2OjLFUWBm2zlNGXBpuyUZScmXQM+1jQgIOY1sMFjgsmzE6Q3H8fDN8VDpyFdHqe8fxqOoeQNZeHQqshwHv7Kgk3HWogBt3MVYo+yT18q1RbknYyYGFcdH7P8hYywj8uAMqlId7pgRijSi0FT6ioA6hX6tLSmHQDsV7J7ui8iGU0bFLNjHQzg4KloK6B5MooKSSpL4hLZZEc71Dpr3pSENcFLjGfN5SmUwHXLWPBfAlJSn8byNwBUj3h6yr00vf2BniS4fMA6dRYAIal5opT32PSLoaMisTl/NugPzeV6DZ8oIB02GMbThj4xYLIB2pW+ODpzmBDs5gNrenN7Xs0zca2bnrOijqAeFgs761BWV54wK748NTzuYdkorntVq+BIEqvJoby1WhxtG+jgpsksQqMruzYjqyuEXe/JKjsqUaQnkNWOil6DR1zZux0jtGZgaZfA8pg/qqEinEg+vGfJmuS+E+uaOggWs55jpx/rOmU42bNwrah5UH+C1o2JHL1kmYnYMAXuUTJCjmZHS+9o7+9WYT+2C/hQcceWoqFJiXb/bByNcgRHn9TATvDpZK+6jqD/wGpYpYhSqMyoIRvbazVtgYB+GNjCiOhc+E14P/rd013KAG/ik0G/fb5zyXoUdXwYlmj7ssD45nPWUOxwVq73wGoXDp1MLyHLTA64/Z9z7C0dF9hhrDrPd843QLEgE+b7S4RD9fweDrvmpF1qCwQTEKoNAwRuIXrZerOwqIQJ2KDKqn0BWRjivxnrX4KZ7GMRCGwQy3yC79QfpgACRBdinsz4JaXpp6/93Vdc6smSjfAqdIpz/2zoprOdaf60hCZydCcxkK+dLLofA6OyR4V4pUIEZHQ8bC3X2SU/sQ6eMBEWgA/DXWrFZ64Pj+fMX0GtZ8oZlcgaQFiB3ROO7PKzOuqviDSVLeMj7fLlu7ItX57Z6jITOEkFv1qkfPXL9fz6HICij2OMT/40xl053wGkRNAAwXsEwjiy33jPh4pNWwhJC8XGZ2V66Cg4r1Y+P9z97/vx4GKVKJ8ET6+49iDVzT0BEQEeZIkXlcw7Ps7QTdNLgN00Wxj5BJ1DAiIH67nwwfbHkFyPoCSAz0j8bR6tsk9eM5cBUemcWnumoeMAm4irTHJH04Mm9YkPstjPmMRjSm+cR+jsyN0RrkA9HOC2ibE3sZ51N7086AuCAoIyN57lnndc0dFTQgx1TclTQNOakUCrrwUPsg3su2KZGZoArFkgp7vY25qERvnrJ7CADycyOkbOlB5XMPGIKvPR+zawRskVltXvGg3GJjjB7xWKd7AiMfif4G04cZXxIh4dcjhJajx4faJDd+hXAAaYMM/e3oENQpZC1l25C7rJZkZ0R70eJtNevkXUTTiNbzaln2MFyhZB3S3VwbpTqwa9p78WY4+wgUFbyhs4KOsVSdxRSv0mCvADtRwyr24Cn/Yv9bT0OlqJ3VSGpB4C0NeoYUZdaMefYu5jjTTQGB70IP9GFH5ejIp0to039QBkVfOGJUQznt899KeZ7OcRpoXbkEZqs+171tdnhgO8cFUsK/In7Ms7jz/3Zn3P8a//03338zV/0c4ZmSn0Usak/+Jd+7Pg3fvd/e3zX//p96XH9iRvpT+U32YC/X0bFx+OoqIPmJjctQlw1xsMoYnsKKbX1pzh4hwihQYyNIFfRHtP2mIknoIPfq1SOG2KH8AIgi54HBIJZ8oaRDE7DJfMsYOnR40eISHnylLUurZd0oRpiIesM3kE+OwalYefdc2bFynmBOUiBixU2GOEIIIO28c5HaMJqh43WSF7vNUhyt6MCT5FRgbVRmnYKQwGEZfjeL6MCQLqj4pRdEPOzso3MA2XDpDe+g0UNv3p4YSDTRuTFEO2ScagNa+NSO+LIi7CSMqJNChSjH+pjJ4WjiMKZFM3B7CSISBJ710t4VYksK7YwXpEGS4HOQAVFDup1+E61TFNZlGFlIyFpzuuqqBIbY4wymQmX4F8ZtjNgUYAClj6B1F3Ua9Fc/JWZI8Nrx7jEuxwV41lyw3uly+c7aGT2SK5R3lTT+zpzNJIfIiKsopyC/qoXSHuKgQPX2W1R1IyWUp1URIbFYlEZFZQ5qzzldEuaLiDQDkBHTiGdeKPJzmn2ucVNyeTWdbCuCKHORg1x9CsX5+hOBJ5/3jP7oduTitcpDRiGMfp8MDWeZ44RVDR+SEN+5uxIN3O2Q8wNGN+23mgfY71rxdjPnJPvmr/fOSpCQla5qO6UsDOWazhHHPP5vcyfd437WY5byoBPkKNi633gmTefwjxy/9fSZR8Cf15naw8NElDAQ3v25KhIrt4CvyiH7EjrK2ZHxR6UXe0+z56SGJojyRFloNv8/hPjqODzztkRljm7jIriBVVur2llq+ld1tIdbyj+tHwQfl5wuwaCZGQozrvK9kmvCh3DZSHW+hPiMpev7l926TKeiU6jlSlp54lNXzvhMQYhQDxf63dvdT2BSgniyHGxfs6VDIbEn+ZN2eIgHfJOfnj1Opq+n1mPg+flno6KZJQXjoYt2KPAGq9Dk6OrTe1OHgfkGJxGYJLqnjPwowVHWIeSMySlXnMW+czue4as93pXrtg95rALppnYBUeRQvapvJB00Bkkq9PD1UCdevWrQDkUBc7Ma/Uqmiun45/17y8dkJsjtLuH46yz0+k392iat2t203HCrIdYmwgGc+Zq59HOngbIrd4haJ8r/akcMJy9MxcsN5kVwcbcCvHghQZxTRPYG0fs0sHgngaWv3Yk8fiWM4M8gA2cCf4yej2us87vbGnTI0B826QIEmImaDwrAOybJ4/ZR0L2KN4J1WLNa5lx8JKR2Y8eH2G3+t8A/tUrL/4L+/dBAWidbqAtSPdC5ohKD8U1YS/bZoCNhhJC7N1A505l78X1lI/kX8hMDpstIsZfVRN5O28QDPgoShvxN2fV8H104sW4qYOTh0V/iqHPqSciR0XYXbfICuH+48xhiK23jRwVeatk0uBwgRximTVkJdw8OT72sY8l4IrzWco1yyhlkBBtD+57VGBghYa4JtY3GmU/fNR6E8im1kDVl1HBZSr/ZAeUnaum9RijnR+eD7QFlNt5jv4Oz549QykmO1B7jwXKtSZvNKfULe6QsLY/PZ4OzA48zMC2jE7TapS2CjpxyTX2/SOoDZoMmpYdbTwHAPiLF5hj4h8tAyvGwJJOLCvnYCg7dMSS8Y7YG9t3gyyeswOGA9PkfwL2dcFoP/icB2jPTKq4GzxaTsSyXWgrBq2zKsT5s5U5crQyqEI8o7HqgZ9vHBXJ1YNPLl6fpZ+sgWiNslLAnJWg8xP74YwvyK042+ozEr+lgxLO5hYYMvDnxWIMjgpQINl8O99UQ2d5dZ7clSb5trZkvG225a5k8DtHxR1M5pP5cxDv5332Zx6/85t+9fHzvvDzt43KurB4cfvy+Mbf9geO7/yeP6dIhU/mCD9dnm3Jcj9HxVd8bm+mXQZN9D9wZFNFxY6toAAAIABJREFUs8r0b8AdeQGFLv7KBnRmBgSZGOUvYR73t1RArryu9/PE8KncN4aDawts8D/PYBg5XDzGDgQ3Nu5mJRQ2GS2Omo7HE0TlgJEmrmgsKwhmxhA0iirLqH6VlfK7wzD0bxCuaizep024fCxNMQv5GVSHsqO9oAJNRbmvZzJERS21lW7XjYBN3V8gzNXpYCQ/veMGxrFLCRBRFah/p/SR3Vbv70LdgGwZmtwLrLeMCP+WgHszSq30w2XVpygSSkW0l3GQodxTVe3USooOWlZUDQWr5tMXqb0yxoZILzU5c8modEa0++yIqN+4duxDUMZRF2Y0kkjnbSXhkCuDvsZoIyDPow5RxxD8zH62u0GKUUEBWoGyMqhMYUM5qK4WtmyqdoBHV4U3a0W5PRtLPMI2XDca2sRWwJEbwhtIsDHL7CnVC5auxxrKr7LJ4cC7ZJjRMJiNyRaxbbAix1iKE59X544lMcgdsN6JMQls1UGTfXg6pkO/mvarI0fLVeL1E5NuPNf7nor7xGwxXz+7/TZCGGePRd6j8lSMoKzMIEfdWTG0LBgUaAodEFxus3gRoy2bY68125sXqpHL8JMBSfMX87Xcp03I9KjozsBwOUcJG05XJw2PTCvpIAHfc2mNVM5zH8w/1o4Kwit2VBWPQDbHuBKjuMp/cZfp5OVMUmYnww/HKokksxvFy85ypSIAqQqUziGNBucDs8LyzBmZHMt8ovye7jyb+R2nVLpGjk06yXmsjor3eS1Atwz73tfEa5X+cJ/27XjJDdp8+lhWxqMiWNtUzIXbO8bVsf6SM28/X4KaC/oYQ/z8IDnZzdra13mOes8VZBZo381bpENyXtvdXWyRn8NSBL3eeWOmI9iKdRX3MpipLIoOTnb9bLVO+bt2eQjJCccLQDM2n+dzIzNuNbfiH2vn3kgIHD51BgOsBdCS38ykE2/tulTn3XsacE8S87PTxg7hpOQRq1NkEi3hzbM5SpC+MiWL6Kz19az7H8CpwXw2YXX9dciDeHQGI2lAAg7H0a0Hu3WI9csbD09gWsEKxVcEtotPmg9TlytHJEBaZHWyjI6zKGGjIBOWQTLYpyRbAY6isdIDvYqkiKyZnnr1cBRqOTpfmR0uktmevt9VJZdUY15BBz1wzE4mAzmsx08wuX9izUMXQ48KSYAswxRZI48N5FYPBTjkvL2wZxV9L8dbf0V1sTNHKn5R5Ydki2KNWZoF2c/Zc4MlimK/Hj4IJ0NkUYiO5dC2zKlodr0vQGtkpLPxNMvbVHDNrJ8we4P6PUF49Tt4RFsctucjNWTWu+mEEV9Aw3Y2GMd4BRhGlgD1z6IP2pQMAop6/lH6OD5RuspBJcFnik/UyjqDG/crU8KOGAaeqLSyenjAlgpHDRqSG7Q8cyvrhrFGyHJZsBX0LlETdoO/5VABMGC/oabMHicOkPH5QBBXy7CJZ8Rz4WCQ7evz5zmZt+uQZQAHnS/OsOHece3wbTX11jEsMD0cEFHS7Dgeh9MhmpwrkwClslT+OZ0jysygc6yy/wP0j6h2O03MMNJZ0UrTZFS/AhFjjnCCdPwntQs9aQqAg96sIIPZrqNOXY4vZFfIiRWPtXPJWR90MAQdEti3Th7rF+Pyd8wGchYmnWnx/0/few+85cWL58jgYo/JyHJR/xJVa4h3sxeO6KOAi6XwMk2BBiaHgnGCgZepr6bxKPcx6Wco6bvpDis5DL1B78xAFDLIDLxMlaJjEj4xPX5KJfDQkyb3VZUyGg1YzuT6uwS2lPwcZ3fuiK7gvH34AEHB0acCZ8mly5tzz7yKTsVRHJRucN4OoSQ8R6PC0C4uPaNsiovL59eAh9LedI8lnv91AAjk2Vt89o6Kq1Ccdz0q3mKJ15fGQfmCz/2Zxzf/+r/n+OIv+qvvdFL4KbFhf/nHPnp8y3/03x//zR//39OL/nEP6NP6ARLZyahUK27Xo+JznzVRY7uCB5nNzhR9oZJIBNxl0g4GLb/O2voyKG2ABbdxxgJr8U01QwfFVM2dZBx2w9RCwdHuUvMWO1oPHASkxl4lG3irr6lyG4pizVqSSZW8vnl+O1PXjxlB4nJSbuyHSCil/54G/UZNtyJVWA2kCJKrfp8UO7gDIDyLhVtodLDazo8ceTxTe+R1Q01RCLYrC/IMDvSSV16P03x2gkLfGxi2YW2jHUxf/0OQpoOyC6BCe+q+EXQGRfSLFDQZcl1wJU14LL2fh2qlouGflSJHdkohzz0B0FARezvWYsCzouoqHbiLyB0oAANDD7fgA3y1jconVVOgMuuGafSjEpLjxTpUfwmCCoyQqmgAOtN4/qsWeh+znUvYPgTGuvRQ7upmidp5HXjB/L2jXevcOsJ4dLzMrxlLGvVfZ2DTzwPvajXgtUTkjUnD9aQtgNYdJZMFzlPXFSefzPaLaTMnWGADVhXbwfJP8xhcl9lj9+/xPXlwU6KQKUSDn6BJcbYYTXdC1uq3+fdF9c3tGfWzeY2cMBM4Z16Wbz+BdyOKQTDOoLHKazjDSFqfjYDzHvFZuUUTlpbAVnOOM4uj5nAi6FaqxYaK50R5aNniNV0fiQXu5WVf3NDXZDQJk78u7oIEccS16Cu+2/Zm3ZzeNBCG3wXAQo9QSYjueBjkQz/nHaTz/pAfrUK7PFuul67DsRrppC+enRzex3JyadXbvaun5DQbmGTeSJLr9DGWRePPOt93NAzmjHxtnUdzidV2nBrM66JegqLf5+9X520njzZksFcjpoQi9A2Vwb571v77a11lvs9nv/hKP7/3f3twRRrpBPIccEI5UWMa9U1GTePTdAyCK4wGdnk7kO6gU694zESNk1VrZ8DggHbWqLIGdlGYjrguXZLrNMiI03Ltzpgchr3XmDLjlit+l/453TSud/1ofhb95OITzTtRdgc+ofNYHZEcIBf4oMB0l25Znq+7xppgn5zkoo3xtl5aaB4XgbjIlHAkfJRFiRIlV3vh/hzWuWLsc6Zv6RpeD7475s6M6PU6Qf+UI8TOL/MgZ+6EzeKzFuMP8JARyipvoz4R1iNY9oXOlysea90j6NPR4sxU1rk6sQM640C9CR7RMUggvDv+zF+Zae+1oJym/et1JDBVvSNev2Zjb2QyvLoFjbkUFXs1yDGg0j+l5klSadx8pgFB1qcnuBtOA6+Me6hQYoUtHb9FdDnYkQBzw1UOlHFpFYC3KDH0mE6AgGoFSLpMju1SZJHENdLdM+Ph9lZ19BXhrpK2rEggG1UKk8+nzyPkmNYTASlp0/ZSUZxjAPZ2LDo7ZQQBi1quJEHxuXG9Zx2CYyU/j7mwOXuVpqnsB5aPI7BK+616SpReB8eGe560DB3T1pqnYIW43/Fc9JRwibrKuLVnhdUG2Icj1jUaUTODp7LHWQaNZa5dNQIOz9bYOjMWpnJ0sHthBFTTb/DIFkyJ+bTJ2AEe60l8gEGFdqT1q8uUaXpf20zSKD/IAHLD7wkMHm3PekBKznjIQ2ZjeBxZejkCO1FRo8oCwgkT5xllvao3jen3TnngHkktoGKg0TtkBx2HlLths79UpYZYefLfCj6wdUrHGgMmB/kwtV+Ip7oEEcYEVtgA/XDSvSRG4K+JW0h5631HHwXvYd8T8lQ701mGy7Q8i9xuOtnOzDVd8PHd+d7rpefSxTONzHpA6uLS0a722jTf7SaWchx7lHY6cSl2f2fZssMLLnXuxYKU7SVZ/gu/5lveTkNeUfVPs++CUD/8Mz/j+De/4auPL/nr7++kqE09jo89e378q7/rjx3f/if+j3fOijvpRyR6b0dFZVQMwJQYaggIlBYKR0WkoOEiK7c1mHI6M3sChpwi/m2ohYCPQ+gUzmEqg6bqJlVjBNxscNZBXx1LjZGqJ1/VuObOUZFOgC5oWipolVaqVM2cRwc3HtJT78wMp6X7v/M2QgYBPGRjbmcn9OscreExRsROPt9CqWdrNJCVzJcGw8wg50iH4Z0L4w5GDaLNqcT7eQPA2PZzVm5yO6SUGbgBZfW+Gi2mDnuPSewdFQYQkFrbepJ0JXcGEUgdFNYFeCkDwvWClZ7ZM2GsaDtC+MqAtJNifBeVUq+dFbcrRwUNNkfOxV9uRCYF98Qb1KzRfSlUt9eXnddCoGCLfAy6dMTHXAMeDbg2kdfYKjgqqvH0HTra4hh1QKkptFlFVK64xpMKQD4zyivl5kzzvbSKVkpDwPnTuehs6+N2VOQgqm57RXhbYex7rf3Cf85NwTq/PPMb0nj/vFF9VPDyhaNiBn7nufvfUIjtqJ7w4hgTz0qBt33d+h7178e1bYZqNlqkXKISKEBCzva41z1fzvQxCJ7qt2RiTYDV5zXOn+lyvFdCpqKZxFvMr2s/VLJJjxkboa8F/PCm1Wstk7u806PIN9eqazoue8YWuMzblUBalZMJsMbNkKNJYHzc/BBZlnMcZE/JHrLxDGrHgt6hgvd5Xjgqcq+GpRHgfF8nBRl68sDBUaG1Lx5rHYRbMTvjroyTD+KoWPGi7hxZU9nb8Mz7PmGMtDR5Yl1cn3gCPO568n3lSMq5oUzL3K/orrfV73ZUeO+63nOSqe2MWv8dszlEN815EcAIjfz2Tkx24LTjgNVMu+sujqbswRhJmy2KfjnzdMJYzzdINp+7/Zhcjs+AtPU/Ayur916VU1ixu3LEtKfp3LoOfsg3gtsvs+78/O6MRFeJtsp+2AMPOx2DIBACtTNzZz7XCeBamW22lOmayZgPMvI59Fk7La6olfc3+08lc873SE4CzFezXQNkAsnWe1RZ0QZE4chSXw9mm/N8JaAvcAtfulSSnEIBigXNnwCr6eXUewtE06OyKe5JjGBMEQynkkRekmy03pfJdL12VNgpk7X3pb+kI0ChLBgf+lBE/7pYU0bOu1G6+Z7pgQ5F6W/KDo+RwMEjJxuzlTsv4LgDaH72/jOAt0+fPKlSPxn5z0hfrhPnZ/uE4LUcSlpIRNm/UH+AqB6gPhwu6esz4SwHOK2URRNy3b0F+lhJwrTZCFqX3cZodpZno85Guk361bVQj/Cu7tTjPf5caQPjWauzgXusR9Rx4ToBtKa+6LVzlL/1ODp0o1T0YwC7tgW7Uyn31sQqPWOpkqQOohKzKI1TtvpKN4CDIgLqokyq5oA+GgFu497KtLETMkolxwfOqttbAdAuzXUO5HqQ5arseFDQWQLW40G1fVrALZ110SPn1cs5Z0l7r0d0tc7aNUpjwZkZDgX2f4Fl4e1vm5/nSvTe6QL6teVaAPpQ2g7w13hufIBVRbP0CCQF3+DZs6wH9pXVQqZ5650eFs68vzNukQR7rb/S2UseikwtyC7RhW7NXk7ipx6jHRUeK/STySwkDXMwb9T33iPyHqRjOZ20jN7iGrPEOZvLM7sP59xl4CJzbRO0kQ27/X4FxO0P88lCqEu3SmCvIjHywL6fww66/LkP5x1lvpwlBhn4+jWwMDthR8rQOrtnrPUTZ79tmME7R8VqFT+J38U+fP5nf9bxzb/hq+Ck6ClFfm1s+o9/9Nnx/vOXx8/68Gctsy2CJn/kxz92/M5v+87j93379xwvHUnxSRz7T91HN0XV0YVOK3/98njzKhoI3R6vXz4/Xt0+O1z6Kc+MQD9ErCAljko30uSUQp0YzhIwqSgDK0vB322AZZoaGga1VR6eZUeFoj3FCFlHv5SWt3JUTExh56iA/ewyVhpTGhCIMJGhu2KUk6PCyp+VQ0fnrEAEChU2Kou/IxIMER6t98HsqLAh6DrslD59WRUBr2VGOmECiC1N/CKe6eTU0BxXgOLKUZEG9AAgcUCZUWFBgS+tvorJSy29j6PCBk80kotPpCbH1B41BWPrqOCA8HH0Be8lmBsKg9fCGRSx/nc5Kk5OCu0Fm9LPZUE055Mu40ij5qjAXjsD4gwsUhmnkRDr4rIBVUarHDPajIqckGFIFK6MnbERlUtI7GvfJ++Q8SudZmKtpUyMR3RUMroTdYjMSUN/w4za2+7jqOAe+/+ZUSLcIJ8kOFNEXPT68Toq+gzcl6HIcgUMaY3wn1Ej3Y5Fs4goHMvjBNDvcFR0Wp6oJ1dMHj/HhiXJ3McZgVk0PlFOPM9daz1ttenK8wiad93k2M6KitwZCTaNeKb6p/a6zquBONLkPBgB0Y7OVJaSeWOCxXKOEq+4Nl7yDXkIVtebTkW7bR2JA6zfkXxV19jYPM1rOrXzPyuqx8eC8swO4FUxprMZ4vrWyuiYnBVjqZ7FgOY5Xjoq6oz3J/UyXHdzlL2jonGFzoEIzLRvrpyJvuxtHRXnhoHUo+azNfPDmZ4vDaYNPazuwckRiDYEGvSzfgd9DWfy+ricnsQgAN60ci7c/9UV1dizI04A/Ik/MS9vBlgAgqoElMvILCvJTTrduBYFADl7K5mvLiyHhfu2rWdc4L8DKFjiQFJmKbd12keeaQBWTXQ/WY6KYZm7XhrAr5zwrnWOc7dJE3MpTgOxDBaK69mM9cTrNrzUjoq43jrnrPPUreKYcmyA7wqwtRPANFHqKwOEVh+CRqJviTOWD1lxMUdtO+qZQCTmDcBuX6qC56jRh+rshzMlfmJ2gRr8yn7JnggC/5jxzGhr944YbId5gpKzUdM9eg7E/Sg7FE1w46UTP4jnIpvjhnYkQCQ1eUamgPXa4ca1oyIeXk4Z8TFlpscwXRLY+oYzFxhNXuBeXNvlHf8u/ZoBWlw/1KSH+BTf6BJEjpBYi3gHS5EKRA07OzM2i+cbqGb2R8/ciP4Xr4+bJ0+SP87ZL87I4RoUvWQJZEVxGySlreEIeOqkzr5HqalwwjgzRUDqeJxiZdzk2TSt0lOgfcvtZG7qgyFO1LLSrvT9QfeQsdT7yEFeqcSvMyqQiaDsuV4ZwWWXLWds92BEV6Bn31eVJatybozy7x/bJvk9qmRF9QUCxvE7HRXFt8xTaKs+CgLDCkZ/jdiP954+JchMYtUiKuMozqf4KM6N+/DpzM2cBbqTmBVLl6mROTI6OBeUI4voe9N4nMbp/Pq5Br+d/YPG4b0H5uSU9VoN+x76v5yhdqSifFTYOio3xpJTdGqj5JMajLvE9M1j9s04Z6fpjQO2wbWjs1wl/EaBvRa++hbloNRzlLriG/A8n0usoQKAunPGe0OSa7qOt9RDJVFy5RSEhQSzkI3Rz6hl2RPvC157y543yrZPTEG8x3qNwfoTT9aG0rYofm28JhdkhXtsVuvybPf5e265VdVvcni0BDVE5z36kTArjDNi+T/2B1p9fHZwtuUj/8C69UL3LdtLVse7jIrLM3b68bN/xoeOf/mf/LuOj/ytP2/ppIh9/nM/8P8ev/nf+aPHD/ylHzv+pa//yPGVv/ivVUTC+Li4Nhwav/U//h+OP/wdfwrOio2++HaD/LS7WpR8z4yKj3xe61FR3grsAbz2lDeN+ckNO0XKSsKRFWWzYTVlAhOQ08HlZcgv6zNIvXqHe0F0JjgbnesIpwm4aZBSvPZuR4VS7NJM878jij1qHnLwcyOvNAofPgCDD+ZkBt9B4pnsMuKtpQ5CliAUxauriIbsPdDWVeWH2MSr+lR0YH7pqJDA2mVV7JwquQetaVWfU96XWsd5rz1nRtOUcDVZmKlDNb1HRoVpFu+G3kWhH+J+mEdbzxxVoz8rfBl5pJqE2bCwz8n9AzbMKOtGThuObT0BnTJedDBGo7aaw5cy0lPYxwjoBIdc+kl1bDtgtcuoGIfqchftlMmgZkzPbAxXynsZtIY6Sknx3M1ySnDXRnS+U/xFBLvauLeMzPUjzrZ8BzENOda4XkVmUr9Jf+/6QXRBNZzHNgc/nX1ngjfuHUCFeNWYAHZPlsOVs4Jgvso8uUY6SvTw/TxzuUI0q4eIopFjDOZjW5tVOaq3Ebk1B+1DGxOfU7zDJRTqfLD5Y0YaLUAN09XgQGiE4Sg6Ur9LTPWxTIsue6+Dfj0Sj0pwyZYZ4N+uTXPgkj/OGmvfjwaG36UkTcTv9XZPnNN4NiCx5zHSnM69wC3zT5ZbYbr6OnPDmTEOVNAoNnPZRnCd1mjFO/r+VcmQOpq2sjYTv8io4I6UsNAyNDzAZfE2z5ZhV7KxzqNpf0kvDe2eHYQrh+HMJz6IEXV1pj27LK1Slm1lFN6TKXzQsRkwvo9jaO+kI3Bw0j+7wqJ5zBkO1n8NnFqfdTkKg3lmusM87+GoKF1q75TMZ1+stdcJIAn0nlfHoyXY3R8y6h6QXLI/AKA4023Ww/wI2yrtkde+WwIE+ExjQwbFS5ZAQRQuSt6yOfvq46a3APhcqzxKfmDMa6fAnqW6OTHtAuov4xCv2LGBD4Ok7g2A7GU14t1lnnRQdaTxFW8ppw0iiiNDWkDkSrLUulU0rufW1xSNl1twlWvLB+0zG5n3u25+nCVk60fwnHSP1R65jFM0BnfPgZcv3Zx44ajQGWVpHJYlYkARgbdBLOTZXTsqAKZZ9ipThj0R3O+B+m+XbdIUKkMg6XTci8KFKSecpWDeEI2i7eCkE5JkH9dF6ae4H3XeFT0fbN/OMtoX7tck0F1As9/jbI8+x/gtelBEw2Xbq56/eddsx7oHQuyjA2DocFHvFGXYuOfAcAYiEAjr2+SkHBUEpkOHu8GvzsTtNAJbHhnO1hHqUdkzsQxo/qUBjM4K9fYQ8Ii5KuPPIHD8l1kz5diL71A5QfwlS/ds9aQ986WDkCW54u85S9/9T6xDxmTsACDNqGm0nQsqCRS/IVANvRcIyvM79jQ08JzAcRplFd3vDA8Hq86aVPw7ymajLxL0OlbUcFki05qznAzqskTa+Im7kUEm2cFeEqancIa0673OC3AZMlQqZmblmEzCMQv5UL1mYtgsV/dY/UDIW1wqa+uosHMAJdik8wKflJNzINi9rheXhZMJZ/s1ZUm8E2s24UKmz3AsxMe0kva9DDjIUYvK/HNyVEjPjGvpcFUWpZxgQTuUZ+QjphcG0gZvZTCz7ZpZd0kx72bXGk/SW9MDRko4hzLlpTtBiuwZZcIssKnO65KGXX3DtHGHcxE73PqKOYC4MqvGWVQZt7Gf3ny+95yBv2BdF+TzzlFx18ptfg8+91mf8fT4bd/49x1f8vO/8HjcmrP4ljiE3/8Df/n4dd/8bccP/fCPg8g/870nxzd+3Zcd/8BX/A1bZ8WzF7fHv/tt33n8J3/0T4Kp3GWHf8Ap/BS+zVzA3ksiJ2A+i4wKOypmQIjgTkWMQ+FT6acTCN2i432QnPobaawxIkRZtIyEGI/Bfiz2gPckbEdHgNLVWQuvmgReb9LoqJjgpIoubABQZ4IGemloMVLFf1NR4JBPNmoHlNDQjJE1znpg7c/WJ8A4iPRn1B598waCOv7rOqIcW0UypRDWoCmgmA2A2ooGSbohB68TnjJ4tv3d1XrOYAb+3RZ1F61Gnj6tvv4JBh/AqJjwvEdgzo6huYejAu9BrUTWY3WDuFkVWtFvnzs931RAHW0XvwPYdap3q0u9c/LEPStHBQ20ciZ1ujNQbKOulGr3IpDwNuoloTmDK+aLFvVu5t0N+5Oj4iQE6U1JATnISbjrsENpyGEiVH7ZnE21Lr0vTsEV4diYSiHcCKocGLUz6di5AG5WNHQXM185KnyefG9fKzgqJrq2srJ61x5IHZ/eHQGp7KWA6zMr/pi04w4mbTJYdjcNTUxHinQaZM0h0pvbLRwVme2UQxkpfzhnOq91aY1/Xu8y2C0IiqueeMcUFW2j3vtho7JHBlpmOEJo3COOixl/c2Nml7O2tt8dFeZMa+rqYObOwLdRsZpjnYkF/8Qr58PamfHUa2bFg9uw+5PM17c+nZ2dtUQW3U8meASNnfjQ0Fml0svARWkFGXraE0Yw3aMpXZMtBv7m/TbgY8fTCJK0CQ6yczPxqx4V0B14KkwDPfrMtHoXf5rB+Q4cre/lIuzoqsub+br5XXeN7T6/+6RQWrQyBh0EvM+DdM0HGWPpYHzItZG4liJ2IufZ7npUu2V0RpNuDDgCaESWgvYoG1FS1+v9I2qe60a1JKze/6IWcUmtBuguhOQAVknX3jrg83VzkMTozOlnd0WT5DXjiIchriaDC84/BKhy+zL6BUR06OME71a83cOnXs8ymTF/1313nfqZNHe6LiJ1lcHaeUqdVz6pnNj9KgKovYxS0IP7MrDnw2g79HElQLWQjzP/I9nYtlAJHjkrrvjGfO76v7Fu0dDWzYsBVLKslHsY+O8A1wLYorO66qrvyJKObdqiBchVWcHT/jgISNH8Dh9G+aYu2AbBN9pytkm8Hp5rZg742S4riVI82l/pvlhn87glvY58miA/yyzHmQs986xXMho8nos+YzePj4j4vo0qCQIz/c4uJzpAF+tOe4Bli+LMxLXIhlFU8KmXonRJOI0EWpqPGnxe0YczTuqs0baqHhWkkW5NP3rM79jYmyBolYseqSTWfHBUNGJwlpEYcPJc2CzeK+/a4Nxn2Sef8zivsMtUfoxO3NdY+1C70fcBpXAikj4aW4fzbeJndxom5D8xHGcA2NFCnkxb2WAx7Fzxc76bZykqMkRFgVgzZJOh181tNnz3GY1rw2ERJaCQNdEqVVjPZw8ZXufhx56APtWIvJ89Osmo10He6uyjxCycKgW6w7kT2Ijl4MTKY86gy9TNyTdJY3XxXbpA0IZ7TQa2AloL2YDeFDxfKOUjezycbZGpFWvn80uefmTj+Jnf4DpnUMS6KBOh6KfdcQdgiabgcjTFGrMMnJqOE4GvrFA9lk71yuBwNkva5cmYPA5B2y6JKUwonMyJb7jPCALUhLu9ImYXS5j9QI0JSvYlYNPEs+UdhhEbqvGkrlHDmpb27R0VdKDrBS2I1N91PjjIurYvOPurTe783TqdsupQhUNOo/lWuuinAJIsgXzxosVPK93jnaPi7dYwr/7MDz05vunrv/L4e3/pz99mUvyFv/gjx2/67X/o+N4/+0MmS3qJAAAgAElEQVSDch4Ojn/+13758dW/7BccN5uN/9izF8e3/t7vOL7t27/neP5inW7zAYf+aXCbucD9HRWj8SAgK3iiGiIZrJ2VtWqUO6W2qwFSjMDNpnj4yWRdLsfN28zcKgot1Zqlo2LFRDoD4t9qjmctpTSlFMpgVK0ngpV9M5VBIRtiPmRgqEbdQDTpqOiKBRWduAuphVN0l6OTzCtHh04XzFXXPeZohSbfDyO4K5IUMPWR0ez64EYQGtO9OgADnbSeDhY+2OMmSPuzVs6B7qg4pZ1aKHjdO3Ld1g/U2gCwUG4sbGEYIcprDdx0466Ptc8BjiIZ0mxUTlo3PVP2jk6b/iw611KjyJ9gHrZIrVmOMapBGTuKVnGIHh+nHGc3wnWYiTTKbvx7nR0VM/Y9aIrDeZiYXQJ7k6PCxZ+6wDcwB0PEjgopozAoEOXSS145Y4svx5K0aMwOYuvWqu07n+3Z33lPbn52VNDBQn7XAHb93R0VJ2dPrmHdB0XiRAPTc3NN+IDegDUVuxyN7+3vcBvF5SZm9s54jFh+IVmj1tMKZK2LaGBygiTt25mYD1pYZROtj+fNez/etwNa+/cwaGRIrRRMZOSJiKJG7xAVlZF1YwR/LQis8+y9WWt3p9U5Zoi1xpwey10g8t2kO0tBzoE8rZhngmKdyCVwOhhzGleXUQvntvlgrdUWTZRj3NmVdN462nWcJ2Wkm/oG3acMDtlGF+h5aaaz5TM5N9P02nB94n/cP6fDFu35bc1yfZJJ2fCgXlNngc8iGG0QRo6KAJKmZrWOTu0yZ3ZEzMb4J9pRUfy7Iqb7Ils/uZsmxbt83lTnu9vJ3VHRT9HdJ6revgInUja0Qc7r1M/cECRzz4l1R0V3PJxB9on3Nx0BY0fkovpRWNa1oA0Pp+Z55ajQmUg9YJxMP9c870qRXs25GegG7ym7rHGcS9HwJBHoz3HrPJimZ0fFrCOu9nMe3kwfOygBevFQG3+O2F5MHCA75WBGqKo0ySALzFYvS0jZ5uGy2fHQqHcYQHGeclTEeXP/hiphyAztB9BHzzxwpct6nZ2tk7Kh0Uo0RI3rGKE/ZTbrPTPg3SdgmQv4OSKfI5hHDoEATSM6P94fenhEKltvjhn0huWOyOXcqATir8zICQD0YWYQMOpZfUTacuD2h8zaIP6t/X/Duv/UbehARl+lJjssL/pa9kA580k70V+8jFJUN9A/AgwmT1CJpOPcJPrcX6mdGUUB99JPDOJy6Sr1AwwbspX5sigDXxW/reysEpedBuyoyKbacoLFmsan75Udb3Zk2B3j53WAnHK9ejuAbqZIbDuvnMnEvnd25ssBA0dKlcJiKRxnN50dFcgkySyacmZ1vpL8CaQlntn1Bjkq7DTxveiToKjxbm8jU0Cl+9icmeWxI8MlzpLLk3fZuYp74Ps4EPfWSTkl2ZA0q/cx2l7akGzE+Dfe+/KlGkEzayIykAh+c128J7cqMe1sAWdwENMxrXFkyGxRbwsbgwBMIXQHgZu9Pwzuu3ydS+Pw2cxIcZaHz6DPXTzSAZfxGxoVg7/wzOa+ply6EODKMoqzjWys4EWxHnJMOCsgxpRZUW9eg//G2rjZNvanNUzuGQx08lASOpPE+1nfSjcq4b4etDAL9ystnqw+Ia1EHH9j1Qjwpvj/2OdwKIg+sD0aW48l4gloELcI1RlR3guXW7eET9ltOz3o4KGCX1W+jMazHUuVUYhhFLkTS8kvmSjTbZIuA7wOg5zrYlB0ODsqcrkls7vuYV0hl6gP78JZQRbC1WO/EDkZN2QIfUTOdks3vHODle2o2brj/PtJ/3xX+umCIeinz3jvyfFbfsNXHb/si/8aRVSM98SB/sEf/tHjn/jX//PjL/zFHx2cFFQEjuPJzePj13/t33l83Vd9yTIbI657cfvq+Pf/y+86fs8f/BPHrZtP3T28nwZX6PTes/TTV37+i9OaoC57CiCxKNe7f/0GHnsozQ8fME3Okeeb1fUBcwpfCouoCwhPLA89G1iZWZEWuhLTH98BzC5Y4xp6/OPZ56h1PwNCW8IXQjVSAW9uhlqA/X12AJhhOm3SvDevzYVT9G1L2bOSsCPCPXi1M+PPRicUcKRfOn3d4DC94CFsXfIFjDoimlqE32lsGwM41xFAoRryudm6wZikwRFBHpTG/sJJk+tMnZKYufS0ZfSU9l8DXN1A5uNphHZjejbsLkFRLL8l82b3uuOmEUWfq8ENOzpSsbECirR4Ng8jnXHKjHx5uSg93ugCaacdGNuzui7YMG+VyeoOtNQBunNiKKAdT2Hxp/HTx+Rm6+2KublY+wlnUA0QKzqvw1y20Xvk++AqwNN8x2xkriNDF6U8lI3EKJUCYRKobsZjpvoqHdx0RAObhLAFYto13WkFHqha1HgO6kZ3xYaAro8E5rytlbHhHe3rbhhBObQxL7rHWWnrynUY172v7QC+LJwbNXZeWUpo8fu34ZG51lrPJd/wA3vkTL57YEJDJDpooEUQ0oG448fjqOd97zymgz873nMN4JHKDT752gSjcr7FexM0s1GiKLx5rfPEaSENFvFs6bz4txabOBitJMoG4lOhr48a8fmmTo+QYRw3eKUcfblm3XO3IhQ9K9YEpUVU2xpRyW4AiLULMIkPsKGJer1u8qcfqb/Ueg/AnTOZ8kTwgQQFyI95O+8P+mGzRhnrip6z4Ysx67u6Z+axHPPb6gudnvocdmdtfseOHvs4OC+ONxp9RkRgNZ4d31RcbD2Cuwy5Pp7uqJjX5focXc1+/A3TOtG96GflQLv/o/PK5U4PX868Z00bfiADBpgNGp+IyjewcT73GzqT4y3WOEudSgcrPaXkpA14lCyCIV/nYXCMNyfyCFRPIzsN61zmsBZQFw+8xtikgySGQz/uXJ5TcjudtGJdF167ACejeoD/G+cAgTKwQ84yQ9JPOBJtoG7X4Pw5yMMZZg0I7ufz6mw6Gj3OhWun+9k8N1Emi2CwZXF3oLo8GfnXmkYMBPp39yTEGVe0fvwGW7FXWGiPY48Qlh9xGRsDmxgXAjh4CHufqIhe55kn77l58ui4DWC7OdgAiGs340g4u9JA+0vpW6Rv61Y9Q6ZokvbVg8OOirQJQ09/GWWsVMJHmQrMCHGpw07b9R7Xzzfvgu0apVK0Zi715OVnw17JSJ8j9Vf0HqRTIKLKb+Pc0zYMmgwHEkH4XXkzar7M8FD5LNiK3DCD3qaNKx2X++VlrRJLCCrL40rblGNsDZObXB3sE9xXQCt6q0h2RpNk0h15Dz7pEKawx/+ptJPLNnksPhO4TQAjnhf9FSKDIvaynRmXjPvMz/jM4/1n7wMTiTJljWIae5IeoHf3uv8eJ+043mLnhVkRyza9hlwtnh58ViWjlNkEXi38gzy390iqscVfduxyXbQ+whAy0yKcUC0IBhUxnEGlnjboQRJVO6wryXnJdVQfjDLjqQs9jLWifR6OBJbLdgYH6Z/6l/Z7pzQoU9F0Zp0V9D5k0EjZU4ZWNkrHjUXX/ZSmHqYsNI+HjkFiR/F3jDsyVIhzRTk9OVLJbCVKGobRX+K/F/06433xvNvI9gDexjUCT6E39vQkWuZ2BOgKO0NhUypQIhY2q1WUjtuHDOzLus/EvqDfGuNK3dm9ZOkYSx1gJTtEiqAFOciqTwd1R+vw3gdid2VbYKzun9L08WEPF8EFK56Vz2lO+9U2cd5ZF19N2KljzZ8H7gHTOUJbi1lfpc0wytk6A+fnv3NULJd9/+VnfejJ8Rv/4S89ftVH/sbjyc1502Ltw0nxr/yu//r4n//Unx9L/7THxtn7GZ/x3vGP//2/+Pg1v+KLj6dI2RrfGxv3sWe3x3/6X/3J43f/ge8+3n/+YhVo8pYz+HS43CdfYlxG9q7001d+3tlRMbnJqz6dPLjR3IfRLAS/6ago4TquIhmpjU7Xrox7InWyR1u5SbGVDuJhVDBjVgFi2luMmBhlKQjHSHZN5eshDYQVI1d6dzzXqcpIFVftxjOnUWSUFD3osjYYOkPpoNzrilZ2Q6pe53FNaWsAbAVIIIoEYEg9iUKBERRUuCnwDSyytwbBYCvPbrJ8hntLsO5gORg+qaQwAoZRh5U2G0+B8tnMwSH6Tg/Pd4zIUQn35u2WTpG/pQ7glMvMKnEGhARwj45fNBfdCSR83xTetTTScCbgbeWowJVExPBcKso2tAhwMeL4NRSfcKChLMFpI9oX3VHhaIYdOxuEJNcohC6arXFweecAyvYBoN7kWnvJvX49OSpmJt4FtyLsUK7BdBVOzEFgyzLL4ZVR6S2yok3WoVRpPePKUTGeMfMsZynYoPSAO4DhckAEHv1eQAzanj38M9GM+B04d3+WnUnlnjg5Ks7Reh7r+vQOWzkM1GeFK1rgcINtyJjHYKoJODXP7kenO2O4UGoudqG0aUFPqvgwK+3z6ohe8RVQr4ygMpj7kx+gvFk5Kmw4jY788zHrkemr3W/rGsbGok4vT+Gacmx0J43b9mrAWr/V7kQY5g/Nb3TSV8aD9reviZVn/xfr1hzSS/qTo4IO2rkAnx0VOgNJU1x/2vE6W3YkLDYYxlinjs4SBVwwWtrZJryA+kjpLJyral3XxL1Imc5veqw96BlJ5Bt5qsHibXSQd7mnT61jd2iQhxSQ7Oy9M4VdfnPBZ5Mr6JrSIXZSfnzTFeg/OHAUBOESIhs7d2Fiv+Vc2+XWMecn7Ma8wVxPtoafl3jJift98DGfxqoGl4MxM7CB1T6d+USCRc4Yzj5Eq5JrOcPNRKpxpIMtCJJOvWQaqB66N4BHRRxWAEY53IUtH69HMT4E6hboNdHhdsn7WtRaDc9Z6ZhN6+G1k0bcz9SGcFgChiV1CiTc8HByIearNoDQvGP23ybgpibUpV9Q0u5ouZ8Jn0/2g2DkbTwH9kDYRGGTqXFrAoQCMh2otTpbfgeaW78iqB2layOgLbIq4pl8H3t7ZZGktjSWdSwv3DLdW0YFViwjY2mTaRllCx4AcB9GQ1hkSwwvwKW08XgbbMmwY1Ee50XWrIcuLGfK2VGu2vFCRGNNXVrHdfSZVeIAGNupzLI7fyzvWqZ2ZlwF6Msxx5rE1MPhEPY3dRdRSzoqbEOwoE4F0TAavGrKP4BNEXuzExXuGYL1ev0GNiWAXL005u3SaM+fP1+WuI3RQc6lvLVC7BJnDEignh7AqXs9jI5InkSWpqJ8Nc3zOeFkQjZI2FJHAboIQMzAm1l/Lf2KtF5O6DS0MsCAP8b+BU3HOY+MnSc3T6pU1quXx9MnT7MvpWCXLp1Ic8pqEPkwqwDOBQP8lW1OIHQM1rAtDV7z8DFoF5lC1oN0vUtu+RzDVh/or84GsxseH1Fyi3tNZxv0I9sATX74DNpR4ixl4BwPwhl5K6fRY8UWEg/oPXisb7npfKwvMpNe3Apvar0ORez4D7Z/zVNzrt1BEmvrc0KChLZt3AmZOqhOQbvTZ3nkp+NaIdvh5jH27vmL57w/8K8A/8H7mVmGTJS9Cr+WYD2rUSTp4BY7PuCoQBb53rbrZU+zfSEC4DigLC/mXjZTNp0HF2/YOSoc4JplWkUjFQjrYGMGMcCWmtdDerfLcNlmp+P8JZbPspR7RjmVVV60wLkWD+9e8JM+qEFR6pcnbfkk9StNh7LsGmBuQw/H2t7uqOg68kwAM863dFZs9J5+7YN3GRXrVQph996Tm+Nf+Ee/HP0lVj0pghZ++Ef+yvENv/X3H9/7f/7Q1kmRB+QBPaz/7Nf+HcisePKYTG/+RDbF7/mD3338B7//jx8vIur4Si/cbPKn19elvDESUYrwpkfFlaMCCqgUA0b1UmDH2SwFgwofBMDyoLphZGv407yk9tKXJ9MpjamFyZNPYCGcEPAwy8MPhpyX0uvveuOOKFl5nF3blxEcNJ5cY3ZLD0q7tpIxGMaOwtHN0AmghLk3h6NzpsDSfNlkrbVB7GoEs0dAGSoQkHBURKomhcMAxkjZQsSHoqe2zpl2EHcQhssiBRDEQDOmkIfgohHUmLUPrx5mwTIApv3wT5vQx5BnfM72yH4KirDKPSGBdME+e61XzqAazj1AnHbJ/B69fBqDnHeQiwTMXIeXaet8YAA9VI6pjI4fgW7xpRT+HiIcAOvqQ3C2RRfK448alQMD7cCbtUQ9UdoP0ueHD5kDozkETt4DOHN9XJQ9U91i1sNdNcFsTcSnMmDUe7Tfeq9XzZFT43htofRv/U6qLj7v5/t6ZsfZUXEf+jFlkj77h7udilP8VYT/8TsqpheC3hp5Jdza1tA/2/HZx5uUsgJ0Jt6Ys/T3+aBzj4i+hqZNRz2S89Ua+d8zzV+dXunJovvzlQGiGZAv8Gae+fzGsxJiw6zLTZLqm4/fUWFHVvbNqb2c3YmWWZC3MkJOPIJENwAhJD+mOmMdmmHM+xeK18DcVQs9rySQVGIhKQ5PGxwVQ8m5JUvjl5NsCTlE4C0c9G4MaX0k+Na1o8IgCw1ZlTSZjJloNpw0miCKjB0ti4FPggw1FgZtsKyCG8+ixnPjaRm8sZj2Vtfd8Nsu864MposV5k5fKNkFhjKaLvQM6AQRmTrIyC3ecPn6u4y5u8bef9+Vf9qJq/tmUr3NGE6cQ2s0rHEerR0nW/EbyneXvsPzMuhnZyRtvlcTYpx5A8fSpxBZi0wLRS+rVIczpR0shJrkqGteDX6lugK47v2ZcJQ1FIAkK9p/y0WmLaPPHY6KenS9edA/N+/OLFAEcVWQxprOZEs1kESHazAQLP9j/LSMWilD1YLfomEA49X7ROWCqJ8TFET0v1C8Xrse2fICmZ2l28s0kdcmodL5IMCfMoKAEhrBqll3lJqJ0T997z0E30A0pKnKPzJyVmBuZdmklTM4KizLMntDUcwA4bD8XXBwvKy7H/2SKMdYoobGWujZATiFM4CZvR1Yq7KKcQ7QH1PRyJBjCNQrZ4x1TfA92c1jv8GSGlz7wDeqWW38GmAo+gxgr+K/MSb2e2TlnVavPr0WLboYoF70oVANfpUoQR/E4ziePbtyMPD53RkCeQU7hLa87essKbQ9p+W0oXNSto8yhUlOBNJZVWHtqOB8x6xx6yIuDfX0vaeYM3vkua8fB5Z2wMPR4QKgFRCG7KnGBsmH/UXYtxHk9+aIrA3Yu49vAPoCYM8MhtRKJzxK5XuagPGer+Sae1RkkAi9FgLZ+Q5kBMBx4ubNPEd0Sphrqb+LdJWaHv9KOnLWidaYpdLkNPTeAuzmu6KSgrNS+JzKsM9+Gq9eA49wpjz2WjKA56/KhpsnwT2S9sjohH394LpPmWmx6zfB4ixPzdfg0ArAv++FSpcVv/b6cPIBkKP/pypTVPkyrgn3gvwWJbdevkx+1emPa7D+gNqafkX5aiuR++/92umGLoVW/K+1LE9MT3gcF2Sp0/U1XGVUxKhQ/WF2fsjpkbaGAxiU5dFnThiBJbpjKA5siGuQXYMer8b7mNHVS3CZfvOZ28oC7a1dzVnJ383eeA8pF3T+4FVXWdvNfXc5Kj5enbbsUg7gnaNisRGxT3Eov+HXfOnxtb/8bzree0oh2D+xp//fj33s+Kbf8YeP7/7eP5/1QC/oIX96+uTx8Y/8ir/l+HW/+pfAGbJzVvy+b/+e47f/3u84Pvr+85/mzorU/lQy4YM5KtzUt/Xqk9Bi/U+WViK7pbAt0GHeeyhXaiptBSfrempD3dAL3nkpbGAFMrb8TDNx1BNUg6bCXZmqSqB0LA8z0xrMpWxyXRjg0giPSI2Yq5t8ZlSEDSytQ3tJiIaurKYyQET/TPpYh7X42jsquOYGwfjQbN0DLa2XzsoyTy0TYtcIrRj/2m+PxljKiDGAboGVjHcyRnaRryIi/ue0Uee1zQZcCwaSyqjrnjpq7eNwVPTXXDk0xgnIxdcZVgdqEG0swSJg0JEZTAMnLaOpl3qKnHmfFOt4DA9LU7Y35REyi7aAi7gdTpLT6k80OWVUQGlaOSowHlkJ93BSmIewZ02kejLLw4b5af0H4HJFHzoJerfBjrXToxsi3g/XzL2WUAbsOd0d+CMD6EzYfLgUnn53kYMUVKe1UovVKTHvNRHt3r/mKbh6+qmv5GlVmx9j5ajw4/KRnc91Y0DDPc+XkWTrPfI+BPBWBqUV7HGszcFDwhqOZZqQbXwEIPM09m2haq3+IWW4a5a5F51O9JzFsheNjOf0fO5EGptwLIy2EIThzFuB5iT0HEdN6b4yIC4gLoFN3FeVDZAztKIUe2+eBf2hIYPOVMsawZUA5JsBNjLPhaOijP/p0uGQdhnTHRV0AJCfFWBfm1RbWe5gGstFTwRFCgiK33aOilyN9AkHPydfefmKjRpdf34F9KQxiizBHR9an/k1tNuBmAK4rjhc52lrx8Z1JDf0DWVwoqFul38NjL7msubJ/UBNtGCecsGDV+94W0cFQOLFUb/P+O97TRexnV/U/TNj2csde9hBty5PgRrW63IvW27gKH4tO4EmAU55PhovEIjJ0hTMas7giyzBonPYwi8au/jAjopZ3bgkiXaerZOPculCdi421M1iHR1q8bNzVODpm8M9SCOiuwSnk7E7k7Mx+sWYDOzi/GXDT5atCD7hBtXU52/Art1gt0rnqk59Dwxqme7xWtbpp4PCzjGWn1WzYTXlRRQ/ei/40EpGxfzk7Ajbzu9G0JXANQbeWfZVlj6i/dXsFnbow4Ml/hpoBbngaknhTEPzWwK4KON0+wKgc9ifKGMVjoosM8U1Ties6Caui/+r0iR2ImBluWcRSY7sWI5r/ISeyw+ziA1kc0yPHj1QdjyrFkS2Mc6ewTVX9GlA4yyjgnS873Hbixd0TqC8js7lijdBD1Plgdwq12VX5YEut3Z2EVVW9y6UDGr9INC4HqW4eNZYSorZG/44WNIltUzTPuvMnOB7GITHQC+sU1PtkuYCNwBoT1uDEeGVaXrmGTp1ARoLkMbahUPk8DtpsznjIR7fA8v8TDabVnNiZU1D1lvHkn7R15xEotpZjUEhmCPLBld/yHJa1CLScVx8f9a/HRXv/qGD/iInBPiZ9Dhke2h9nQH6Oso+yel8Ak97mT8D1whoLCe1g0oiKL5nwiQhxLnNTP6Jaq2Sq6RWBkJKDa4MJ96Xv4v/usScfzVXqn1gVlIfC+hVfXRf3TLK3z1ZWVKKNMHtE+/SA9aSRWelTY3rSPpm/001KVffjtXZtaMi7nL2SGZViJToJHqNMnw+K5c2LA7Y+W0OYAYv7WUJm5znK/1/4zMyIAEVHVqPmzdv6EhSXxGfrdqfGszg2NmUfjqN3LdPhz33arWwIBxSDmSOtSDZrb2s5XB7y1YxljcvpWVb0tucKb4bT+OvyS/fZVScV+vpzePjn/maX3L8Y7/yF217UvzIX3n/+M2/448c3/k933dnJsVqP6KpdpSB+vqv/kVH9MBYfaIuaJSB+vf+i+86fvyjzy+29dP9Jx0BMQoySDG7ECSR1vfq9nj98vnx6vbZscuooAAPA0dYj4z2MLZD2SSDphbQa5jOqwsP6Csqfq4/2VN2rZC4kVEopmHA93Qy1+GzEwNwQ6adh7LJ9EkIDtXitSjit2exYEdF/Jo9AaDkLiK4DfRI6QvGaNBhMCjEyMCY4cY3OMA68+5r4RIx81rtUvl2FBsZFY7GLwZL44PMu6JPXCOVnmsald2RsgXgNz0q7HDClNGAi5712D9mcoxgnJ8/vGfelgnQlF0s2dQAR6f0LBYG97R3U7h+8B4VKTiGJuV38JA2r3UUv6NKpMDY6IPip7UTzbqGLBTcXtu30TX2mhMvvVzPWo30ZATbkGjnxKBej+Abak9dZVTgAJD+Unjqj4Wug1+omPIiNKkLehpSzUUGjPVr0WRebP/XRkWVdpmjbOY1metmF7+w9tuMDkQYSUfHz+SB6YjcxsosdiIBcL+nVifeYYBjOEswnrkGjd1chCfvwJYCXec9amp8Dhrgp0F/zTtX3GdDV+cbFw4K8wvsdVcSTfcbx5bXIMHjRS1XEhLnNTh3p2dy+LW3tTO1rgkGhGGU2+Nay+47MDUwb6t12p9uMacTXXSz6XnRDd1OPTNobM7YIPbBqLDDj+nSvVbwzlwCU89SAWX0OTJPTUhbX56zwzL2ossZvstAih0VNYJeQ5mAFxxX6lfh6FWPpW/pEHHWtjbqREcQjXtUMNuyg/Q+u51wm6OrOSpMWySdMj77vA2odHrqho9rZpvfzPuYDqQWSMA63juuudm/C+dwgUaTU3slKNp3WyBqNvTav1333mUy51lg9PdwLszv9np0R/GZp+/W7I6JdifgfGkLJkmZe2aed7/g4opkBWlIz/jAvOcX82xAvOspX2cNr5+FCFJFKGMvcC4oguy8tc5Hg5sR3NWjgiAZy3yMvIPwxQjqWf7wdK5F264nU+dVd5JXd1QsLxbP8n6JVndnIcodIWNB2cQzUDpuu92JtlBqXw3SAaBXWZy4N/R9l9omb2R2isGxFVmhlJL1c3ljg6cAsEYvCJb7zDPlrIOpT046t2wP9H5QqtdtUAljFUhn8Mp6edo+U7yWAf+4F6VnkPnAcioV0N5q1lv/UbkVgNQ34VxgBDKAaC2p+TKku+rsB7AY98SYGYSmOvpuOCznC/d6tPKQMR578ygy4lhSKZ4V4BXA1oiklu1nh0A849wPwjoc5YlLuyDLHdnUEaXfrsEwlJWkveR55M4bJIcTZtL/nb0X44nSUe8/e4Z7yl4eqYdgP/X3OMtBQ1FWCz1XHkfT7YoivsqoII+I/6euBHpuWVXWce3UNkawclTUEXVQC/U190rwnF9ludzWeLm7+KLp9Ws1iHb2AYL6plJ2KUcJ6ro8U4wR5bgATCuKIPoLqrwWbOMsozvyNpZZIl6xigy3DtCzVbC+KmdkwD3GGs44OmdiLOxdAQeKqiWkfe8sp6kc2kkem9YCCDkAACAASURBVKeoj0ngMNhnz7HxCTfTds8MjBsOSK255EPnlQ5ktCrMrA9WnMC66BzFXO3cM8WbOl/FHDZqT/LN7ojAA1pzZzcB13lhGSEGlTKzRo4kvbCrJ9FzKwIHM5MCfmZn205OCa0bMgJEuIQitOobHY0OZE1R+md3iCI7JfpUqFSYcbN+epeOiqCfZnNZD4dDWJlWJz3Tk48zSyE9fNjvypmDChJWthWdwlWWFe/DQ8bNi68ow+iosH0HOlbQMvh0K7WOnp3oZzQ+i+f/HnqfLukyb6hEYUaz2CO/ETiag2GVBX2no0JlxxxdzO0Yx7vTK2dbYZb1/TnvMiqm1QknxT/1q/7249d+1Zdssx2QSfGtf+T47u/9fjQZ+6CfyNT4lV/6C45/7uu+DM6K1TmPBtt/7H/6M8dv+Q//u5/GzgqfQgnID+iokPaaCpcVohCKqEnpzAUpiHtlhaCOBToVIyrXrHHpzAYpe4ocWTkqLHPAR8TwDWChGZpKU1gwlVHVQRDKLckATNMRDhGJYAfETKeI2lBfCETvRDZB1ovl1VBpwdTJzqzco/yT0iQt0A1w1p0FD973jEAxevRIzfoq0qhjYnBkAPTEqiGaM5RVp+SHUsuGf5tGQAIl5zHZOeXofyuaaPoW/6cG6amctAekgJkVjguApYOfQ9T1CuhQA6e4B2LfURMTED8w9zvAHdLevjRNAdWaqI2HKYzKYGLUpU8QS2vsZ6DpK1LQme799OmT4/bV7SKgocC/2VFxGs+0gYMylHVcO2xII8Ayu24vw20JTqZ1GMqhjCzdTM5kRU1AppeLViRT8eEwpEHjKFxvT4KBOYHWByMjDsso6o6W3RbPwGF3BHjICQLLUTGvB9d77NNzJwaX9KSVsTIo/pQlA1ozTqZaa5/CuHKJgy3TWGv1Boj6DvX18V05h57t0ABq0odB5XG/52wGMknXGqbx2nThNGTnqcS5s/MKfBXOb0azZaNSkSWVP5UlMCO8clSIJLPmacuugOgMMn4YZcxUp13LD3tn0aAtBUFO4tzPgvJHzmTJ5/X5Wm+qmx8OinZGOVMSdScH1st1dIfItmWQFF+qXkN8mqJDs/ST9u0T4qho9JlEt3ZUWG6UE5VDda1cr5a32yUvQu90oACaO/cMpeYgNf468kbSt4MMzP0MiPGdZ7AxAwig+1REaVyJEjjNGVEACftT4DdH/Hag7kQOG4t987V54V2yYUV1O3DW+lutfYE3vUEvnBXtwTnESybJnRgcEq2GM9nJdrKXWW5bdnnhqPj/2XsToN2yqzrs/uN7PWhqSa0WAglNRsgSKAQLTHCIMQiEMcSOje3EFSBgF+CpIBTYgDEgE4PLxiRgbDwV5UocQgiJwWDjgKscY5IIAwbEoIFopLulllpCre73/jm191pr733OPef7v//RErS6P5Wq3/8N9557zj777L3WHlCKRi8E8az3+6YrX/5Zw1nqZo0vO3retXNenWCV6JCNnlRcBxyEMlbNFLAElxEVIiQzShVOvKLsXZ6ZXRGRgwVoR5yFiHNoHFkfPsIR9sA39QT6r4Bo7UsG2MYutRh/3as5fOIeaykNO4282qwWtYgKB2V8z0NPjmWUfQRi4xTZILCrfRqACKp8e9+bXX9+Zp425GsrYzojDNyy57YSNXY9A91snpGxsLMcHFjJ2Av0mCjAkHRfE1wVwTQUf5awc3utlH4SaKosd/Xw8PmMxqtcKQN6DfhyvxLRy6YzUAoI0duSaew77AMnR84MQEfZoJOTU89y291HfX0Dx+z8CoDJfTzcQ3OjZuMWwWtj9rny6Pm+SgD9Om9mfLocXr++nJwc+7UMvBcpZNc9t2h73lR9FfcO9pN5Kxv97BRjQhNe2LOeebJnthLKPiHb49wDBM9O0S8BRBb6Vzhw7TXdLYhuPysY+HpaCUQQaMoesPm9fv26kyN5hqVuUZNhDzyjvIhUQK156WY2FB7ocWEGvh/0fbfr0b9GiKyD+pblUMHHxiyANpDNJFnUGQtg+8z3nJUWE6GATOpiW0td75t/hfr3IFShyNXDw/2PsFNx4qvci/m3Ji9mR+wf7C1nJ2dOikFm2PvFsw3yARpbjESF3U9gJ6pNAKzVuR86g02i7e84TwWOszSw3RvlcjGnAuydQCMI7PMXFW3rKUZ7mZlvWCeW3OUesbdUatszYAjoi7Ax8N4zJw/2vDeN/d6wHdk43o80MpQElMBuQ2UMI8FOlz3qMyjrHGMN4PSMCh0I3fGlPV3fhu7G/z1uxucT8ug9eQ4OfK/Yetpzefk3f4bUS7LvJMeZQcIsGvZptesYYRS/JdCOQGGeb87Te/rO0Bi4cLuPHmjX38X0g821jVFyguVqD0gQFUmguSw7EZc6D/gD5Nyaw0sHQs82JQsQAMk5bAatAN5i3yLASP5p8hLx/L0vVg5wP7tJNIN0NnIXDcNNH0W5ciPaT46DvJP+gooZGQtFxcW6tt/LMXO3dkRvfW6QCReuix3bZCWIy4iKBj/qGmxXLKr367aJfXyCqBhup2WxLAcjKP7sF3zqsHG2/eyhR46Wv/6Pf2L5sX/3q1cq9zS55WJloKy8lJWBuvP2a23UJH9kPSt++N/88vJd3/9vvdxURO/PLvph9z434JYZFZ/5jEH2iWv0uQOohsk2daop2SiowZzWyB772P72en9t6IT/0iAoRICgxrR5hP79GqUfylEp5MnV5kGFz7z+Mw8/NwjI/rvRoegXY/W910IyxGj2CkMF0Q/lwSKqTDX6kDVRQQA7i5DaimgffzZGGqUDbu/iwrOSDXAwk723f2caLCNpvCEXiBYngbyxVYn4ILstUkJstwx9BEwjetONPpbF8mcuDy4XUoZnv9SRqaISLfZ7As/5/HCUPEW1pFS39+mu3IwhPxvJT0bdToyBqOW+vo4OrDgsKHNIL0ZE8WWv6pi6PBCY6sdqBqY5RyZ3Jh/o9TImrMAzJUjdQcKrSAW3K7aJLmhP4MGjZfQkJJW1qAkIr9kTzrkLbD//NioaUP4RyIi6CvV6+HkF5uWs1prYmUViXzejy3u1MMIIzoNFDsIYtr3h9YAV+WHz7fmxxXBBxzYMS151M0/tkPWX7XVsl5JRROMr5YnPzej2dsI1dyKZOa5mHtfAt12jzb7QVet310sLHRD+4vCh2mMgx1fXTdFycVf+KHRpvTWzSEbPnZKQhGDYvFyeHA9G3o5PGQ99skaWyUCdaDnZXGIdmX6mYOlTD3AtmgEz8k7ysTLMM/KzguoJuObsBWAdzhe9qc7/8F9ERFJXgqZf2m7fwfUo5J2iR0nojPQZ7Ka5DbD5s3JFbasQnbEDf5lOrTpCuk8OVerbdrxT/UcHXPu0BlEItND94GDNeuVgLwf3isOSoMzYYUp5GDVc3zTf284Qyl0IWKny1+jZTp63vXp+TyAs9dmqomX3LNMGmOM7yyKKT6mH5SQ6oFnKoPj3rjh9aLKerxkAffW5yV9UB7JVg3xCggzCGnT0KOp4XRloffKPxid7d/UZ0AoCu3vRNBh2n2S2hXqmZFBHGq3upYwANny1vZUZTgIG2XB7BtyMiKw5zkOgDiPR2Ya/eDZkqER8Xs/B+rtLAw36B44gBtxZvXEMJBZYBfB2UP71srn0e2UN+P7UxlgrqYczRg108TnWV+BWzR6HTzGQJE6Cypp4poM3ci3NrHsjgkSLro+zC7f38aihdq3McylhmWPH+DP6HXXjzX9DE2DPkOcZrybSAPIha6gUgEhomwwDV9UYurE/GVm+v2skjwV0wQfVTArwtHeQzQDQSsB0BFTJ3+C5K99LAQUaCxr7luaxDmCzrBHLQpm/bfYrSBX0CLD/eSaHkzscn9u5Ku9kIH7RSY0i0h/deR/HVxv04P0Y7N7uL8NPt3vbe07YsP+hXVXAurIjpaDTDsKeNMDPZMR8cWT+qxwN7DD5zPase064IFvGGkCb3jKySIEI8PURyOL6xvED2GMaD45sZZai0gHODvgI9v+Dg8Pod+nzTAC50Q8l+r4/elAahr6AppiR66ZnDw8OnCxRaTzv4cOMebc5FKzV9Q9wP7QSieyJ4PLNfobWY+X0vK1sEJlNNXu+7snJIZdxOx14XQh9B5i5f4Wt2P2MFJVf63JjPQdKxQr72wk41vy3jAovAb67s1jGk+kJNbv2deQzLnvAXGx9PTCSv1fmiT2K3c/JDzaDt/dEDCGzVs3lkbnlWS7eTwYkuz8Ty7pBttmjJrZL0k82FicD9/a5D0Hm1LJGXlrPM9hAkhkJOXpNg5+KOYmxKZtxbGeqX4gIN7ubA/0bgjtcp7PfiZMuJLJFckuP+9wz4234DJ6plsSCsgx9P7ouVaAy8KbExAqRwpJ8jkVRKdf+eGvcgaf8pJSigoX8uVhmj6DgeB02BKx0hkXIvuTK/QpmBaEc4jhAf2ZXzWxG9YNRtZvU3G0J1icyKjgzZgh84ef+nuXL/9h/stw26Ulx8/hk+Zrv/BEv92TkwaP1MkH7g5/6scs3fOmrnLgY1e83ofyJ175h+fq/82PL8bEdfhtYtkdrYL9jrvPBJSoEvOpxFS2zaY4d9HYDvaSK94Bs0dsexUqDet8iSqwcVEQrs260DOhAqvo1ruWH5BTCxHRDwCJn9i0ah2WB3JnKOtZp9JsRwxq/9WwhURE1CT0SUkSEkQWIDkKmARq4+WFBb6AqKdn5M6JCzoX8GxkqiKxVkzc4RgBfMsXZ/o0oTR1C1rgtWX9EvqH5tqIbUlH6KgyJihT3DhzqDpY2daXU1RXorp8L3Jzto0pUbAC/4udlWH5slN8LfAr7kQhH/x0ZmvpejdydOu+dIRBEhZy10KEwBKKkggPX61TA6kY0U0NQLKMpunV4VImKFUoc6dvr5SpETk9URFgGrpdxkyTDRiVweoBLVa4ClVqDkzIyHXhhpoPuhxRpvu+Nu5nC/igQFeGNR1miksnlT5wAuYzNJhpmqstSUisRinfTMcWfLZHRAvn9as3OxZzTIVExMXablZB89vihlFjdz/HDoBinhN2YqFg/RwIzOgcA0OzuJ/HmexiigNVxp18+KwaFc627PuVUUlxnVdFsXArqHTWmrpHKdbbGhqzG1T4zx7oJle2JCju/XN9yz8U5PCde0w2rT6eSRyl3M3Wdequdu5aYvOzX7ecBAAWxn1qk7oXZveN9lu7wwAf2UXA9UbMKKacCfOf6XmUW6xkz792wfuI6P2Pn9UqzpEjzi+qUlgYzRWdARrNperPSkwaLkj7YCOvMtRlpNIt0m5nmQyqO4KSNAYBH1wTyitM3cggr6HKleZ98+TKiotEdihqvz1H0k2R828ccaXfgcegdEplZpdzN8DFmN5wsXjjmbMTqIJmDQAAhnRhkVhkAj3lg1Gz+puEikyNtrM/Wqj11x4igpvTPjk3atMFb04nJOt7lbOnnbgsfNQnnVif72VWBLEwujy18UJ9f342StwLhCjitfZ46k8FRjCS190X0NbqxnC06X0PP0PeyscEGZ0CAg6cYJTR6syswdq8RopKLICr8OgQJTYT8rHYQVx4V3pOOQ/YATvhwP0w2zW+ST1Tm0cfYnf+aO6MPVN5KJIf7dqUeOR6G/UD8fCn+rxrLs9qAMu5rGa/dPQNUs1SaTwNLoJivCpA2a+djnmD/eb8LA0tZ/tdlsrFbOMcrArlxcrvVAMlkIK+IEQXyaJ8aUeFNhMN4wYr2NgyOV5ZHZlkpJ1yYzSJbzDP3GbEMPw5llxqAs7HdU3Y8sIz6Rj6zAs6wNVVaDcCifd+D55SxwGdwcvVUAVbCEmq517XWjHJJnV9ra3bzyIJDbWx7voaWPeMBhKX3R9j5InJ2dvx7Rnqq/LY/EzNznRCgjs21gJ9vcu/APGVHgRe5SzacdJwDBYXEBi2+ak9UaN5xTiMjSGP18ZyfOUEBwFpZ1SgT5AC79a0gbuGZTcQ1vESUX5T6o6TLgahE8KvKHKJJ/V5kPvu4PHMEuks9daInopdMs6BBrIltLsvQQVNs1UBPZRswRGcroX8H5tQba++iVJNALQum+5AQFSSFPSNBaz8jxD1LHTLuxIKCg9msXVlGQTjzLB9JjjK/RLjFmV8yz0AiUj4teJcYjf3G702bRDozMRwGGk/8n032lhGhro2iXFWS9v1zzI/4tu9N/Z2IHpx7uILJ/xnLzG3YZVt9lFglyt3JV/X/FgLwCaKCtZ+/4FWvWL7qT/1nQ5LCZvzo5HT59u/718sP/etf3CqTAml7pkiRwnbZyxTW53/ay5a/+Cf/0+XpT71j+HWTk5987RuWb/++n1zuf89Dl13yw+hzoS6KyoXxhnS9dY+Kq2ZUePRsAZl0uK4BNEwpHCM0Gap1cuG8cKwtwoWDhOVE9nZQT9XS3RLI9dAcGmU9GJhLGcx42BiZ/uapwpa6pRJSdTwFBC0mb5vC3REVmAc2lfPoGqQi49lF1OFqtXSRHh1w2MwjxAEuhW8K6/DaNTRaZikJj0IRgMOsEUU6K71VyxYNx2mt+6Htacds1uSGviKW0OBYrwCXsbCrfeNPWEikMEgZ9Y3SWoiecVLF5oqX2eiAj4iKfgiBMgoEpwzKWOR/RVRU0KwHouoz6CHXJUbGI+4JD5Uxqky8IoUiGkwH/9TRLlMdxi/SNyMMvHzF5emKGRVTcEjXDctsk7pkRpJ9ZUBUwD3N2pWQLYJ8fv3eTSWRGN5//7jrNfBazkrf9ugG1B/1Jo0WjXZyjEgulz1G5T8KRIXLMsmRrLEPMqQBu/teIrG5qjYYzXGbsVU0bAAVI4dwvlozc6zs914382I90QplX/VE6rP2El00aUNYtERFq3O0l/NdWv6pmzpRCDAi9r1F7zHluUR5BlFBx1nOvoMAG4iKOv91iyh7AUC4ARUZ2dr2eblsvecg9iZSu9930AMiYWot5nlT5XHbjAIMj78wFLWeYJDszJyKmbzWyKqY70aE1xDXNtequt7Xu+qaIXhWr2pERZ4zOu/muONsz43P002advhZlMRRaRDo43Y8mKdch/ZKl6+PALwPPVERYCZrgLeA2JVni4Er+btNAQhXlddNo5nZGx6l3evcCgrpfGzQ8PGdhpLGzAlFWuo7ZpdlGZjuejPD7DKigpdBdiPsf/QxgD1s76uB8pxIGO+XjbbiaDqUYd5/tsHemo1ptrd7+ZDvI9zCfaR6Ts4vNNGjJv1ozNyfPe2lSm+wOGLaB80STQJm9RvYY9AZ9TeI8raX9yggoCTAV6iJQEv9Fs+cPpr8RBy1bQ3z8Zqi1Is/N4kKN3mtdIkaVe9YhQfLWLcSJixNUzK17bo2dJQVNV8HoK7AYmWL4KFz6jVWLwXjEfzIVrf3DcyUHBtof3xygtJVJRBGVwrCwwMGcLxg/+OJUY7Q6uRjnjSHtlcM1A2QnVH99qx2PxsrSl7tOehn5Y/t/95TgtHn5tOZzeP2sM1fL1lbEhVuwe4g+tls6QNWCBDpg2dcnMDI0kysMz+QZnBKVgHAotCtnPSxX9vL2thzMLvE7uNj99JFAKHdz2alAvNbvQwz5VV9QKJ2PiObYw4ZpKAAvwguYrNinzcHbElaqDyRZZJz8Xw/M6hl9Wjzg9+/CpLnwGXg6OZRyhKzAvpzwUFfZg8KBzHc4vim+TAATZGxde6ZQTZ/psdVas/uKXLGA+OIMrjvrR43l4yZyiB1QufOVDmvJUP1fs1YNezCMhSuHV6LIEuVnzbh9OwGEukqx4pMm9Sddj6K3M5KHbsolWz7wPcTnltl3jSWDGJDTwSoYxCCwlhUAkwVPKzUOUhBUMXD46UjKKXnvUG0MkFYpcKuEKWZuos9WhkVe+y7g7Vvsy+GNg6JCmQmWQ8VEESanwYPKWUbR3Oh7BGXd2YWYd4wF9Chkuv8jjKp7KueZRMZ/5jzCCzb0Gh6ZqMZ2ejl3tiHNm1cnH/bvuBJrQzq+LmvO3Wb/dNtnAlRsf1dcXmdIy7Dfn7xnPa+LeXMf7w3097f210+79NetnzDl34mGvgMLIsbN4+X1/zD/3P50Z/6FU7sRAQuLpbjo0eWB978uuWR990PFnv/YHnqR7xouevZL1h22bBpJkBmWH/GK1+8vOYrPmdKmNiG+OlffMvy1X/7ny0P3zjeVhYf49+j+H+wSj95E+ZMPesjFvrJc3OMjYq8WQ5rjorRDr+rAJReY48Hk230k+NjPyjctBWYJFzMHpcG3vrerEfr3IpFYjDtKxpZlc3NWtBQdFWw9W9lW/AuJCoU1ePkAw8rNWhTxID9ArXUS7p0vQs30kxfwqhDA29nnC111OsUwuGrhydK21iDqhZACUafzc8j8ofRAIg8oOHLBnOIdmiJqcuICjsgZbRqPWAkWhqnyvKgrBeiWAdERWGk8wTgOuCUGJYM6/23ICL408raVydpBk6ImBgBN5sAjdVnTS13HrpG1jDiA2nUbHo4ixSowv0hIyoUfc4sJh7CEZndyR6GmPWAZ0RF7K44QK5AVPiBXS3l7hBy3QGiwvYc0vtxsMs57Jt8WuTao1H6iZsx9qQcdKXjN0s4MniaA7U3YxI8aOVrBtkIjNx0nD2KREVHUmiX2n9b3G1MVECFp/PeWn5JPLZETJiNtEX6uYAuV0kX06O21rH34U1kxBV1P+4hPTZyTUbnQ51n7nGWYfDoRpc/kLTr12wd1oAUVOMVSz/Rem6eu5Q/GknIo0lU5PXbUmRXBX7lmLfl92pUfTu3M6cSkcRwZLWX5Ph6P4u6D3nezHcRzlnJTB5dM4dWSnS1MzZt1O0/C1KqOHema0rSTtPjiVeuZEsjyUMQA/sOzTuzTEdd59WAr0iae3DwChSo6ysCRs/ZYIzbz1cXWLFRW24D6Gx555n94IBJeUzpxNgrsnd1nyuPKbMXHMyxuvUsYTK3aa7mUguQB0BCvVdsYy+vQeDxt52o2LBec/xiPh/gtUUKwzep4L0DhDJlNwEkMxJoQFKk3ZGCgxFmjf7eWY9ysnwUZVnLv9ITVoAKwW5sHsvxAeRDyaJq5wj8qUQiIqZBjisAoAZXNfaR3DAn7vh/xeSQqPAnZOaA/A7vT+AAETMoPYBLZyaeyoFIl3vUmFewTM4jRpJkS9trxJ+BpUTttwDB4IupLEdzthHgVFARZMC0m2wh2bPsBcXyPg76srSPl0I2AJpnlk0/mh1j+E4goJVxNL9WKWPPGvTxCdiSuXuZ/Ye5SXvdzXuPMPeeAyKDLuDLIGMK/T1EhDooOQF3JYPeP4Nld1CKGDXz7XceeU9QDpHa1iMCZY3QL8JKcp1EpLxKYQUQT0IN+gZPAhCUVR46n9zWDX4qqiGEmj3jXHH/yifX3MRM5kEqIWo0jHqpgIAC+Ir9kJUdHF9hSRztq0r+gKhDtoh0i8/Zxfly3QIYj0+QTdM1Lq9ZEZB7yPjWFUc6ndTbb/63So/xu5LfPK6sN4T190DZLjWjryXLzFRQ6SrHjLgXlU1kkh59e/zsgt9ghIYTFSdo8uzyaIGRsnVZtUClplQGDnsdwK8RY8gIwr4y0N6yK1wWVq5mK0+9V6B5lUes81Ug/OjoebSIigtm1IYMX1ZaUATqgj4YXo5tZ8fJtINDw97wCp+2KSvePQnPgpBh6tzs1YZejsoGSvljhpOyK1hyPQKdiLlV7Kafw5lPoYbt8gcTo5pkP0/s/qoxV/fq+nNEdpBl8Q9et+L/VDtQJcVFRsUaPZ6JCiMpPvtTPnb52i/69OUpd942JCluHp0s3/0DP7V8/4///HJ0nA1pVsJ0fr489J57lwfe8rrl9OiRkvYJpX3bk+9anvWCj1+u3fGUJkqzv471yfjUVzx/+fov+czl7rueNByTOZ4/+ytvX77pe//lcu8D799eKQ9F67HwJrfStkTF0wc9KhDWAb1cdqYz2YoS5UaOg9LA6AEIA7AeDHjWzDz1pmdWp5EhRjmx0fAHxqyYUJT4SoASYIXKtsxi+3kQm7FnoCVLOwDwyOiW/DWNmfrM/m+775ioQC8NM9R3lh0eipo4RH8AjEfGw+DVgJNjhSYjxdZERozfl9E0MjZUCkpkBQ4VAHVisQWOh1Lz6AWUpvLD3mop8pCyAzsAGE1DAyauxwugJsEDGAEJ5NB6K2vZZ8RA7nrjNhwav0AuUM2K4EmaByofUgdbdcRH7+WcwFDsiYq6er1TXw+dEVERv5W9S6MpmkZ7mvZ4/fXEA9iyDKkH6brNu43qGgtoRjKoXjvlqgvT5R14EReE3rIrnmYlKWJsfYmSzAppwcN0uNbWY9cfwLdu68C78Uuy1RE8Vy3VBOnH3k9M913JWXHeG1mp9berI9ODEVUXrEpe8ZmrMVQFfrK+twY+5fO2wQj1/fLvdmOsRtLIdZnKlnTQSq5cP55FeL9/np2Yp6zPHUAQl0kgNHRxqg9FbKk2O/ZwlvBxY9Y9xW79vTbhejfqwcOwbogKEMhRfqE6DjMQt4hZg51fkaiAJoBzXudwo6G80gX9G5dnvqaqHszhNvqo+45KxiRRkXuCT9b+Yq5OQ7+rFIDPC5vB1gjgXm+vh5310AEMMPJp+nwFxMwojZItegsT0+y/Vu+Hc+xRqXhK/385dhs15F/a/BwMU+nkqd8T/Xk0Lm82O/I28xoV/E2ZHsNuc1A59munh+c6s53by1ZqWw6h3k9173VtAFls+FobMxc1eTWHV2cnbGJ7KXJyg/lx2aO2n5d63sqi9mOYpAXeU7QhoslnYObsxjuTyZ3ZUBWkq9cUoD+6zxUCLQc/LzXdVRqEhvBmogLW7+xVtUd+p9pNlbgVSFxsS97cQV81uKePguClvHvKFc5FkBgMLop/ow+efyN6CGaNfZytJatC7mk5P6Uz/Xv9o3tj2CQqPOjEtyGAQz+jo7kGCASPYPZ+FZAtP79Zfvj4+ATlYPwaeBbpfZ/PxvdDYAS2tAAAIABJREFUgAEy79GjwkoTKUJdpaZkS0YwmogGV6X1jKqNckFwCyAFyA9wEIPYcbDWXvKbkVmAZ0aZXxgz3nvBxncBskTAH3xzSEn6z/URB/PNM8JtJdn5UbrJgknRyNaD5rhBQJpgDJbBEWVbAoBPZZX7HOdFnOlODGQpLyccWOseZWfgp+7vW8YFZcr0omW77Mrf5H2UrRP7TkcePvdodsmqgHrKPXx2lgtlJnRD8pPwqHsBcsMnK2VfJWN1L0cfido4nEUU1YxXmIpAfMm5k0MXFw6ky0ax927evBm9HQIrqHLjWUbSdO1ezP4hcxXfbMmid4GjwFpwf9nWxbcbdILIAiOiDOy3ubW9VOXDn5WBPPK3TZY88r5E9GvPyR7Hvs+MYD2f90YgERKBKApKGZRX1vPr915qjNk6Jm9WucK2oxGRVvUlXtzX0B1GljBwQiWivFm3EfLswcKId2FCs2oHjx5RoX6X2O8hr0HMduutMmgkKoxIMpLm5lHKljJw4BJd0nuhZIFSpXil0HR/SZSVqiqQXehvqGJHD6UOm4ohW0prfC0xKVzb9afdbdobq88onNyx2Q8Eu9hDxuYI+mn829kpP7PnXCdzv1Si8gmigvNrh9IfeOWLl7/25a9ebrt+uJp1W6uj45Pl7/zATy3/07/4uY09KWyyH37wvuW+1//scnY2yXLYWZZrtz91ec5LP3k5vHb7RrLCxvb7P/FFyzf+6VctT3nSbdOeFa993VuXr/7OH17e//DNMb42l/zH2CeyBAn20qCcln6aEBXhPHW7yQFeRiS6AVTqBdYIhDppuhaAn2LQJoIdusyVCMscqZk2DkE23ePv1XjKDjOAzv0LqaJumHjTL9TpE2DvSpDlpcJ595qCiFIJc051PRmh0BxUTFX01OAFTcWgBFEL1c4mgSrqTdEQFnHY6apjZEV1VuVc+D3oHHhK4vkFGsWx7qkaZtukKLJcabPe74MOit3NnleEBKJhQA7Z/MCo91iUnNwgjDRFHSBBYxkECQBhmwsYD0if9LJP3hQOGSIJ+fXgRgpfHUN1ansQNMGYDF5Oo1sQDCNSBo2xq6yOiIoGxCjDrQbGZUSFG+AxN5xaOl0zR9tdHGyeslfqfPVzV2R4Ww02FD/Vt0xjxy6XQP/As8QX5kRFFadm566JCnMqNJ+5NrmOPVGBMgGlpIBN2jnTxs3juKAeoJOEUmRwfIqQd5Hv/cT036XGoD5JoxVRx4jGUW+dDcfZb4Go4OXXWnCsUi6RiPzRNkSFL3er8Jvr959Nr1l+tVqNSNNudSWIikJS9KQQyd3YDV7rmo6rInRoVMsQrOCuj2O1/PN9Z8aFnV/aIyJ6FRnn2UDwYMN53KZ+v+bMHSPaw9NFHKRDOFFRiLSY3xmaujLg+0m4NaIiIYttlVJ+rycqsE5wivFqx1iPqno3e2Qv28FoWD9Pw5nPnib9b8YjxvkW602yYwY2xrxXPa6a7dsi25dOHccjPS2nMRDSPrOlaL56plFOh7fzxy7lN8VBx5f78+hqDQWH80e51p5y26GSixNddxmQ33++mai4dPKbL1x279BmApC7ev0oP0Giosh4Q8ZeRW6UDc0yTN4A0su5WP3u8QTOHOrZ0SJ71bVcqQOvfapI9q1KP02m+0NBVMyBhPGggpTp9hAIcZZO6sD8tH3TtgvQc3Cbxr7tdB62K/QRtgX8JvdFak9AAYkhcwCIBC46cRQy1c6CgjzMx0B5zSxrWKPWUWIjsxKTxEAdJtn9OkVWe7Dc9tyeg+c83VknKppIW+8ZgRIxyA4hoBu6tTSppo4WeGe638tZ4ViOl4PCZ6fL9WvXPWvEIo0PDw7hw5Sa/ziXMogs9BKJa9jK5bznUeXmKMsfeZYAA2g0r3XmPQrbm0mj7BZ8TKwTyiOdL6cXaKatsywyDixzmz192kc0oqJ38CFhqGjAoA1G5ps8qZl27XOIDAT41mq86/fxbJcMUhAQL72ArAU2y2YgnzeVFuir7JsCegMbT9sDpBOywqRr8vryL9X/QONh6SA+p/zDBKtJRpUeCJAVYhdFrt1XLmXlQo4DN8j5dbk5O1uuXbsGsodlwrwsrRFgpfyTR5uzh4MwDvuO7TfgDQBZrZ+DrYnNg7/P20XpJ5apEtmhz0WGKPPislOtkRKRHh1R4SqHPTltPSwbxso8qU+EYRbXrh36OG0e7HMDwg03USlwERIWxGqZITZn0bvDiAsjuFmy2+9xCExBfVFcDq00tpXAYtk0ZQ2GXDEbpcm0qGWKbE+RXLEJNYzE9VzpC5B+OMtpqXcMgz5NQtUk2svBnZ85BuKlrSzrw/uCrl+PFlEBPgKBvEGoln21urPkm7ItOXG9VRq2i0BkNOlUbLQPlNGC7BarbqBeR/hpEkWZfaneITq3pOe3aaY9tbuphlDWC2uhrJGRjYZzZmYBwNPofSjTl6bH1T/I+/icWX+YyVpPZi/t2vYLtp5RwYbnqxNG5rtUTOXxmlHxu573zOV7/tIfXZ719CcN5duE8O/+4E8v/+Sf/8xy4wh188evi+Whd9+73P/r/2E5O765WTfu7CwH1+5YnvOxn7RcvySzwjblK1/2vOU1X/5qH+OwwfbFhffM+LZ//JPeQ+PD98Xts2VGxWfchXWoYGCNxNDhrPlyEBBWL6NZCAxGs+tuc9HYUTaDKejKuI8AriaiYHfX0wRFMIy1exqBHiEjhEIRsRZ9U/wAN2TQlokgF0YBAHnPDT03/siK69DrnyyUuStB3dcMNEshyW/H3PaDL2CFQ6UyhOpgS6QG5j3HmilzLG+yqqmegMQwSrSOJ3BwPkcQCF2kP+cWBzdkAWWmGOXD5+7XNUmsmmonkLEHNRJM1BA3ZRs00zoFwVscq79eBSfqARUOFk+m3hiOA3lTb53RmPhejKNH8LrfiJgSy4pxWe8F7HdPY5UhZ4YRo4ammpil1SKF1oV5DfiZU9BEQZULjoGKUrDDIpP4fTimStNdbYSM9l35TQUEpPz7wWyEmtfDxX5zGWz2dYm+ZxNWgVqtvLBHxUiIGL3grlGJjhcpANlnfDENB60PlqWBIVZLga3UlUKCSroEHJ+tqn5MzUaiEuqkbSgfYEanF6EH9f3+eh0QrLWdEBXx7QKA5dzlzl5LQxUyXCXP9B5IzjmO+eTP6/1DDkchmxuMUqfABcqGLCcxUhcq9MYwHJyA+oBEUJZHJdg2puMPAcUaSduRCEbKcW+P1mQkTWMjvWa/lQxBLupK2v39ug/aO83cgCiDIK1Qzrz2CoTtuvmAYwYwwgFYgiH2W0UljnwQ1x+TMGqV9MBeYhShg0+94tbeyxKIAtbtE0UUqlSI2zokWmb92VZ3KITTcO0a0jX3GdSNjUul/HD+btQmVE/QH7T5IsCj/lJ2yWRfX7X0E1CEbmh1rO24zT4029LAuWrLzpw+u3BEXDbqJvdRDbwRyD4jMXqbYeOk8t7Sy/W74z2RY6r3j0jwiUMdq8u1U0RkI+LFvpyNWfa4j9fta3zTI2g33Ls+n4C+RytrwzL8Bcz5vuFzOPBbAMDMokZkpvyXKNU63Ct4vjPPxIadpXI3BkTM98x49aJUq4HdxycIUlG9fV1NvoDMgY3z2u/ZWkKolSa5QgLyssQT7HpbWweHvVwsevaFHheRYWV5DOxm/wEHxw2EYfCYnS2bQJ1ernz0thZ2XWbZRBSts8hElZjVvFjJ3j0AMifs56B+FRkRW7N1E2RC4+ETB9DVv8IiyNzXY2NdgG/QB+ZrHh+h1IueCT0QAKgH8KdNILJW4S6cGyM1oucCy/YaOG2vLMcCv7GfOy29gbAPP/KwA7Xmg964cYNlq86Wg4ND1j8XSH/uZI6ImvBTLhbvXSB/wfckswL8veUieh2a7jw5PnUg3er9m/zLVzfgNgIqdpXRgSoJ6DFgPrOVIz4PPax1t88yih4BajYH3kSaJbPs+URSjHStfHOfG0EcmigGJ+nZVqRQty09tFGkgFU7KJknPL1XqnCTfOuMSWInSy32fmXFPmxYNs8etGcAO4mJOEFpswvw1pllc2dzJQBfgTcqe7UpYNQJLRIdWFPYPH5ND2JkPyHiPCM7NDM/1DMEuImaXXvP2aK/UKf/zPefGiir1LEdJsgQQVaO7T3PYFKjcJY6s3GbXFoQkPWMQB8WVqrY3XG9igSgzLbE+bPr8q37WlkolIc6ceAc8sTAQa88AVmNIAweWAn4Y5zKIML7ls0Em9PLi5uuMCL3VD1X0O/B+0AZtnSI/jYgYfaXM282vizXb7vue8J0rQV1qjeGBXZaVop9X+WT4mydnBPKroLrQh/aZR1Avd73efay3/OKDrGfaFC4TPu/0dRZfTY9g0Slv+gP2/0s48ebiu+hVJvdu5bksusry03lzKMsdpQnY49JVjCBLlYGHbNZcMBPXuMPQoWUc7faTbBbmMng5xaIQZybKB1oz2PyZ6Rl8+KFzPvyEvYmhwcgL0a2n357lbOUR2nDsD8um2mb8vkH3/AFyye+9LkB1tTFMMPh+37kZ5bv+YGfYkOauaA88r53L/e+/meWUycpphKVF9jZWQ6v37l8xEtEVsyuDSDjk1/+vOUb/8xnLc+5+ymDg2ZZ7n/P+5cv/Zb/ZXnb/e+dX+gx/4lOcRjlzC+dN9N2oiJLAQgMb9MdE83yTUS8XKzjGgTr9muNqjLlzPqBTf1L7Fz8MBh7gA12kMdhPfOri/OOVPIadqof8b8ybMLIzIuinmebUujPN4owDYOJEd6hpC0KPJ+nEhVD6DIAHZpJBXhpn4OpakpTzaDGcM5hNOk6Mrv03JcItwEYJSUWejab9uThqLQ/ZFvo+SAb3c0F7DTZC11dwBrthXiwiHr2e0Ktb7czy9dW5MaGz3qDUqBhBT1kvNSBhBEwBA/5zdF9Z+912JGeodjnuUfo5EDUzOhSc1MaJxumLMcdMW0NeZczfmtEBQ54gcoaCLKf1q95jwqUaKOhpZqrkXrKKCcvrabIgrx+rCnLBWB+WhDXaQZ5zjEwn1EYKKoD29XaDUdQIC2N3ZGxMQO3INYfHKIiVWnOnbQBBWggzm6+htBWvR7PWxZPq9qJbJf1E0hMPO5o/ZsdPtynhXTtiI/QckXnttcrhNlvI1GRIHi3MZnlsTVRgRjZDfpwTVQkMa/lbc/a4cWaW+CPlI6GiQ+gsP3JrRMVWrEZgdzKciEleSYKkPRoRZZJNIF3YEVbfvDQM4LGjvYoqRHkVT2mcjfAh2ujiatqaeymUtN55HP2qzzNJmyeZaxjae40Z2lN519NRzySglPqM/XfljyNz2of95ZHuPTTajwNydfvoZzzjGRcg4D1mjNyoQLz+n4lNUb6fCs7oNx85oyOvaJyRgjQhjadAsRhB5JbhF0PeXU9VJR32lsbDQb/rUq/2t1VMm+9TmuwW0TC7A7jnjhzN9EjVtljAGBvZuxE5KVKGrlOuCJRYcC1MhP43ABsNqjdyUcOgHvJE5YSEpjFMWkt6nnqSqp7zW/dln7KnxlwbZnoGTwiYjQCXAh6ojQu++1w2qtdH/1omM0t2wBEQ7HZt50eNkVu5MHNOawTAr/gCp4tZzDbPOBEQKQF6bAsSASoJKjkfco8O9xAXZsDNKb2zG4DaOlnSP8ZQGtAkpNSJDzRy8Iy77Bn7JkBeKq0VBvF73uC/q3AKJtTRZVralSKV6VOxvpk8ah7A/AFbnspIJ5liOQHeRKnspE5rMufZXHs+Q3EtZAj+sW1xx97ECLzV0F6Bz4X3giYDe/h0KIElxP/LI/jZalKCTnPqti3Btn7KPdTLH5lCbguKNkFmhevjc/MAsiA7OMsGxehw8IIXA3mXbSe8D9aYZRWyn2cfr7KDHnUd39QlYyJ/pg1wNkIPDQJZi8T90Vod5dAF9e9BQtBxgl6Vfh4nRRtNWSQICr5IvyFJYf8eiKeBKpPsDUjBIyc8EwM6hf088usdUwrMyVn6rdBd3PPOoju8gESwUF8B/6zv2bvU/jninZnLxXJuxph24wY2Ra95ir4XnrJqWa/5kw9UStR4QD4LrNPSr8RNc72yhdNiWNaIyJO4iwx3xCZWzZlqHiAEmW2hAims1JxRjBgHnx/OUGSZeucVFJGCCXPdAiaoqMXDPZilqvD0b/ZfveA4F00Wvf5tMj+s+zJozJ1KCGH7I+291s9RZgNSNMubHPTA8wSMdGzZxYBEX+TALOfOtlyxpLaKstGez17uEIWld2nc732XNG5LzFXCd+wY4Zn0Pj07LGyapv7ThD2oL1QSi9bsJGN25q/S9+Pbi3sUL0/nBwqgQqrc/6KRgaerOAej7eMChPgj7z7qcv//rf+m+XaoUri5LSakP/gT/7C8h3/479ZbhwdT404W5gbv2kkxWuX05OjaRTO2MbZWfav3bY85yWvXK4/6a6VIq+/McbSyIq/+ZWfv9x527pElfXQ+OJv+p+X1/36/duaU4/B7wk9346oeNVdR6HzFMq7dtTK4ckqJs0m3gTS6iAha28KzA4KNWCrNkGAsuUwjgZKTLV1c2nto+Y6ReRwiUJrDA/7sccAxeZGdBUugWdndoWYczKgrTCkc5DKTg0e28jxnqgQoKz76bp4rNJsT0aDHIcgBdRfQ4ZnAjU9yH8lAaYT0ByCfckrn0ukFEYWSUlxFpPP2Yzbz8DadPB5CnZKtyzsdo8yBDn50w2fXUZUxBrR4Y/BUFY2g9H1KZpB5Pz03iojnygSCQoUA0XN+GD8qXk6j60OOK+TFwRmpHQzUrYedj7MQfmmS1eBgKY7I9jRqAPMfhO+WarRwPkIsq7f3G3KPDKDLJPBjM0TTwNHlDKipBp9EnNV27KuoT/CN+XJIOOYAtVmxnPYGYPG9AnZQheyZvAAifH1GaB02N6T+v2THhWXTj91mL7XkDycjxkYW69dHYrZPSuw0jx2A6a1ft9on9T36nXW36WGjC/VEjb8dyUxctMmLncpUbE+XGKdeD2AJdJX+f2Y10lGxYyo8OOHRFgLDo1nfgpmxtf7skzcG1KDlQifGMVjfVYBwWwuuAK7taUvcZxnwNvVQN9s0JpnDmutG4BhdZFVnoHZFSitMdiol9DhAcyWjIpxuZyqAwEKI509CeQaBe66UbpgtOR9AMf6OGt/NZzYZmcx8lBqrNfJ3eVKhlUFTtpvlesPUOfskDLXYHVJhoT2lkRF6OJJ1sRUn0lvdaW4KunU2AHbKOMrfmemm6U7GrndYHdHiQaqqbCtRfwPdMCsXjNqS2NFeqBp+HgFRMTZV34/mY+rEhXWW8odfgOG6PTHpQv5H2sXYdjY5BsJugLUe/mQ84vlwCO+Ad6Ogy3mbq2AQICKyKqyf9cSWXVaZiRW2ByD/d0S13kyWwYIoo+pk5yoQsCI5s/AOfs8+hho/oq94OP16Fn0UbC/LevcwJdaurA9TsYaXiCerYIB7l5+zAHCtIf23M7GmC2K2pLizbwTsMnKfdl3EAURYxEAwLL3ng8KffpUctWbaRs4z6wKA5b1fZdZBr6AnQsHDJG0JwYCZuS2zy3nTGtn/1X2noGsiJjHMyrTDxyB/NRqTUEaPBtwbzdL4LA8lUeDe+Q7/VSRTFZi91wVC5QNtIc66fQRRBLgDpABjw4XiFnsVPWb0DOZ3B4dHy17+2riHNqQ55sFIRpxwXJOtNWVeWO/xxLh/HUCh305lGEh/VIDxfCcme1dZcwlrJZ75WGqc0ojDJJCyTpe0oY18YOkY5+Fla2+IXNM0dYsBwbSwIQ1M8/q0Y7MLK0dwGsbm2c5sI+nyziz420+VEJGNqL6XMRZTKIC9+lKjBXFgh4riPoOstoTmDC3AMXRl1IlZkbq2rcpdYivn2UQkHDR1GmNXY6pXwCYAxsRBqSsNXc1WX5QPSuclDtF9Lnrm/395dT7lCgqHXtGpQQly5o/71djQLk/U+5pZY94Rkb1F1wPqek8iaaiA23snsXvZ8+CrDI2sXeywvtMgmSNceHB/G9lH6FEIEhr+8TKXLk/e2ZNvKFncR/oKyP89naBv4bbgVN1mgHs/VIpVw7671j2ExrdIxsH5ay0ThuJiipTpSeJryebmXt2J9fZ15G9QrzfiPq48js2HSg/DpJNerieSSImYMslluffoR5Pf4uqf0P41uxMHREVo7O4wQJEKLGSw74/H0rzjV7nFyh17uvHIO3pGV/IkeHFBm8+QVTsLMvLXvjs5fu++b9cDg+6tJbF+lKcLp/3lf9oufeB35zOqS3IzYceXO57w79fjm8+PLTmqhE1Zjt2loPrdyzPfvEnLLc95RlTJ9M248te9Ozl737dH12efMf11Zis5NMX/9V/uvzSm54gKs5Pj5azk5vLZ0WPChlKbeocJrEARCWzoB6KMDBGYgCQrtZCRORGNoTSr+RMISIKdT/9kOoi7FdERXHk0TwNY5ZjIAImRrdryu4MjpcOeZaHQcQl+ih4czOLiDk59rTW9pXpb+lE1ijTwnAW4A62+KDEDh26NpojG34Lz4TSxpzY4aXeBdVY7ldh5ljVeeexTGCZTdj8Rl0TcRIViG6A8Y9IEjo7+5qDHlTsRyUwp5bg2qSax8DS6hfla7eaUeEyt2pazJ0wICouPVCuMqbJdz2CqUT4Q0+qsSAluYvinaUA4/lKQzlssiwPE2PAGk8CdCaPXcqTKaoonE6t9ZqocPkdoRW1BjKjirycA6NELKrFfmv6xJ1Or7GZPQKgQFqQrh04x1LBZdVCdwAEu0fyjmgjOgRNZGpLOLRA6IimKODkANhf7dkpktNppQ3gVQXBV7qsBOmkvs95G+2H6lo3u/MKREVPUuTf6/0+erT6ff+8Oh6h4Mr8rzF86rFxn4MQ/+Id3zJR4fqUe6oswI6dR1Dqof43G7KVeBusfycrOHMYTdXt2tl91kA+xp1n1weXqJgRCWulMyIqqNAIcqmOtCZ4VPInz8KxWhMo5J8WoDMzP9ZXcPuIzpirN0ahy4GOMgMdubg+08pe2CbaakJUqHwVbAmdvyApNqgNcql96ad+f9YxrvfuVYkKzEH/IHM9LptIZ7dK3NSyGSsLZPLQcsD1fZ2jsHNaAGN29s917dxa6O9LiwMzQSe42ReXLFot25GZmd6tpvGh4pkmjSURyU6wrmTczp7EZ6ibp3hv05gHF5zZrjskdt1Gj5r6DCwgiKYIUd27+hHbEhXeRJURrh4YccXx51Rkg+kGBBxcb677e8C0ns918vJ9nRTaSVV+EV1cso5wgHLrFXuGtrDZoOpvZ/6RRZI7eRN9vvKn4/2Ldz2ohKCWg9emp61muBrOSmfS97PjDOWlqo2IaObM6rHVTftSuhUZQACSRMTAZ7EyJTAG8CwHzCAAMGzrbmVovJSY9S3ktAiQq2Yx3M2okedAo71sfgDo4mMnTzyCOckJkQRly4TeM1AWWQ27JCysVBLAUmW/KCsDHiGbUxMctu8oehz+OUDxWmc+IpZJ6NuzevQ6g2ssG0UNhvcO2GjYSpnYuLzHIGxh9dXwjIiz8+X45MRL9ahMkd3fS6ZwIj3T5OQkQXK/L4hAvepeU5393pfH6aU+lcQuSMBU4LDqEW05u6aaGyNAsJSNbnTRnKgw+XXSi43bTRaAi6yJCuw9gM8OcDP7xAFlI4p8H5lPbZ+RRHPZyoh3kynHJvZQ6lcAPPaVIvfH/cO0jup5ofJm0oUW8Q4SzMhflGQavZyY4BjV6B183o6bt/actpb2PfUSbQBxyqWTwNxXtu5B6Jn8HCubKAF+Wy/TN9YnRiXE/blJfkQPF3+PpYGIS4mkVFkxROUj8EzkmV+rK2spebX3rQeOzZFk0cv4nJ55bxhl6bgGtf2qIB2dm+5DipSVLX7hJIp6jLje8AbMatoNh8B8W8vMqK96xo7WCPLenZ4KICCOIJJGOkhZRf31AucrlS/0nuRPetF1wYWVgTuIDAvTQV7SCkNy3QLdkX6PsiKctKC+dp24QAf29pTbSiWjLsc8Jgu2Iyp89/qlZGYLQ6wlraov7PJh2Al7DI3W4vTsxHEJ9e+BvuxxtfIE29j45UZPEBU7y/Lce+5a/re/+UXLtYNxRsVP/8Kbl6/62z/szbRX82skxcO/ubz9l/4vr8M2VHo7O8vtT717eeo9z18eeMsvLyc3PzBJZ95Z9g+vLR/50k9ert1pmRXU4Lyo/X3n7deW7/36L3Bypbf/bGwPvO8Dy5d88/cvb7n3weFYPjze5EZVuiIVpddkPD9dLrzZy8mSREXf0Lx1MnvHSOw7mmgng49armsHVUCnO+xk1J1ttZp93mQ2Z12Hgko1aIkB0Kq0zSCjIop8d80dk2KRlOC/HoGRabsYN9IhsxGuMf+o6YdnHjjmTFFOkKnW8Iaa9dtdQlTUz/M+jAotabrAezuiQmBIiZhpD7Sx4q7fSSe2rf/uht6EqGh+z4h5P+jDWcj9CRte48A8JreUZMxmJ3AkW4MdO5Cn+NaGz67igPp3da3Lp3co483Itxhzg2OK1JJjp5Tjki5/mT8tE8YNDZJ6aFytkVWn9SqasRAVSnCgE2dpwYTHygUlD5uJigoWoem7nNKSxUQ9UJ8NVscc4AowbEhUYA6kH8yQRFkANJ2HA8qI0S4SYryn23ms4E04uxjwOmrzEqLiMvmtn8/2Yju6SlhLj/Vls/CLgq9Tv3JNqyhJA1cioRPS2oei6oi17s2RVnndhqgYRw0rbX/1JMnTfVCJChKHDVFRo6falRkH7hQZnzTTvsouHn/3Q5NRsf04qU2CVBaYnmJo4Jp0h2QF6e7j82TTKaPeFwB94MyErimZkNAZBHCiSTGcIIsgdKKj1NW/7ChJ94kzc5kjsyVR4eCZ+mMM5yOdtnxmOJfr+dNT9P/FmGU3blrb9RC2JypkVNjY+tJPl+lG12HdnFZHXPIzcnYTdKw6KaVoE+G8IIktAAAgAElEQVQ4mov19ynjt0BU6Pr10QAkMQioZhZsWBi3D0jYN+fUBjnU2QZbqSU6tt/fK6glfrpL0fD5dyIH9rr9jT4SyNz2zwKgYdR+iQqF3IxGpHHDztimkeeUVIka+KXUDKO5R/fenqjoDtjVvmcUMfe4oukBLmWde7+K1tIVF+esbkhmgPhcVHKDuek5gxXomRjHsgc59YqgBmnigwlA22V117Iq6Ce4rWoiBTwi1lYZFfEeop69HAsjs70Hg4Ovlj2CTFyTG6sFf3jtevShAPgMsNitO+pJj+Ql2K7o394GNFFynUq7EKWYrI8DsjCiATn7YrRz2cZxnlp2hEdi7/s5Y2DftWvXWQqGvYZog0InY29Dr6t/oNXjt4wKk2HuBxJ5LgcGGFI+7Bo2Vouqt3971PvZ+XL92rXl6PjY/WaPuncsR2VuMJcI6LP30bciosgt29lB3vWZq8bSDnp7n4szB6FHNdxBSNn/WyLD3vHySREQkDYBbPTEQySjyDohSM3gC5VqYr2pTiFszqiwe4Q8sYzPzpKBvZJpn1PP7hTBBoPPI/SphxSNj/lVkCeJtcicR/Q2Ivixx3UONWX9uqfAGS6cA/OkWv+Sw3aM474FAolVnidsCIsWZ5ZSlOfhPfTcwFiKb2H9JU5OHNg2+XbimbpIZY80bhEkfak/6QB8TyXjSNoZMG4ZQ+rpQXlwG4FESs0+lBxVuw72i60x54yBmchqYv83GYS+jpbnz/ODOsTIJz+T9vbZlwQEjIhM2y82j9lDKIlin+9Tykg9c1eGYdXClH1eBmuGZ0idCf1pgTwehDHJCIjzqOnNltiWdGQlHkR+uO20gx4OICEhryLrTb/YC6URmXHm+CDmy/a2y3gZd2AB6jNDHb0poLKWhqzboh57PagjfNNRgNJ7w3AAlzOTY9u/RlR6DydkjFWTwv/cBREp0tbJvUEYjsZ1ZZsRJ2E81uO2R8X3fdOfXD7+Y54zbFJtgvZj/+5Xlm/9Rz+xPHyjBb2PHnn/cu+vvnY5emSecXHn05+z3POiVzgJcXzj4eX+N/7s8sj7370OpuLy7x9cW+558Scsd9x1T+Ms3fXk25dv+wufu3zyyz96GB1mm/THf/rXlr/69/7lJQ2/O+3+mPszD2ZEEOH/M6Lis5/REki5cQXGtqCTRXlIsWBjq27rLOUQv8+UWxgJYCpbYL/GHatBrn3XU0fJwPqW7BwLOKJZk7JpUGaHF6zJXEl/g+P18wQKFMZe1uz3GxVyYC0KZqSx+RSsZyNOPfJHjDbOrZzD6ji1YKaunrCFmHv03NBBSUPMMyr2woBHjcX2GhFBRuhT812BkWZu1KMCDxFy0zr6fBavJ0knjs2F/NCmAK3GUg7Y+hlInjRe5tttE4RUflWXufcCN3xWnxHOdbmmthQjAGQ4uSzG824Y3+C+vSG0Ij7633DSBADAEYJjrkZlim6BzJnMZN3mfl6x/2rJMAEYVYZIYsQh2D3jEKiQfGJLynDE9mxLM5UNOSyNpM/N+DWj1V5KW5UTKacw0mo9ZEP3lsnADKGVcEFv7Gwss6S9jLlyA8tJXxiCchSqLGjP132GWw9khHrDP6mkh/SZ9y+4XPZHYNwMoJsTFWPzScvcZ+g0eqTObdF3/WNjTF32HW+riMcWsKxllnSTEQCyXeknRXg1omC1nnmurfaJTMAe7cOCYW00EazROwO+oOvw/M10+ZHTAsBy6EYyI9Jyvaf7M4R/s5F9//1NAO64mXftpzLKqCDTwserUdwjvT6Bsda7VLpvpW+oazqiIi6ws8BB4JkusH0TUTFzdqqjhOFAaL1sCu0YOFTc6ZHdJtMjz23MEmOdTXxIePj7ZbvjbM7piD8LQdJOFjfScGILmOHlR9jXRyDmaIFKdJnmrgL463tXHdfK+AebqPC95SUrQGInOI0SKEP5IyiaYqWgCcwjVHNPfs2uVRzFRoFp1drF3EwQdaO9AJGqcyXlu+7H7jcBKrTve4gO56rf/zOgIkGs1oyefR/aLPeB/y07CU+xWg63h0ZTO1ES/lWenWjKjN53pt8FzKLUBUu8BDheLih1VUq/1oFZORM/89m3wKPFvRHpRAYmyiNInhLdKwC9tTOT6hhPhcDagTQL6dRHuQCMzgZwpjIgyhRHCZCOSCpERVgEAvyVueolkAxgtKxukgJ+75zfGeDiolBjfWryhgg5zjKsrIvllKAs+kYYaIfo/JwxgcnVr9PzIlr7tuvX/TzwCNhajoZ18i3iVU3TAcYXgoplWMzOtGsJ+ErXMs8iNR4XWG8g7I2bN2AvegkWApzuPw32QkzhhZe6sd94uRuVwdHpQ8BboB/cNjXAbhvBO4Fgmcgs9eM2hBFAnrWx40CxETYezWw9BZxIt94AJ8sdt9/pILJtE7eTrHwzSwipoSwC+jBwB5vplwjMle4KPcDyUDYmrYXmXmcF3LASeS3bkeenm1/sVZO2eAYuNfJXt30pEavmxI5POGnQKxydqXy/M5Hlj+n+GYGX6woXV4GRu65DbP4MnEU2BkgHl2r1xHMZZdkjWw8j1Ux3n6Lhu4gAlFFLUmNGltr8i1iAa5HN5L3RM8t67e/u+/VNh8Yz9cdRKbdkz4E9BTzCsgtUMcP+a3KE7Acr4wTCDLKBAJLd/X3fG9evWSPpIxA+hvWc2TNbKap1A3q7nuZJ//XsD+tnw54yKtEnO1qypTNPpbV877g+KeRonP2w03zuhIeQoEMpTzbeNrks/UlpVvgv4bsegJCwRtpOllrWSjXsUgGaTrXn1tlW+z6I8BLYH3M68sNJWko2lIFlcqhSf44LGklAomJm+1asws8KZmVB22f5KQH3ssWiIXboOID6sNOYyUd9lAHBKEGmNUnkH3027H7WZ8XkxzNySs+X7vhppHZboiL5JgYK99e3PSjcy8gK2TYRGE67h3f382F3QcmyvX3vOxSk3SRG4qpEhdZBEYOPS6LCJuHFz33m8g//yh9f7nrK7WsDk0bNT//im5ev+64fXd770A0X3+ObN5a3/fxPLmdnlmmxtjZN4O942j3Lcz72k8lWweg+Obm5/MYv/9/L0cPvm2ZW7B0c+u9us54Vu7vLwf7e8t1f+0eWT3rZ85DK1b3sIHjLve9Z/utv/KfLQw8fDQ6jgeH3mH2Lc71lRsWr7z6O1LnTU8tygJGBw4YpiJay5tEgUDJNX2QqIR0AWOvqlOHfOAjgpMiP81ReMu52fU+xVURKl54uQweqUUoe10baWDZWi5JRlE0xsjp2PJXYmX9GY5E0EYjlQAZgXJbbYaaBM6gNd5mRP376CxzuHMgA7sYODqclorM9/RAPvEoRq1fQrpKSF0NPayAkOH+DZ7rayxpkrX8hMsiZc6aIKhtF367+eqa7Zm+LBvChA2GHtCKC6l178LK9h5yENCwwp3jfDR8/2Mw4gmyvHM56AxEubn8g9doPg67+5yagT9PshhKJj0rMpePOyY3/lMnu5704nzk3jICT8R4T4zupkwFIbxo8PYFXJUX/Ls6gC0LR5e2ixL1cA1Riqu7X8pu5JPaflHHxn3b5rEGsiAczHtVcsADcqqrTKq4AG2tZuio3jdTLT1FTXVmj2rzSQ/G3fi0CVyRoGsTNGvZbzC2mGGIzty7aq80xQXT4PekT/XbkjrmMQ9CDNEnittW8uGy7TkOiNO6PKE4YdkBkHQQkQKWzQRFz0g3NfzvZibH2c+fGIWuCFjJO4+2vKan2hnMEBEH8kpSSLMeZas9Cks91vs5cdQVEiSSRsCAz6lzN5buXOYEb4WD5+AjfCEglMydgtZcrOfMBsEWZwcHE+bIm2DPaA3ivtbOSmNddWr02BSdXQ7CIP/Z7KXrDHRLP4oTc2H/NUXHwha8MNMgsPYjzvCdFe/sZoYlv9aS0xjSZxeHbkJQLBk9wiyfa1dgXVduO/i37qd/Tfk4RCKx2Wd3zVR9AfG/BLgidmOfK5EiQSilzovtxRjqF5OSxR38iIrmC0T3RytWZuX0oGSMyuvy7VBdtFC3mbGDDblSxo/lre8PUOU7bp8y9SgqOJKfxoXJ8CSJk0AFKmnD8BAUkvzZ3s6aZKnuRekIbS81CUbbBXn6PrueLl3Pd2U3gw3WvAXOYhwzwaOcKHkNvq7R7rp+Sqe1F8GU1hav5S6mZyv8O+x50FwvSSHvmssyUgdzIS5IsAygFsYp5HZRv8WkDiOwZ6Vb+hdHq8tcA3Blgh3rpvncIsikNzO7tYKnXRQdQHRlenYlXH126q+pblwcHm/ApTN20GQ1cN3DOXgbwexk+hXEVxn2TjnZ9FmesgvUFJFWVksahZe/6GWHNsw8OAJieolY9ZlGGCH6/a6WHTqz5M4A7zYvIqQB5uUb2nRPDNqx8z4E1zEVteQSb2D06Gfc9CdvUvm/zf3qCKFuVOvFsBosq954R2Ev2UhNt87WMTHAgzxu0m78MW8MDeJjtoIhdlLuxEj4AYq18jK2XlWWy8XqvhGUpZXZKtDVJEC87s39AcO3c1xDVlfO7XtLGI+NRLtnnQpmMrI3vwDrlwiPHiTNEI9wSBBaZ3TaF5ylLdQv7uc/MEScs+Pss+6qSZuPzJXslIHrbrm37yQgZK/Ns/7a5tn9b6RYB1bv7ewGU3rx55Otp3zG5Up3/g8ODiCC3nh4mI1YGSzrYtZ35o14aF1kq9k/0LjBCCY1A5VdL31rmwfXr1wPkTfJae4CyPQk+EBnc43Gyp5Tto3EKaHZyUP08PAAOO0h2vGEvUYaHQZ+5K2UbDJQg96hlDh3s7bv82r5wOYp9lDvJ9RbPNiNTlFVi90IAmxEjaJStrA2Qe2GoBD5YiX+QbTirrLSUSLjw16nfvD+hkZTn596zyEYG2TkHRqKSmh4cC/LJXsrsE9Duw1GGmKsK9AcyvWDXl86yj2zN1fzc+RDKhkpbYZ6rrkEgAs4IkEbAU1BKTP01em8EJiiyW0w+brvtNupLZGfJR/ZnYdaQ35nZEeozJDJVJf0C1C8YSj0/6vnS/1ty2pBvNGtivyvLjb2DbHzSQciyzDLm9lNUfjGbhPYG+9vUe2tufD/oPDg98znA80OfBpZZSQrinzhneBarFHWLnjTBJ/GsOkfLfDkeW2yuVVwls3qsZ4qP6vHWTFuLt7+3u7zq975k+YYv+czlSXdA4favk9Oz5d/+3K8v3/wP/tXy3vc/spwcHy3vfOPPLx948L5SpoPbyss9PWu558X/0XJweFvnxF8sJ0c3lne96T8sH3jv/VOyYv/gcHnmCz5uefIzP8qJij/2Ga9Y/vyf+H1e/qk6SyZs73jX+5b/9jv+2fKGtz7wYU5S4ADhOYLNJCZ4VvrpGUdMOTPFhtREGEcA/uVcBMjkb65c3kI+6LPqiGa2BQzwVJOZ/aCIv945qN8dqzU5lhVIgBNfo+ISuPI7GFHBZ4Wqx/3BkqPZT3WGPCqATgAOcs5NGOUV5KhhkWX8G8AAAT1ef5+Hhv1SwFl/HCl7QzNi4zOD0h0WNk8LYC6mbW1AbzooMJBJjIbYeNbMXLxMVgv01H1oB5ga8en5dMiDYYbsIhKC0f2NnIyOki5a1YPyyhEcA5CxmlFG3tOAUTSc8GYqqixFuRhFmvGbQ2eZt49IjBK5hftwew6B/AQb6ndjYLG1OjOjvp82GZ1/OpBlXvzZ6jTxj4sGCNYXbp2oiFtM0KvWlZtJYiuzcSn1qKjZRqpbSR0o3eXcRcz9GgBoJHyGtJXh9YZ+AuA5Z/n1SlTMdMF6JtrmmBO9N94S0y3td9HzSf74d9XWugBsaM3/wNHoCON6eZHTmHZco4m4YV18OAjY+wC/Vdu3zRDDMOr8cR9NnhYkCJc9nkF/c1S8pp8U4ehiLPH36Pqxx2xvxIZOGauAo5+/vzWiAvOK+0D2kqiIBqgByPfyDUAhIgU3rHc+qoz47uEzaXEACqd85CrV0o4jGR/L1JqokHyQLCtzISdbczPSyVchKqabR1F1YSuonvF2Wiyuy3NudJ+NxPfgB9jC7Vmgs3NEVDSXKHLgMjxaik2TEfKmMbTkUP9Tcp/l7bXGqUCUERVujxHwkgw3NfUvGZ8+nj5ae8O42mxFMU9XWW9ldtSQ8XXma6zh1kRFPngQFYxUtU+8goLKODAL0EYtcmEmZ/VIaMgKZfywvrTfoxAV9jsDAJSpZKKl+uZqAqpSNHnvnEdoszVRIb08XObJOb0+m/nrCVEBvdGvqd95WSZERc6tVD518zwkdfgIqueu+ZO8Zzbd+meow242PnosVIBDfR/ST8FzVFlwXoF95RwYZBNlgWHQH+MdM/IE8OSZ8SMiSxHbEW1tvhaj7DHnJJBxuG3cyUFU1OA7AuUYafp2eVLgrFB2g9fAt/r7CmTkM+pJw95nLXHvCccSSRGpKpKOZYrsWva8p+4rGxEHEsZffZ8oi2RmRLkRN+qNYL0xjJyw/XLtOsBBmxzzTazckhpy2/gUiWty4hkOJOxFThmDYM9o8uGyVPph4PlohzVHhjW1BoGEdVGj61NvFhw6lPvdSAQEccgewVoCAL1YDg8Mf0H0s5XrUh8G+ywCAc0XpH/tJWdK2abIuibRDnmsCB+eAYGTJEC5D2CzKfOslKls7BbOAudQoKyNwwBrA8qVvW3+6eEh+iE4SG3fMeBYjYkJYtZGujYPIud8pAbkEiCOklbyt8JPAZlrmSwAo7PBvOw9z/Zh+RgHr6P8L3dgrCnI/dFL5F3/Wez9su+x5wDMYn/b6ZfYDexJRse7+YCsqvOmj0y900CnEEfyNS9Zok5oRWZVPeuoa7xvTJbQ8vOGvR5UXsfBXVV94H2qDR1l3Xh5+fgim/Jchf1s/6/Eja8zm17rc6pCEIxB3LZli/Q0tYeGi7dwAjZb1tnnwZV8lmYGaVBl7yqqnWJfmrygPxuJw9r/pRMCAe/IdLBnw35WqbvaXydkmj1RfFW87whLL7KUm0gMv39X+m16TvfjqiR1Ue5a/1rmE2SMsrmgv3FGInNNuk3ZMAhEQ5ZGffncn7NcE7PZ7G9knzEYmfMfWeOu/1PniGR222Z2nnbvx/csY83LVqrnEAOkReYOtpLtoQgRe7wSFbaIpqg/7RNeuHzjn3nVcteT7xjaFibc/+/r3rr8le/5F94PwoTo/tf/++WhB+8N5WnK4vanPHP5iJe8ctk7GJMeprVOjm8u9/3aa5cb739PGwEcErXjDOyzP+b3LHc87VnL4eHB8qde/R8vf/oP/94gK0yZvu2+9y5//m/80PLW+x6U7thoFD32P5ShBEPtMqLiVU+/6RsJ0fgwkKTrACyV1Eu3v/rGi+1Bmax8dUSzrIUaVsFQhXGX2BkMm72aFre1X1gdZRgziorze2phadw5Q0xwHR+ls+FlUYshJQLDo2WaZIkWJOBRoaOvJWQuiViUQvNoCh8ObuQHJ2vaxfthPWZDZAPezSmUOYpJlRtRDvuRvdABea3W3kxUoOQOxujnSLl+9T9E7NiaI5oFkUT4Lf6NA18Hbnd4NHKQf+AeaTSPiQoocYdCaWTD6FP009pZAmueBNZILzQOP4fURyOqZmjNpsC25PN1vxtdM+6tKSlGaY6rOmt0UFm3dxQhORLHCo4XmDdvH0uisY83Zy9i9VvrR+Cnk8NczlXZvv5PM+adPCRRKGPOyjXkd7kHGoJpA1GxBUkxPx8ywqyRQcLKHkU9JIJSfuu1p0RFRzDEr7fUk9Ovdc+u720GT6uOX1+5/a3633Ce3BHFWZJciF2jJyrK+TIgKjaBHO0zrHWGyA+dFCE3JOoRBQiSIEXfdFQtDZcHgrCAdcm11MX1rMn1nqxKAWbC8C1lC+Tg46jLBp2tjCprsMW0Y+VG+06BCP2wPlREhcpC8lzWMAwkUV3mmuUWx2FJ067OwVWIin7vxrVxukWAAk+pW8H3h6TAraieNVEBbcCqySG7npkgx7kKRxhe7bndys8M5s9dA8AM8zN70a8rH1fdMf4VarqXzNdCWsz18Paf5Bm8tpNGV7lloiLO+F7Xh4YKtQCAaDqLkw/wiwBizjPCHaBelihA1sTk3J4c6zpjHVAXWMuSSgLLPbqfZR0U1WqXU4a7asAn8Z3a9kNCVAzFk3aSP3edE8q2ExX9q0M9608nCzdfUZSaCQDFM8O1duOLOVGhiH9Fi4b5CoDYh0TAS1njfgKpPMkFiCQv2yQAidlLGznLuWAmQGwXkJNEotEAI2RKo0GvehBKZt0G8Aa9Bliub2LvwJctWjeIANYw6kTabXdG3KvMit1bgWC9jjtjbX0HMBl1iwj3DH6qoBP8svSN0aiYgJyvY+pcPKemBZZdbaZs628guYPip6dRfsoyH7wprYPo6FdhF7L3lB0i30vVDox0cIKhEhX0ezyz4sIyALAWHj3Niag6QTX9fb0sYpy1891fCyKAdpGV22GTdWT5INuj6lYvfUPyxeYQMgB/MUoA0e914FC97OKIgP0EIg8+ccpOlrgVpqDPYgzdlnXyynxql0dExOtvb7quc8eqdRwcLDePbnoWiT2bqky4OinBipD53GPKhrDfhLwzC1TjkyzaHHhmFCIoM6CPASY2Xie3+LdF/aucECeiE+fxRm37R3IvaV26agEhszYXnvkBLEiAr68xsSD41LCNWBVnrTUndqaD6fvwyUQeqPqCz2d/JRLitWeQSvMpCNbmHiA5Kicosl7EnvQtMjKYWUSsxW4XZaMYXyC5kgz7GRhl9HYX9zlpq4NAwqils5peIgpspU+K7Cf0VfIeErV6Q+m7JL0umfbfee+d0vA8gTQfD8oNMQPC5tn3HG3Ybl5trC77e0Y4wLf20uJdSVyfO+7FJAvLQrGsqGWnmc9iOs2uoUyLqmeCDAr8ZqD7g1Du8CD+RkSnGm6LuEFPmyxRZ/OXWX9JWqDqY39tTI7Kqjlx6bJdmpwHEcWM+qZsfMKPG0uedhhQYF/U17AN2NvHM67Y366bJp/THZw97hM+nokKWzjLXHjl737u8jf+4h9a7rzj2rRnxS++8d7lq7/zh5cH3vuB5fT4aHnXm1+3vP9db3VxsHJNRlIcXFuXkVoZD6cny/1v/LnlA++5d+oI7e0dLM984cctT7n7ecvhwd7yOZ/60uUvf/EfWG67frg89PDN5Sv++g8uv/Qmy+pY6c4P0zfCmtuKqPisZ9zk4QgDw5V52OdsfINcTxrRZrzVyUwgKQ2FjLgQQIfDAel1cmzFhsIIyeXIf7fg0iYWNhxxptElIFpAoogCYSpbyZpQQyU3PklU6PB0wfWAIBxCWceyd256kcpDa2sgggcgDkxkeESqfgfUyZEXZIAyTEw/HhAVMyxh7TyW55hkVOjQT7JBtUZrs7O8jlh1S2+057KUWDRhgyMNAyjrMFfSQkZTkZD453ZEhRrNweDy+/UKYbBAYWBUoKeuQSO06dDAeExDsCEpYMHAkA8Ao8p53QhVnrSvO5A0vtKScbjJOjJaoAOG2N7XIqD0aoiKxKRggOXmulyH9vO6ickaXq3s38InubPOxoiI3kP5gkzLzGywC0sf75pvtzNbGpdd/kSNWZOGV6kj3pnXMIQ+OERFQF1j7GmLp2lJuv4y2xAVwiVW2o/AC97PMwHAPxx2x06C/PZ3+N2yiTTEDyJR0WdrIAqpRsMwy0L7Vw+rbRlbx2PL8MT+bHRgm2yz1SxP18n1hIxgRlzjLC5EqgFW59qkdJKKsudohveYubQYfP9pBV/6Z6i6Q7e6tYwK1hTgRUqpyBKdVKPjYik6okJnVOi0osfHE17tlvU3YGPUYIVNoPLsDtttyfZbuO94Adv3PaCxREXDiUnH7ApCcAn5kPKW/vHcyJ4RFWm3tfvdnsJAbtScxmnUN4O8lZls9X7+tZ36HJTj6YIz2jGpREBdPZ1ndU3DENgQzT57Ws15ni+1CqpOeZGtm2zo2R1mRIXONAQXsTwIgVCAb8hMdhDktOjE1fmIiNzYp7HzqYEGgNU0sWXi6OHu3T6qYPdwf+HcHr2GO38i/pu0BMAIAdnwFwCIT1aDX7Z9YYA0AE5EjxoZUMvHGAhYTwUQFdAFDnYSVJaO8HKo8vXGD73hnKLtXogKAfsCqlHOCL0SfGz0B0VG1uzxZp+OwKpGANa71+0LnrmwTwBw1/K0bVCTlX9iQ2g24IXIYCFQE13ltHCueR1/q0FPn0ZEQBK3+RQI0MoyNNJlVnLKwEb4JFr7zGpQ5HCdDy8/4wArMh4A7BrQCQLEyuLYSyWjFIBogzZgXmCoZ5XvWamULIWi66KxMXtJqtQiG8aCiECwmeTJAFE0xoV82djs/1jnbI6rucw67SDe1KvCGl1LhDKCMdfXwHz1blDZLANVBVBUHGBGVNiaiiBxn1mN03mQyW4QeeG+6h5qXgswtnULv5v9ObQuHg1tpblIBHok/sH+suelhWyd2NuREe7420gg6ahyLtlvvPwP/Dv3+dnrwLOVhvt0ZtWNMy0qgG+XC99+D5kNGRCRGYWRUeHy56vq2RTIThvsxyFRAULLSzOLxGH/GMc8SsXGeMwo4cZGhMyuEZbkuEE07IY/KHkBtoXDZJSpZPtZ5UWFP1TbRrJinxkA7099du6gPlaO5WyZUQFiKdc6yuvRpvcSaL7/0HDeMxlO1ZSZBLaCDLguDrgz86Y9yzHn4XP42OxaOBNcL8R9BmFw0ZaU5eI8G8PK4TELjUenSJwgHqxku5dbykwMW08r32Wvqr8q2YzBclWLuGILtPKr56znqIgJfL2Q/ewZa7rN9R77b9RxaN96uaoLlHSqL7htkK8zluerewQZQLJnkqhofchS/ncG/gVRwYwJPrvvrShnx3JfVa677S2oz20H84Ee70SFH4o7O8unfPxHL6/5is9Znv6UcWaFTfTP/srbl7/83T+6vOvBh/wgfuf/9wvL8cMPLc9+ySuXw5VibZwAACAASURBVOu3zR2vRmTMwD1Z7n/Dzy4feNDKQI0U7Y4bGHe/4BXLk+/+qOXw4GD5vE972fLHX/WK5Zu+98eX17/lXY+Dck910oScbJdR8epnHkG4TYm5ISfQQ4cmiIV0+tmsNm5ZDqWSplXBb+DC2th5kOVhgPdsw4EFF0s8B0PW53Ne3+/tRp904cANtecsn6P2oR382Oyou4mUTPr69CakGKumzWi2CvAWPTQ2KLp3Bb6kEcsapU4+5P30NHv7MKydPTYH8fCQabICXnl4jdZqNaKJqz4hKhSp5VLCOtKqiahLt+STNd+zOqqY15NjHIBqtixgUDUEUeM9B9nq+hzrNkQFWGnUWgQAwvJa1aDqCIhqBPSAVz5fmbPmnwk8SMgiyqI4Xb2jhBUeXzPDyVqiIh1RZeJITkhUDMZVD/x6v6pdV0SFL7TuxnN6O3SnTe3vNkUYgipVMZTLfr1Re9kjZ5zMU1PrNjoi9NZlREVZrtwq84cTGFDlYE5g3lrppxkwuYIs5VxNAJUAdDXYgVKqTzqTdZeqlcEl43htcdptFHGIoeV3cR02v/WPlKVn76v0HXdDO7i1JpsZgcXC6IlY6QwZ9TBMmTVRwG6cCdJDqomNv9OgxgBTVyE+GF6ldlHf+6CXrbGsVeO4JTsJgDKzAw6Y5hfzFsY9wfUo61aU6hT+HtRtxcTXdMK+R8WoxvytERU6tXr970AbS5fAZpEjnTaPahO3z9/K7hys3YaoyEjSdSzW5cf8tiqzvZIOwpncrK9qEcKxZ8kkrnRBCK4L62DwY8A0nXdKBX+K9ZoAu6X6UchSQ6i0+90BjH3U4reXB22whveVo44mOiJs0vrkM9ZV8j8EYWbrrrImzQ0CVMs5z7mfgdoz3LpUcM8yfaVmsjoiVf02Jb1WahyjmREVyHxGJLxnVHgpCAAdNTrWNSL104osIMDT2iQpIX7/wcN/8IkK3XQ282X3z7ZnnLlj+bBnbsHJ2r9v/RuJppcb8p4EWTIVTVeRnR66z0G51NmRUVEiidXLQhHC6zM+H2Iqgyz9A33D7J3Sa9BAPRvf8fHJYvX7HZQ0281LJ6nJ7lz31kyGnBX1ZkNpxX7c2XdM53OChtQ0aUvsLMsJI4hlM6ongT2zAZ0RoctMcO8LYaVAGOzm/ow1D3ZyNZtk51kDH00lOkAOYa5uHh0thweHbFiNICqcb1naS7aA+rLpuio/I0LXon4dhLUsDGYOqNY6sh1g0wBoBpBnzyBiwn/DZ7QJEqBv9wfRAwBO84FsFfV5gN9sl7Zy4V7zn3ME0oz9JEuT8jijeC/LqHC/kP0gIb9YQ/N1rc+G5Filn5QFE8cZS0mFTukyKkTy2RyiJ4WVTAaJIBJH48JcnbustjIGvScQ2J7bsCePcreyVyen3pfC/m0NdEUKas9GWTEemb7WFqSjElsFL6nN2e17Dh43PWywM+P4nZG1RZGO/FuXueasVCktk1P0w4FFq6xoAd4m1ejzsexYw/a1LTG0uSxjzcZk0f8E+9UoWZtzpfvZc0WZfbAJrZ8HSMCIOu+eQ0G4OqOsP0vf2Bm4D84xYVPInujNGpyKHkSq7zPjK3xOPoDNnIcUxbqizJUCPKEHoKM19yIAnfyhX6yG55Cb/H3KfNGMLAOpDDK7vJ/RpTdDv0LQBmiIbvvbiAaTVZNbmwtrAK5sPtgSlDnJKe2iKkNeDo6kkRMZNfCLA4BtQemVGT+T34KdKHMiSFfD7jzjkz2QaIeYzkN/UsusYe9FJ16ZqeDHSHuyhRnEEomeSxRN7qHDGzyzlC3z54fyoL6f2YYFE9X3+dUMVMC41BdEfTVGPSpEHLs4PUFUYCbtMP6Y5929fNfX/OHlmU970rD6gnpDfNm3/q/L29/5XnRs9xS7gxa4mq9jfGJkxbve9PPL+9/zG5P6eyQrnv9xy1Pveb4fdHfedm35wA3rvzA3NLe49WPwK+m0g8GUkjSlcbpcWOSFNYc6PVrOTm4uRlTIGIGxCwMDPiGNPNaRRKriuEeFb/cuOkgOkdhWBgNFTVgALDDIoHDRo0ApinnWrDyowbpA0Wd0/iWh3wQ57EJSdh4ZxgZ1yvxAuJMZjBYZkkZv65NXQznH2pIzcfQOZUpYHuYkGw/6nJZf1AMGDaSsbBJS9Xx93Gh3zVfAwc333ijklyArGq9Hz1iEe2luWm0FrD1S0+2Z0IAOCr86woiuMFlIY7/T4w2osg1RYcRXplSinjJmqDxcB2aoOVgYHg3RhhkbOnX1kh4S0t4nDLb+e6NFaOZ+pMeUsdM/hyyrCh4WMCTA6rypA+2NnOn7hRjpmmnPNOtYXsMyibs08nFFokIOAbKOZECziaxuFYhajQQfR8W2y79Z6CMCowDRac2OjXR3UMtNGtnrwa8NzY5hIvO1AaTXV2TQS7/2mErvfOF3rRGat+ufDX9rP+Ee+nZxtKXcuOfgaBYCmP/ue1Ss9n0zfxu1ViEJtE9z7COiogoleu2wr4OM4ygfBnDJ97FIgPLMVCxBVGg6W9v7EqXKwSiiUcRYAs1q1N2W8wBIlIRLvSfqoefa5Nk03g8zdFDQ5Wr2meEBvRrSV4V1/ZMhqI0z3M89V0gpsbaHkPFYS0lmJpN0cj2nJfdVzudERTv6fsA6q/SAa8f+Epm85Y/Hun8MOGNvCYjy82sErtOxxtbse6iUgY6cxs4J87mVnTJzMnsqpNhSmvVYI9pA3mTU7IWSCo/9dEWbfqInw6lMBYd/Ta8/3rfz4cD9r7olSduqyRtjYCglU5n1n+Z+AJOXRGolKupuGt1kZWV3pCbsc3wrslsIMCpCVc60uwm0sxzgdJDS6yx0L0aRlw+K5aE4j9XvrtQq5BKZmfeomMhZrZsd7ta8pNaEu8M88GFxnpRNMrg1pOnCm/kKOLI5NjDJgRidRwTaAIqSbJTzRT/LbmufeyNZ6YBLyo7Ndp1jjWFTZnSoa6IavMasSi8FYlHh+/sAiBkRPzNneh+oThwAK9rzRad49kP0UsisFRGf1S63nwkn0G9U+sTujVJDADGjDrndkk1qI4K7KZPclosE2Gl1zq0HBfaGTVk2n0XfCm+obYA8yYbM3gdpYP/XXrN5QAmvg8gWEZHhzbqtkbg3WGVZlx0jUpD5LnBfUd3WD8OAdoH1MQ8sLaPgLiMS2vOVvQDYeFYBjyAsjMxJEtM9oVKOq+pNe19R9F5yk2tXfVnPTCARUiPVjWTqz3cROyM9ZziHZYA4+cJyLvq++0GUHWTRoBm7/beJyqbf4XgFyXStqfpcKCNXY1PGEp4NMqd+EjqH5QvrDJJ0G9mHviQov9WCxXrKsd1eDqDSQ6WdGegJZQSoLwOIdq/7v9g+RXUH9+N9jhwaob1BMs+IisFrHGRs5wjmVedGNMPmXl4RFVayjIRS7m9kD0mHqkdPnEUkMLwJPbMWEOSCrCDohAxg1FxALaLRtbJS3S9gwKPvRRt7BYO88THONL9/0bt2PW8i7+WrpK8zI0BguGdYsdy396gwHUmdIAIVjcfpsfe2F8dsesTGHeXEWb5oZBEqGwTXR8ZJZGR5s/Rk+/q9Jt2PgATIkBFBNnZk/4AgzfWA7qx2aSUVQ5o7w6raQMoi82bhzDLKdYPvYIEu3rM1Mo+IEXIPyY7pbSuqah+G1jLPcO4xvtEHoGZpPGKChcTvt4X0TJy/slPCxsL6KkNLZ9rEY4tAnieIijLTBk580suet3zLl3328qynP3lKVvz869+xfMvf/1fLm+9Vr4mhHrv0zbPT4+WBt/zy8pvvfMu0WZBt7mc896XLUz/ihZNalJfe5sPgC2E5b1X66bOfgR4VEfsZ/SG0HWQEwqp2nzRKMMgRw3fqhk9lVprYqDSLkSBkWHHNzlEbhVBtWJkEXcoY6cng0qUcEVpAUQGwrj9LlLiB6I3OOId0wKmx/D+hmHA+M+OifYbLQJE6NwEKOlg3qp/fwRFlriwDBKnaZjiYw5FrVgH8eoURIKtDG4RVTQVOEknTH0aXlD8vGBkWzQ1yXcFgI53Ozh/VN0zvLNMmq6GQ960CMAZMA4CMOvdYsdMzRKDU5QRQStnuCYvisA3JCA4lgZVeOFtoCMYeyThG+8Qv+CiKmA7ZK5eEEQGBE+EDcKj47/Lc3QBQqTbU2K1ya/9WSat+DK4FCNLCiIMxP3O0V6nKZe2nUGz9TvclZQb5PbU2RhLSMIz3fRJQ2SqGJy96N93pXLta6ku6KgEpASr9Pkl91oLcHmlfZaDx4EdPjij7KksVUIbVVu6xSdfpvs12SHCgMYwLeLC6JJ9BRpL73THn0NlNIzca49rDMjpFDOf1O2AuPsjSZLgGHR0XTtX2MKcge93IoQNXTKS9NHIMcHQAgobTtSIUk8j1xw0dUGZIa1EcAPAShIo8xb02bQSxCpxoXadEzYqr071hiS/9CNLXErn6kYNuTUkTbF/E+WwP8I4ju6uL08o5giJUaq5CjTozB99fjUfKKpsp5p5c76FLJ2rTPipOUAVecsvUPb+2b1wbb6j3f6tj66+JvyuCCW2er7W+yYgs6v7BGcDTxL8w6ocT6rQ1GPj9ztbbRrI6hz3Gzz1Wy4w0cys9VQ7v0L26CD/bXrr5wxnD0D9zfM8VxmBpN5TqAYobxOkYFK/a82pPIdK3tZmwTx1UsfJLBILsb/SiQ6SmN91V5DvJcaj5Lv2Fz99LoUbqBAbLacqNh5RirtQXI5368rzhrpQwiULUwzdZC5gnk5HQivt3Pki/UCgvNdk7A+bD666nYl2tO3Se9tjU4mn8opleWEd1Euzyfm5YT5WEUKa3bGc1Mo9143oZqSubanVf9duLKFPFtFHPpuFYhXM8/JU91NLZfm52wRcAXWo9+LncAyPrPy/zvWpcjW975D/LEBkhoIA5kwGU1IW9i74EJMdLNH7uoZKdFjKGeVK2ArJHUQrGQTQC94q4hopShLoibmGL56OpDwPuV0kK6UT7r4gM28v6t5fVYn9JB9jZa8Ej+WG8lFKW8uPzDFOwohbYQPFr169H0+8A1ZhRIcLGLh39ORw4xbqgZ5xFN2MNRFxk4Gj6RP4DAZdOAGRJo9QtmCYPyitlZZx0IR5h47CsHQt2c71GvSRg3YkOLzNlwC/K/HjE+HKxHB+xcTn3tPwgt3OZySnCCmV/0C9DvhRMw8QN3L/1nh3woQxcb3xJEgPSIVZ21/t2WPQ7fWsB5DbW22677sSTEyc+Zu6J0M19f8e+Zyf1VC3HamQJ+wr5Y5fzEGeHkWJsps0+FR6xzrGDcZPfjuAIbyzf2NyynZgZ6T4le7ScnS+H1w6cqAywm0EoEcEewbPMmnCCIdW4+ggoENHmGEGbavxtcm8kyrlnuKBJMj7PZsstiI5zpdM3HLPIkerhq6SdQPOYRxGSbMSsbDMnxziHyIITRqZeHSAxXG6p/xW8at+vzdLr+dS4e+o5xM3lJo3OWjbLtuurNCP2GQijyFKgHEJ/AzAPEo/ZEiLv/HcMIoI7y+BAZo+4P8kSa3Z9EA1oZN2XcVqd23yw1k4HsVYJFZFnvQmD9Sh92sLPxZZFCekFpdqM5I/sRNsgKQfy/9Z2Ba0eLUCcd5B9JznZL8X2COYcJLWX6Su+tnt28R3obK8ywt5VLn+56KlydgvZ/kRGRbtENoHPuutJyz95zX+13H3XncOeFTbRVv7pS1/zA8vb73/vb6EMkzULOVveaZkVD7wjQINeaOywfubzPm552nOez4NhbkDOjMbH9vth+W9JVNzA4zYNQpHCiw1vBkfOoZeH2sMB70qzKKDaY6B1CJTtoOZGKvHEZtCwUqJJj6URjl+ztQRINALn8V5tNAySxBSlpWRKMdvzeOSE1//koV0AqwBEOU43FCKys00LhULNk6EaAOtDvETDDUCB1TyMgIMKuqwcsfWc5SX0mYwcKHQbf2QgdA5CQ1TUscgRGZAtFLDptqrgEK4PZr6aCu1jj+SgAJClIa/d9PxCNUw1BD1nYfW3mfvuCRrDsxuSDBnNowzQi7ML3z/Zd4Rj4O+TJOPNgBxwO3VERbGNA5xUHxjEucSIm+iFmPB8IDnCMITgUCGqAwb56CXAPh59K7C9lq5KfF7P7T1LSL75Ie8pvb5r3BDy2VAkyWBQ8Fn76EZFcibUUh2LnqjIba/nrqAlHXq6zkEYNdjOQD478rWNxCjETF32DQdRc4cByOS7qAJxHSDvzga1VE9QSH+Zo4JoHESe2TXVAFC6vjecmyFXeZBeYGaVrGYDg1JdwrnVS3V5qzEuRwHbohBG8SM5RnSgwmmSPsbn+cwADfr5jEGEUyagoV0UIwVF3Aeg4o0Fq4EL+b0qUaFrNHrGb6/a92s5A1fQvg+ndnZ2jvf2LREVEzAJs9vfH0BPP5v6O6cvz6jpI2zYJ5s+6ucXDji1TSHtckzteD80RAUAvZZElYyv1xrab7ymo8wK/77qE2tfSOYrKVgncmPk9dUXQ2BUzSRFltwWr3puV31XfjqejXp4dlLIaza/o7P7WyUq0mHW060Mh+FD9zZkfin3UR7rzEqijYqodYA1ERXM0nw6JxoQQNJW7N/RoGbzKodewEwqdAU9pI6GvK5lNna9ycHgRg5wsIF3Q1TMRMYnB7Xgx6+BLq37qMsMyNIOKjtppMCsZvz4jrN9igjtnajdbvaJl7DwEhzZPLUV/Ykeny+SFJ3/V9fyKG8F06xV9uRByjlcSMNNJw4CHWCBOCi5gWQSED07K/pSMwBZRRCyBCUzL6CzW5JZJVL0FE4LOUbFczxsJZWBgX0s+zfKw5itHKQHbQwDOC1rhQB/PEPoE8q/bwIsVox/MNs6cwQEGqFgwLn9FNkByFZXhrsB8MiesDJbyHIQCGxr3TfLDbvI/OOjIwfxbr/9dhI6VoJY/mqWpZLP6PvQAk0cAEfzWicxlAHA81VBajXbN85YzwbM7GN8h+V92O/CffadXb+2QH2TERE32RgbmRmeNbSzLNevX/esBC9ho+bd3ttlz0sRKwMJp2pbZnL3QFiHmgyzzJ35JAOS03v2+BywasDOjpf3sr9rJoX0iMicKGfJPWhEgZUG814GpX8MegdYBQXKDIPYMI+1ukX21HLZqZUkWK6vgsqxDsz+MTnyLI5TBFLWLBGUMaPuYLlQI+jyjEyLw3S1kWeqoiCd7ftM2U+FRAGxyP3kVSOQuWL6zx7Znl29LfSZyerhtcPAdG7evOnraGSIzZee09ffSj/xvvWZYy6qPqIORbURZJPUrBvoT5HJKAfmPoVnNrB8N8Fq4QDImMKFUZYIv7FxWqaZ95YovocTjb6f9pdzlsmyPd1kKax8jrHGNFmyLAebY9sP6oPqK0f8QPcWuasMSgDnCDj1Rujsc+QkIDP4wieu54hlaTgojzJfruMqCb/Jp58QFTaXdn97Btg14+Ctur7CBqpPZfrBXpaZ5vuTOtx3Uke89WRFPcOnNhrPD99/9KGR2WPZcIfMeAOJ6qSFk0YMNHEZzUDLEVEhIknP+URGRZF7K4WDDb+/vPxFz16+7S/8oeU5dz9lTFZcXCxvetu7l2/4nh+7pZ4RVu/w+rWD5eEbR6783/3WX1ne+xtvmvSsAMj+9I/6mOXpz33JMEp9Zst+eLxPrRp1ai8p/fR0EhXVWiWYJCbSNzUtWRy8WaPNFDEARAFBdRYTFPLDhemS9o2MCiKMEQaJuRNXJSoIxTRgczWTe6KC0RDnZ66c3Mjz6AcBoZ0kCGcJppTmQANqqLmTSB6MKQ2wtXQVCMY/XANSI4nM52rWZ/RVhJ3h2nQGdRjh6/hMZI0MPXvPDh2w/oOMFzrAzUq7jBSP5wqbKcEhMfEtCFlFs467vQWBQD5zZAj5I8L5qvfB03MuO4B9CmwMnmm1ZrE8jHKncSgDx0TCU1B1MNcUyFJfuCEWmFFRgTX6gzmiaixHneA1UeHjMEegwEBBPnFfViPFvhfp8t3z9x2DtgKWdI2OGDLHxh0oGkEiHq1BoRn90QRxAkbFPuN6t+uyzqhwqaBRraGEk8aLKaKtJ6QwBElJ/9RdBkpgM61UNRkVNGbrlWYgRkxfu/makj8BOpXvBCwWehzjwZZN0Mx1O9/vHdpqeMvgU8TgcLtvICoAhrTln0CKi6gAMVUdh4hMFpAoA3YiU/lsa8kU+JuPnnoSE8PfVFA2gIQSPMc0b5cIGaTRTpsD05EcItCOBxHz61evr1L3zUF+nQlxtQtGaU2zKSb3Hi9o0RvtMzCGtfuV5lQHaP14O6KiAqjbIdfDgU/mtyU0e0ej1+0jYuNKOo87btP50pMf6q8Esrqdz9Vax46+ygkGWZcuD5ukZlyNZHP7ad74TT+PqPtFToxLBOEy/ZNtM/9XnI1GzLb67WVnkuxGP7RrwsJ69PNLjUeSvUigzSEibE5qQICXYUCdZgBVsFPtfZWfUDS5St5B/WFsOOquoiO6bJtGZts19MuynOTovLt0bRW1WQm2mbQFUVG/sJm06MuV1DFGoAEzoWHfXY2omA6VoJVFYaq2tvrz1JiRsFuYIXCVLdlEDJdzGmdYZthvuxkEwkhHxd+zQSlzl7YoMux7ixI/hkWSr6r3/N99RgUbSassrpcw8Whf+a3UoxQwzz6ovmm1kSpYGEFqICrS/6LfIqKC5ZN9Lo0M8Eh+ZsRUGrk8lj+GHrHek+/VGXCQj3Nl17ZIcf9be5q15k12sqSVRUTD7/CoYZXX7exwDSHLvrBML3+nCHqpBJtjs9Hlj2TUOOYHZV/qvkDgo/dGGdy7ZpHo91YvH+XNcs5rJLirEWYk2DMrQjtKvsD5zaxmzwLB3hfRoybj6zOefQJ2kTmips0CbLEOa02VpaKgP13Hcl85waV+S9Svbudy8u1qvkbS06dnnlFxcnrmJYCciDGQuuvZKv2EtW0xEawXy+xRiaicF4bQ2WOUDxAbOAK8bDsbtmPtsgz4xQJiCkddnY+wKEJmBfIbwXbj5o3sGUlw34Bi+46D4OyLoibO56eQXQWtBTHITBgRAYbrPPLIjeXgEBkzekb3YZg91YD8PEMU6T8/RlQKjg25Dbgn9mF7XeuGMtw4Z7VfNd9+7no/VhINcS7jDLHf2r45unkzgoF9XMzKQa8YkDfQfwOcqQTd6FncCidRhbJQy3KwZ6QISDjbAx4AICyOeABkHvITskIdhd5UIBc1nhlRkdlHIEi9DFY5w0dzXm3y6guEjO0gI0KEUCm4tzozhAH5cvl9Zd+kbsB1MtDMAkv9yRufs853+ffETrJrWqlGu4YCRTDfpteM2IWMeEaV0CpmWdhYkP2TAc3Vaom9XrbcE0QFp9F6Rtz3+p9Z9g5uW+554cuXvf3D5aPuedrynV/9ny8v/Mhn1CoWISymxO574P3LV/6t/+NKZMXhwd7yJz7rE5ZXf8pLvDn3W+970Bmvd735F5bffOfbgl1shRwG+10f9ZLl6R/5u5bdvf2Z3vkwfF+oCKOUqMjcsBr1qJgQFTw/Y5NKoVhTKbzaqFH7XJt/pnBqaaNQssijaJWKXXsI3mSzufoDOPcVeJYDVFV0Cz5FOnppFO7p8EoB5oEbitT1VzbjiVTJqAHNg9tvoyaiawcvDKEYWikePjEae9nW3zjw7cASEFRLECQ4lKYCjuy8jQ4eRM+bokTkAQ4lMOYJHOaQ12l0uYTjo2L+aJi3avRX2avTlPMwcmEriFNmzA2TrGOuKJ7GGcNJBFmnc94brNsoinp4puQxrZNZST0Qpcid6vhiHJlllCAg5CmyXWiQwjDIOakGb12z4TM0U5mlnxBBgQZqM4yzke5+gTeAG3HL7jeIIoCRjuc0EMuMUshyNBLbsE/mGRV1VnJH1Gfbhqhw+aiEUhgwkp76X+pJEmUQM927NeabOemdhsHCtcsGHSqZTflojSxcpjx7c90iPyQr5PC5E8PSbXJIFQ0ZDku5th6xykfo/rIM0hTKqjB4ZHdHZzUjd/KGUL9qssh9OpKlmOFicPdT2IpQNnnsVw+P1TR4CL+gAUmoOGyvwsWsKASeNIGYVn/dElHBJoS9TlyD19TxE5S/OgITccDbdHT7++nvDw5RIZKc59oVS0Juo7O1J6fzwD2LPbB2WkYn0cb7bpDJ3ikT2BDFKuOMoj708axHMAKAfAlnKHghKuR0T0vGbDupW37Pxpr9tSBFsMHGF/C3aYcN9+qW9w2RHunWUGADAGB0/cuICq2S65HNRMVs+LO1k6aB/c2tyhQZ2Bog+aMpLCP17T0DvRT1rGyWUM/UeZNlgEqYPvfQAqknRAGPEkRc6ehNa1l18mC9+p9CsjaUfqr7SC5UBwRKZqIRp96IKNQx0D59jNnkys8oZ5y9ZaRUZn8Wf2dQJkj3nJlKqquPRaHtq/JEV9hDcTZ0Y55uYMqN2yiMTg5Ab3LfCjTW8yd08iCi3ZvH7sOn8Yhbq5nukfW9/cOIczYYt+vXPiyQc5RnSvIOIHBzHlCve58JB5ySCFQJncxekE2ts1l7KTYwrl0Wr+41A7iQGQHfzEBZ71+gxsLMnjKg1wlJ8xMVyUuSAn4tGm7L3xvtZ/vcIrxjv/MMtmvay7IEbDwoBYXzCP4ISFH7p4F0KrMljECA/3qfQv/bnHmE/MHhYv0zrh1eQ/WG0ntEvQIiS40ApIBw6+XyyI1HXAayx0NWiAAoDcLEo5sPD6L/QLWTvbzXXpblSnC19r5bay/vRWDgL0vUaH4jU6fYFuZn+/NZuZ2i23Q+2jzEZ75n00/qTQDsCyinAGR5FsQaF7MBQVMEQgVGM8/NrnJuVQCWXUb5I7AAeiNLEnt5Ja/FO+5RoX2kkmHy8ZoeO2y8rHJO+/sHy7kyyEQS0ucVfiRCDWoMD2Xv2Xo//PDD/t8z64NB0le+kWXQ1ECo6DMzAc4rUC3Zbfq9iAij/FcbzOZcIL29j3liKWpmO/n7+elS1gAAIABJREFUrGRg82tZUUdHR8vhoZGQ0Fveu8LJDWTGDO08nslhJ1Wx5Nxl/01mgkRgI+au2hK2XnrPnsOeWaWSkOjUYkGBb5T5EKii8lAuU8yK8sBnz6wYBw30NrH0kM8H+3xUf3dymTY7RSXsVbpd2QvWu8YziLS3svQTSg8nAahpbf288QEWNq7ZaJ4ZBKIpMnoYFBTYFO+PjJNdZH8pS7CpDwMDAmdFORmfKP2ECIH73vRzy0Pveocrqjuf9qzlWS/+xOXw2jUnKb71z37O8jEfffc0s+Id73yf96z4mV9+26VloCyT4os+75XLl/0Xn7LYv99874PLX/offmR549ve7c7Ng29/w/Ket//ahsyKveWpz37+cvfzXz7dCFe1yX7nf/+qRMUj6ewOECYx5FJIzcYUqkumtgKomCcYLjIovYZflBqXUdY62qpANSIqLnPA7dpJerRAYDXGecqSRbYIhX1EbFBJy//y++kZWa/WIQJGPzTRA16im0Cyg/swZnGgl7EQ8MC1CTBOo11H0tYBnDwsqkGS/mOhgGiY+ookukdFBwfOoxSUrnt+4aRFRl3ImRlAMy1qOnyamcMUuR4x6DH00wOL65kpGRXdhw548/ouozIcGuAnf0Q3JPu2dA7DTA6rsaSDw8BeNahTGrQaToGLyFJIATaXMmjaR9XR3kRU+PeIX2VWCedUW44Nr+KJizzAkCIgx2yK6b6r89wv8AaiwudJvx38zu5ua4aoFO4kRiHRFRqS4a5x/MKj0k8VPOlkrAMg9ekoo8LVQcct2jy31bHq9QElNdGYBazkrur0RBsl09maUCmruc8eDhkR0yMh7bgmZpXPn1J9c5kyYwzGEebZdDvkUfqBv+gM/hVREX1XTB/B0LLvWNRfdbKq0ybfXfo35iH2cftEkFs9c5Ys6FVyu2+bFRlOUbZuzz4p2iNI7T/v20T4OBBZWMeky48BrjyH+mGgaXyraLvzrvzE9dmk++zWREVuLi1wM6hHlahgtFOuxG8vUaEH7YkKf/8SkHolQI1Mtp+OnTKTjbb3h0ppCRjq73GZnbQW6p3lnOJTowPjLBntgvmBPlYrk3dNz8POABjm5YlYw3dkSGzSaNMbz8a6gbiJa5XvbALtNz50OV+wD3lA+496e2d8lzlRAcAoZVSXB5ARARC0OxUxGQCDynwySlsjCxu3Rv6u1NBkRqp9GcAJR9L5GDoZ+6VotNnoNqzJbN9TLwYHSSYLcSWigvs6Qb32TFD0uq9kGfgmu3A8rHEQiEAmgT5e9slLbaDOvWygKj6z8pxToqIYLK0/UGSpniEb9Fw00669RTboRreHrZxL9G27TGWwlFPztQISD8429SfwCGtFIhMcw7wmYWhBWucElH1HckK0tgH6qcQmgSHox9J/hr6uwESRQfY9by7Lptw+NfEsGEi6P/x7AxGo6Gq7hiLPjQwAIYLyJdbXwMrgmKFgJY5B/iJgy2uek1hQaaLZGWKldqIZr/v5kHknKljOBVkjCM/Ys8bLqj/vvqT161D0tPQdysbM9otAW6v9789zbg15jRA5KfqyBC0G4YUod0WL+/WjjHPW2I9zxsopMYjNe3Jcux6ZCJgP6GrIEvwijAWERhBlQ/GFzsA8sUwd683bWoeu6jao24iWvUCSzb5nc+VZKKdWXsdK9pz60FyGisKrwW5hq7C3jZOr1jPEe9LA7wzAWiBs9ZscxDXSxIg7EG827tMTi7oHmeREhY/B5gIZFX6PRl/Tl/QSXNBfGaSK8XtAnGXseN8Y9WmAHZClf0EYevky0GGwF/ib6vdK9q30k5dF4/+CYLA+J9HHAmvhOl298Lr1DNu+9PPwEsUq72WAMvVG1R3S34GdMQDNn9GD8Gx+TQ+iL4ui5l3GDlHCyuXZm6gjC0mVLlodwgH3tkqvs8u6xDi9YTz7BbHxtAJfXb6ZnWVzf3R07GSejdP2gM0h/PPMwPNnrvIkfKP0QLHnNtLdq7GIWZgc3DXzryFFWBYMc4UxAfif2CQcp01JEtHmqzE7h02vq/z5rLJ/by2ZVrX3NkSFzons64N+ICkXad9Lp4gIRr+d9kxQt8fkMzt84fFNVFy4gnzgzb+EhtYEKuxQevIznrM88wUfvxxcu7684CPuWv67P/cHl5c8/1kbyYqv/+4fXX7xjfc1JVmqfrBST5/7+166fO0Xfvpy7fCALNfF8o53vW/52v/+ny+/+pZ3+mH87rf92vK+e9+02KE2Cv014XjqPc9fnvHRv9uV/CgC7TIz6bH1OTfq1qWfjKjgq/YX6JWaWyhg+AB8ZDPRJg2TclEuGhsy6/XhUAAwDg1VzWPfwAOFs9kBz5rkuJ6cCzuVWfqJytBlVwamMirIZkOZYPShsP0E0ygVMVKZTKVH4of+u8aAKOzAgKjQXDVKbyp0LSAFOwcGVSUo8C6/G4Y3y7pUR7KbfUTBpIFXz7rh/NfnrOl0q8N+/EBS1oqOSXCxOvMt1zPewzXCoC60DCk4IMqYkfG3Alg7LdKD/UOwamLY4JzDAeo1RsuhHD0ZZKjGkHnoi4CK0jJMBfaavm4WRfRPzVRKI5hARTWEdQ86qc16MnhA6+ERUIw4mvFovo2kOkKHtNHn/apXM2IF0ZQ9qblTM0CALrifRxrMDBvu01ZWa+mniS4oDqouPSMqPFWT+03kKHtS4nG77BbF2Ne50Jo1EEg81MTYKs5r8/gV/KHhj3VMPe36IK6vmVzvyVa+Aa77vom0d+gHGEmQ7Z6oCMO+AXEYMROPJgcG+xMjsv2ZzbRReqpiwWrcV9LkiyCMRKIfi5zu3oavfZiqcI2uGUQFG1SG82XPwJR97A2dxXSqJmUCAojuluNSoqI9OPudGLYOjrvxhvmdS1Rolktd8IkiujpA2AGMTbTU9OAFuFD6NvjcXZmomJWboeoooDZ0oIgKRdhW8LnRKPOBX/JJo8dd76OZ5FwL3fKtVj+0/WhAmkW/2lZGqT+WotpmAPUg2IZ4qCOYfD+c+DDMMJBthjOcmUpU0OlMG2Z1Ck4uMbl7VBospS0VHCTwJKI8UX7Ealwrk8L1Ls/dkOVy1irTYjSo2Xy4dm5sbammIrsxtwrpaa+mWfGhDW5kEc4o14KzCSVttiEqwlAZ6Es/JeNRE+xrontCDwBgLpH183DOyYaZZKsWoBylTTAmAy+yzG47/BlRsUGbrZ6fZn/7E8ruRtkvugK+A3XHZH8FsRTlTyfGHEciwGy+dcc6FSWOEAUskBK9trL/h2desExLb9sHUbHSySA63Juq4GDJcAaQzaxgA6j3kMFQz9sqrXg/A8vctprMnz8Py7TI/vIodLgFDmh6VLbhHWqqy8a80ajV+1OcL7veLDkmOsaHqPSDKPsa0b++vMjkz2fJPegZXKUMGkgNIyrUrJzA9CBbqVO3K9G1ZwRAij4ADtryJeLAymAdHR/5GIywuG7kw3LhPSjMnlQwXq4tykBZE24rt+N6nsIu29OBWPYssXmxMUhPZPmgVoZVdsrWwO5roK73XWCFgrQl8ACGZVkNf7u3ETJG0HjTb2Yv2BiRBYCI9uinIRe/6i1Fd1GdwU5HfwMnO3ke4Ll01kMX+f6lewBClhn8TnJZoHLxI2i3OzRkTdM9K6nZpSEj0pOynzwoyZ7p5CRKXNn95StLrs9OjNS0/hwgOlA2GQHTlQBADxjYjN5gnmtp3zk9z74+7lPUDJIoQVfK/dDOq0/i17FqE/y9Ty31cqw8IQsngVRijUB/C3SjT4MIOPRFOHNyQmRFkkloBm5+sMmFVYcR9tbY7j1JMVD8fo6ygbo9i82rZN71xwKd4KXF3IZAHx4B+5bZZPvJxu5knREO1OEVM5oRFW76sAeSsED4jiDjRq+Yj45AFtGNsnqoBOJllWblF4s/Vkku9eD1/ivSzyKOOafqDQPMpj0Jt7GSJZcq1VZLZOmMCntHmBEDAJ2sI9kpu7QtZO8aqw2YeDwTFXYwvOvNr1ved9+vrzMYdpbljqfcvTz7Ja9cDg+vL8+8687lO77q85eXvfDZTSPmehC99/2PLF/33T+6/D+ve+uqBropsD/y+1++fM0Xfrr3pugNlLe/873Ln/v2H1recu97HLR68Dd+fXn3W1/XseH5KxPCJ9/9vOWeF72CymWzYTQ37h4LnwgcIVBCZ3pe+imJimygnSmDPlPFGUTaGqJfZdjq0GgBg7ZMk43KFR671+OgzhrkXoNQB4QbBQDV/VghMIgDBq+SK7AsO8YK4xCzx0VambIayEiWAzjk0A3I0sgN1ifvwahsf/YutUrqKqcal6TfgajEmYwpOrR7BipSKEV8x5003iuu5teVF1j8qhjLumlrKkGU1GpHZsAEZ4QHGZ5Fqa4EFEvDOxg4xTkoAPMM+IpUN8qTfS/mqanJ2pI8ayS8MR+aDdnLXyxK+ZYyKmoKcT0kNN+aiijj5dOQzHUjfzGjuFKuFfdOMXyaKS7Npmo0jLIskmiqxOD/z967xfqeX/Vhv33O3uecuXgGz3hsjy+AIbYhGEgKpoUALSIS4KBUahVVqtRUfapU9SEPbZSnqqpURVEfquYl6kNKXqpIjVS1FClVSatCS7EhFy4JBrs1xOA7xjP2zJyz79Van89nrfW9/fZ/jyfBw8yWjs7e///v8r2stb5rrc+61IgvhYU1b42ztK5H/b3uUf289uGFQpm1Edf+uDqjVy8fpWiCPKg8MxJJHB/RDozGwMEP5wcMqVWvTAAViPzoov+bdM5Ce5NptbIQKsqcDrQfGQkO8unrzHfr1Tjd5muZxnTuuUADEd8dm2NxFAUtB3DZOmpDHoZszfJiMlBdkSNoEbI/DPN2LKUGSZlElTq2zkUOyRPli5QAm96j/afoaGRrKxeT9+r2rfhgeK5GO5HdvczEdiKS0C6H8ilwQo5N9PgJhpyUZ8OhcZO6q7cTrDvaz8CYUQ74N0+TcIyAqIdbrqJrQSxKVwu8v2eUjXlWl2fwV0W5jaegZGYhRojeV+8o7mdXtiQE9q4nDg8I/WTOmrf4dK4btLydj7NoRewR7/Px10kkSL8EnobRKcKdjuJiZHO2u/NZU+x6bg0Vx1TMkQBHlvGpO89KwEN9WqWn4O9yeENfrAV+6CxUBiy/l7k5O/exyiWTtpimcEzuLEsZbHE58pxIHhj3qGhozblTZQeZoCFYgkq1DA2Uc4qVbrDFAe76Fx3rI93lRILmqwLQosfjgnAIfnZwPIjk7c4A6lR1Zr2kaJuq53pcM4raI1vddjDnZSvK/G2xBNr1PA0lrdszHPIwQWY8xAO0mLFRV7XRpeI+oxNR4ppepBOsgFbYAJkdOvLcjDtaeQ5nd3JOxDRM6Di+64ccQW98dpO5Tt20R9V3AFwvw0Rn8wFiF2AQdyRnzFrivj2jzPHrGRjgZh0b6JpDWIEX7ohzh2eLN1e54BkBF4gWl+0AisBuuNOechm9B2C0VZvY99DNpfzO77VoXo/ol77Qnoa1RFB//sD5jOxNNY82+WSR2RhA9gtwGsVg/T8DZjzT++oCkc0W3btZiSaUlkGEt/HTNcrP3L/vJYAjW5TBeEGfntVkTW1PmWGbAIKeBcen3p8gR7P//AN6OvQA7aHLEq/LfzdKD3kmDB2leo6VqRJI4OeJgwMESehzcH5WoI1HqeMeBMZg9yvf2bzvHlvJFtP3DCRQ7wQEWiZfEjX2QwSlaSKIpep42huxKvlLTnjtqehT47FxO1BDkKrKqATXSUsE6BDQhl4lAJBQ6srWUYCT98Fxx0ktbyZACnZgBf2iHJDkhJKtqaJ4GTIPCkSPHfgKMK4ovWSOcvVYkM3nPNv1DWMptQS/YBuGQ509rvz7aEKc/R+UFaJ9sDGodJE+Ex/l3rcCMI4tHf+lJ0O9EjTDTSXQ6EviAblaWzjldW6g94bJAnO4H0ffEfAsM9bvHgOocZAJK+n/Rw8MjKKhRAKT8tWp7KwaTqtHi8pN+Z56Ng99YjpTSat4v5WBYyaF+/OSj+Wj01Ej2pQupfnqDBUtQjaug3c0TwDKWEc9G5lrsIUcsJA+0ylp7h/wHhCcI2Ug6J7lr7iyklEwy0Cz8IVAXlPqLw/1VN86xZTZP5Xm7OWS8b0OYO8xOx7vpe+CoBqAxhwChpmS9A3bo8KI/A8//fHtj/7gdxrkpu7W8cn97d1/+oe2x556xhfxve94q5eB+p4PvGuaWWGL+6WvvLT9Z3/r72+//Ju/F4e1MdC/+a9/aPtP//KPbU8+fn9KEC8/PNv++s/8g+1nf8HACQjUr3zuU9uX//lvbdY/Y/ZjhPDMuz+wPfst31kadi7p7XX8RZz2YKoDgQonftXRbxT+Tgn0Ekh8R3BL5RosnQ6kcCBS8YBbEdcLrYUQQY3GTKkD4iwwo9qIYFQ5HC1s5XI7vzj1epY2XVOC/dC3RjjO6bjehWkocBRCjoxT6Y1wgC4jggfwQBSdktKsVAEUsA+6u6o1jWUbkQVC/HEiSYtO8CMNq1FBb51OxeD0R616f8xxFddd2EzIlEI4kNG0DQcaFFLVrNQ61nWCAJbyZ4TFiBsi6GqK1akGsVdpY6UC2frV2jVIAZ6frzAjHfQZYQGB72UoWCdQBn3SzmhaYT/mh63Pv9nmPMDiMFcJsD6SozEIG3V46lxMPxbesTKAZ8JNtl457uKyneCnhA5jjhHiWV5T6HAWHrlnrfLWdi7gYy8PdQRl2AwSi0ix/eubzPnexGGe9JhGO4wyKHWjoTJE2A9zwJxBI5h2jdrQ/aHErLwFjfYx4+2qPPEtSuMujmXuvo8j/Qcpd0HlaRxHKix5uzZT6xWilpdWvJdyq/dvDXQ5YU7fIcprHhukJSpo3T1Jet14ggfm9VxXcmGZUcEbXHmmoaAom8bIcaDZrwjAOedd5Fhy2CIwX/Np5+U7t2zAfbPrp90TnI/9j5r0zuTyVH4UA6I3TkZHoBw9pWlru9GzV0STYH0pmby4WIy4+3X/5Wys4KOb1/VWL5pcXA2jOJuY4t7vg/4W9jnKrX68tZ722Ovr9rNb3TGXW0ngOpswgz0AHPKy6jDS2WCSB6Agoz2upXQLNbXvqSUn3rj7qad182DG4e5R1dwSUmJKFqvnwPCe92KbPUiRzeH46MCH/h7ILakPM4N3fItPi462OId3+MGNbDbMRZkZc9opa84ZfUb9B7MPJWuIrVW1h/q570ajA/ikbgAfGQVvjg1G5Ue5otJHymdDnbh3GuxNCsPJ0kF1XWSnADPjmXETVMt9dccKHcMeJxt7ZfpSZoMetuDcq648UQYqoezLbX5WTbNXPGH0lNmt0A3cQczeWTPd2x1yLDOjkjOwXyhDoGSEQ7/K3pStoDQ4nBEBDoBAulPVlllKR27EAdizjAdcL6e4PUdNoiEM+WbqGeaQhpMsdYbo01aa6crRekXb/J5H/FsGjpWTgX3mwXsbG5YfHbl97HozAQ84yRGEqB4Bitp3/r2w6Gk4KoGRt7tl64J5wU5UaR0LA2wyQ3o5EhE1qZMCcaw/0NmVuSunuV3h8/K+mTWDHDRvPgXLrjDnvvgJzk2j1xCC4A/qL+4892pNKJVkS2/gBPrkYZMs28EafAvYkLMT40lA1p2QpTlxOGvTm4sn0lkrZ7CDRZZNwVJJM94yOjj3aHKUUKu2uIAHoy3QAYJp4LDN80VZPynTW8ROctaeIX8OMnlUbWIcmc1XEfd2jwFdWicBSJqb9zfxSijjT6/btb4bgECeCeVZmOizUrHSaq9Lz5e+4BkpBLmM7tHzBUCkfE7TNSed2D4pkt/3nMG72kvxsveloCy2PUH/A2R82I+N3+avfVJEv12D88bsUutngKBb530pfG4CFPA/2DGECBo4e/YYAL2QJRLplGM2Bsg2VkmJ4ODkc7sUPROOcrzKiOsWK7OMMusE9vUoM6abrw8VwHoNEBVlyMG3tRxdA+CXEk/2GNG9ys8ZL9gaQiZYJsu6r1SUnVIvDgIGqyBkgUv2faMnLQ620U+Bia9b8bWZE4OI5AdvUKDienv08le3T//6L7Bx9WgAGeO++7t/eHv8KWuknYbI4w/ubX/zr/5b2/d/53uXmRUPT8+2v/Y3f277xX/yKSegH//w+7f/4j/6yPbEg3sDPbgT+upq+1t/75e2v/O//Mp27nUleXxcXW0vfOH3ti9+6tdL08q6lUfb8cm97b3f/SPb/See3uWP1/eXWhAe/DcAFR959mEYfQ1QsVoE9/mFBSjWKKZHMikEVlXEITlC8WaEg5pYS7Cb0JQy4geIO62QAoWSNLW+mx2admif4cAmQu2RF0xVrEqMR7j6AQJ7yf9jE1+hvY2jau4rItElhh0GdfF+DWcHVyuMbJdK7ULru1BOO2m0cqTkZfWBo7E9bVLeJTHUZ9l6ubAv6LlSUi3KxpVYCn8oB9VoycWTIlD123DGDHZrUc6p+CHKUnh2HsY6jKAk9IBL6xTpSbrVtWl8REmyahzlAFfO/6Nt3kQsri9zxB4m4FcNyz4SIZwxqVfjMGvRj5ha/fy2QIWv72QvwoAavoQqm7RPgh4O5vLQRfDEyhE4nwPqe3oGlSnfDnodIR3aDfNe+bgBqKAS6O/qQYTCzzGLXaACGzUFKuSUkIHcs/+BQAUuS9p2A4RARaHUSHGm+jPQTBrnKrFUHTf7vKNnNidsI3oUDdeOFfxamWEgOMhkZuxVARkGR92T/JB8QdHMFcK7KlDRyo4qP5KJ5vzejzQiKHmGKIpxu5PANNY4wbvKGknzKXtaGTU/fCA5Vm6d+cE9OvXLbGY1vmcZFaVh+8zZWIFXHwWNhqXzn7pBUIgMqOXU2gguyPyddRhJa6XVTOVnvfhfNlChd9u+VcOv57tXB1QkTzZMc+PqNCuyuHqx6MVZWnlutX2VviNwQ+cejk/qb9TBGjLIP+REgq6R886/GwlWA9MG5cxVx8Ws57oHzsfZz+o5cihITt5Md21D1z5Lon+3j6jRJW5mEnOIYD+Sk6W7zebmdcPp9FGZyssLlDDCvGfvPFyeYVVLuvGELPsjOh1ZdfLjWZCPwnUq1+PR22yCCRAAGd/VO6ZZ3bxneEt/P1YGT8F3ezTerjz0HuhiaTvgAcqqCD2TAPrh7E591XVxlc7EueoFkFaRLAvmPnR9ND6bhek34mWf301ABcvaCLAxG89K53gkcbVB/ZBqwZxKAxZFDKeY9KEsiZLAAveTtnbVIZ1W3SHoM4i1QpkS9ldxZ9nIE+bf8OsUWc2a+HKuGo9Fc1tuhzeuZgS36+YWDe819BHh7mcJo+3N+WdjMsep3WMOU/sdJWlOtrNzlEOy+42GHNzoSrRoL+VUR1UD9jc0x2w5o8dQKwy6dTTOZCauU5Nks+trtkIt0Qrax34aoHB2eor9lrPRtpu9FyoAVMEu20YHQFhFwLJUlPGN52JNTCbAOYkgT9fDGexjf8PxrIhs7G89y1sdDs5XldLRtTXroOdX+GtSFllTYqNXK9ll763ZOgLZDGDBnrGME/uVQFmj7KFYVONfgUHmU7Hy75Lvw9nikwUpC9wz2QC6sewfZBLobDAa6+lJzxz1Vayd0bONw8ogyfHu76IzR+uVtg2eqHW36+CYBy8kOIHMPOcflp/t54cyfMYn2VDa9bMZUFHeiR4cAPGU3aPz3fgNlQsyy8IbKCsINHwrzBoMhyfOntY+zjPUxukAFQOQ0dQd66demXDSIzvFegDDv9KdIQxItWtrmSeTadI1hnUq50HwmMomMZPp0LNH55n3J2HWutG1Zcbl+VB0hwVQYTLCaNf6WSALXvyGnjCznwGoUJDzyofBvjVfP1Cx0BlDKZiMtprUb8zST9fbZ/7ZR7eXvvK5iVGIBrzv+FPftz313HuGCF5zLr7ruae2v/Yf/Pj2I3/225dgxZdeeGn7u//rP3YZ95d/+sPbU08+GLIwjD8N1Pjb/9PHtp/52V9h+lSnrF1dbS9+8dPbF3/3N7arWWbF0dH2/Ae/f3v6be+dh5Afyj3f0NeRyCNdV4qYobMX27XVxrs8364uTrfL80fbR972sIkmcP14bV8xOFknWTpS0naEQuRRMJGW2ZsnapiESBUTCFZTMCJVXDHwxKeIe1ANOQgu1NqVgLlzbM5KO0AR+STnlH2PqIESbRHOE0zSD7sKVDROsDg25zBn7+A5AKRoSKcKFxtNNcAZ/aPDNJCV8oBi0jSKblOWiU5xWPUzR/QeMdteIirDfpQqhzTgdGoiSgtOoz2gAsoBIgMc0Y7DvBfMc6DCaTOiq2Q45PhvC1TIiImoNe5HNIYrfSUEnL1qoMI1kxwr1Wn/oAIVoVAhFCAUsBkw0QIELXixB1LMDEU0iG5LnGG0tbdAb0yloMjxzZwQ5bP9Eu03SlbNS2mnXqf67h2P9DLDynmamWH5sH2gokCvLDsyuoGbWR0CVNQoOA4E67sDNR4AVNRIsOby6MqTzo0Wder2hQYdhiZ+Gw32+o52c5L/pDs31zL1GMbETnbP5AVu6wTAUN9aeb57rgIktNavFVABBuUqtSvgBnIVOhEtWCjKRVtbiqVKOxmNenL6dmpUTu4dOA71ZGc/a77X4YK7xp4VLX2ghES/9m1U/pJZuwikJVDRVEgsc1yCD68voOI2DrnqNNlzTrQniICajIxPB/J4puZ4ZjJ6spsHXnaj0HaCKyM/4LmuJ5D1pkAFHwenpYJy+pHopZX29XJ6gYfB16jSUWYuiq4tgiT2FOn5qs36Iu3T0asAKvYYd0YG1ZFbGgqvZI1lY6kmvYMT7iRAlgV+RgJYyrPJeNT4fdjBWq6hI/8af9DGIqzogEExlPEqMxNz7kq54JiYy7DVOskB3UbktWsTunzjTB8XpQIVsbw2Na6/5IJ4aQ/fHZ9ObZVnWU4T5a1uDVSs6G8FbLA/gHQfBC2pGbBPcjyqCPp48BshBS4xAAAgAElEQVSjii262/s2iASLjQweq2uvni/IHPeMAndwWlQ0qgHgIC1ZuIp61pOIjsG/hGjkSztXrQk1a+3bV+i55lpPzANOQ/xtTjmbB3ojILDOy1HR0eoOQ/bMOD8/i2dA9zKgAme5NboO0MMiu63U0zHKPsmpaYDDY48/tln5nqj/7gDPXXfy2efBWoUH0G8AfUIN8LBr7P45X9d17tHfmczE2tjY1B8igAQ5ist5AJZlXwmLSqddI15Cto3UOmbnWak2DsuqCNSAMXdqHuP97iw3z4QakjP7QtkeNgzvwUKwJGQ3bblGZy8yyp7rJaVKlLrd24MXDaGzLIzKIKmcj/XbUMN0AQFofm1gDxy8CuhEACIAlbacZB7ZtW9CrZTRs7HP1fpE30HvCZV80hoApEBfBNH0WhTk4gi0EI96JoI1FOdaS7Y5basqRtgc8PHUbA7RtT7T/bYmXv5oCqSDT/2dJlMvVSLJAjXRdHxYDytjxR5KzguUGSo3Z3IJ2ToGWiIDLLLNap8ogjsAxXJdfNydzHJRI9HEMk4qwaXG5AJpNG/QHjON+j4lUfIu9Sbzj9h8QpZ2E5dvTqAHxGRmma/2fEpPDGYWUGF7YAGJNROiBTollrEIWh/zJ54+euSyzWjT5mBl4sYgoBwF1rtkhfBvO1NnP83+VCVjbqpNKj/gqZ4pM/nBx4uHlSG9YTMqPvFLP1vS5XIFTQC89d3v397+rR9aOv5tv6yE03/1V/7i9oPf/a1R72skSqRQ1ZSees3p+cX2937+17b/+r//he3sfJ1qenlxtv3zX/s/t7OHL0039blv/a7tmfd88FZlUQ5lrG+M61KBgsC4AahgRkUoXMFgi9l4MAvfEacuuESRG2gKlY1WzbHSSPJw8KdyaNEPnpLpddsYzVBSmG0aqkFoioKEoEoHXW+XXqbISxSx0TDQ8qzVWeLBSBt0HCoKgwdLofDy60RAVKBi4ihLM7k6mgiwVMGiKCqv257pDUKx80BoUzPxytHQGoEKCe9plY9VJhujNSjuqdCo5JPxvjVksp/jk5NQdqsgxfigZBqabYqYxibl2K8Y5D6cdFCqYQioPA2ACgr05j420+o+mz+/PYzsHV4j22sg0g1YDotqaM6PKPt03wMfz+ADaPrhYCp0jg8qBba004MT3J2BZHfc4UsxhZivbgCNItQZ0RXRDPqfrUNH/1qDtRd8Osa6D8rCMoPVaML2D6nWM1fSqwcqNPJV5Eq/8FKm654qEheKJUtEOesuvClFwTr8TBFTVMAKUV6QEpxJgyok2JhGnAxFXN9uUe7jzODqgQrUm0VpPdA7f+q8OxqYr3ctUaLf2zJQLdtz7A3g0dFuvojCsezFYkzDggiY0LQI1s7JmtF25TX6tXVE4lOB6/ijHTtjM2/kkfaCZgcCqMDRN0q1sUcF5MLKwVV1aEQXMkigZlz1I25ERR3DQlH30hWUUFGmso8qa1+y6CG+ZKt12vX8ltuAEXu8XI1x6TQyxuaOzn7PeKJElF2/huMex152NeeDTVdG0eFCKa6cGdR7j0EgBFP3ZwxFtSdAjLUoJT/hhrQfR70J46nrNOOL2ahnpaTEbyvDcnw2+H68Xp+tHd45JtHR3tr6WdAdB7u0WZzkFVBbjcftOEZo4kUWAV1r/M/mvlinycAEVEx3Qs6F8mWcuR1NKTBqSl4yo5g54c4dlgBSWaF4xY7XX86gOdWMOsDQQc4yCyMIaBZIkodPdYqKllCLPiNl/fO9jIroF9XzQVoznYRdZ7XdDg3ZlTZy/EKvwvmYpTO6sz10HjrHGAXv5Xq8TFBZMwcXWp0HEflYKZUz0nrO+EvBGNFTgoKr5Q+WVSp9JRTZCz1J/RHwbgRBQAHrZYI515S5AOevRYKfAaxguRlN8c6G0qj2c3wHdrk5Q8OZzMwnPceDyO7d215++eXt3r17xekMZ6+D6KShChAfH1sZGys1lba+v8vLURX5RHswgbWyH6GizEs/QWzVfhMo5XXkjcopvcNEhv9B0fwNrx5dbyZDRDV+K3tTIuMEAbgCwQFMXaJmvJeGwss8e8GbClNn40s8aj5sqSLTu3O2yp3Inmm7UQP0mJXY8bJmmAFAJmTueAbQXUXkK9scA3OfDOkDTvlSZtDdRM2KlEBCCwC1puCgAYA1k7PRZKX5MJgFqswTL7vDDAYbg/psuJN+pz9BPffEd+Zs954i7NMBUAzrb2Ozz708EcsswYcAx7o9Q1lByqTA9xgzwJss7TaT2d7zhDxpwXG2DLVZd71H469ZUQp4rMGdyK4C8KGm1jVgseF/KUW+3+oBxVO22hb0v8XcWCJM80W/QZQYQ8YMaCXABfKiekRdki5R3QT8IeCjXycBuRVIqUDFTG9Y6dHe40bvJv3hLE4ZMYChC9X37PRsu//gQdCwySx/9hIYoK3RByAs/RY6N6KqIP2vM0piybDJV/uln+bPqvWi3phAxfX19smP/hx7P7QUYAT31Nvevb3zAx/eb4hytG3PPPXE9lf//R/bfuIHvwPpl7f4ubi82n7mf/7Y9t/+j7+8nZ7Na9pREm+vvPiH22c+/tHNAIvZz/Mf/PD29HNvZlRERsWzD6HwlRRF6EfhyWmX0bmoV1phAKKmHg4iNePyFLY4/9r70uiBs9vTCj1FrtTLU81dF1ZoAoVDC5ES1sRLiDCMIVNecGj5OAhU2CSg5DIKiA1J3ZGm5o1RHsCvjnnbNdPIEDvY47LeFC8HOX/NaKbkowqe1Mc1Dk+vyUplAxoH9sBKjPRAhe9j5a8cB8XulC+mxhobCNkNAkt08EU9xagdisfKeGgj7NHQy4ZtQJIOH0TFzOpOYcxAqDN11vdJRkSjJ+X1M8fq6lxRBAXmZIc2DkU0gMuMIBkiOqTnomvueGiuLQMB7deDMPsutOdmqwSDMoOgkigKjSXh3kLI+oMnJ7xvwWxusgiKheCvw7UtN6QCbAZnHf/K2dGPvF6HSBRkUtyxjB/Vx2UNy1v3qBCgW7IdegdDM87VOhXPn9eyjiwVgW7wvNUyZo2SVOljuua5rqM86h227T7MgAqVr/ByeiEzFPnC+yd8NgMkIF/LrjEjDJFnci5MaoI3cx7pFevegROisZ4sO/7yO+P+bj68No+mQvu9wCjGQf9KnErpUHAj1uVy/mD2KuEzqQPcMLye2Cxm8zw5nmbcPTUCIE3jcp0tsa4HARULfYBP9ZNI8lpAhYzABS33cqo6QYe5+evRsDxpbXTi3FLifd2XrwysQ+WaBiDj3p6ntP/aFLQdqGi5z3Cp/DXK8qpv4Xmpj82dtf0zGqKert3KNxmBBv5InmklGrl/WEZpKxuWI6azWXqPztGk6SqHiu7DgSVQMQ+QaL2lLbfD3TuuiaZU1xC63kJvHIRlmX23gOKrFT1JvlU6XNEkOQf6rl7J9+3stBaeftOiay24xwMH3MGmp6LMiDtF/H0zKXo4K+6ta8RQLR7n+p1AzgJcDPSngAK3H9CwGLXesyFtsyfu71jXu75pdqAhrE38Xs5l2Tt7ciUceyynA1lyjNrmRe9SxOt8TDNK0JjyDpCNdNgdAGXykhV97tFgjJmk40dN3DDqp8rs9nI11oRWzFmZlOcTntU21ZaDU5n8ps8BfENmuZeL4tzg5ISzPEqCaT9LZLT3CHRdlXRk0cHMMoeNkbwlSrLrVWI3atuXkrtwGlP5ugO71370v/UBsGtcX94YzKNIfTpvzUF5xxy7zDDxBsjcW/O9nHjPPtjckN4Zua7MkqovwxmLMjOgvNRpZPZArqFnoSjJFchpsBH0J8kvd9Cy/whkgfkdVGYpzwm7xsAWA6hkO3ozdeN/yYDQW/B8OIiPInsF5YaOtkvvSXF3c0DGnNV3jrbT03MARh7gyEa/bJxugR4m76qsgZ9BCkxrI/maBxia9oI7sWc85HsKQNhLCtFP4v0WCGzU7Dz4SljuyJ0eqjZRfD1R0iGWOkBOn4s1YL+056+DQ2yOtj7Gc+Z/UU8DZaPY/ypN5uWJFjJTWaXKiAKJo+QPqm9kI3mtqZzwQRvB3wya9V4e2fsj5GXZF5RMmgRCcxN8HWnbeGkwBypauV/5uL6jbqPmJwBFPTeMV3wMngmk8mOZCRNlhcBAKYLJmXoHqpoYmMb98n6OWd5JWVwCHAyoaHoHUbSrj6wBaR72Rh+MejXNzhCBHwI5dE0TRNjZ2rMzQRyP7ByATOK96l+Y++bKyILWBcwx8FWNqg8INBDvgtfH8ybmWDJ64FZYn2qrHhVFInbLu+5RUdfgjQlUbNfbZ37ro9tLfzQv/WQb+LZv/s7tmfe+fzs6mtdp1zn61BMPtv/8P/zJ7d/4/j/lNdEO+bGD0ppm/42/83946af1vl9vD7/6R9tnPv6x7eLsUWOY64CzHhXf/D0/ut17/KlDXv06vUYSlUYSNTpXoCaln37qmVeaNEfsVaZBTo2KcNTBgWROMDXNMkZWDTz9Tm9zqLU6ecH8YGY1q3Ok1wUBlCE010aWRAIVUCigEEFJ88PLGvbx0PHULs/sSIXWlUGNwubg8+ij7LTtKYwOBSpC4fLR8/4i09x4VXRafF2MaWaeQLjZgXjX52VzEQ2ngmzjZw+QVPXwm5yOWR2Ls+4FrAyNGrFcBXwaKDiUYaTZ+IDCZ4NyzL2ds/ZMxrTSNaXUISrI6p9OImhKOYdGiY/t0dgFNK2iGk0n7eqg8hkebWZ0VBqMyeEBXY7GQ/VujEcHybtGBpV1Lk5OyUEptq5w89AT3bbOpIrQJ6Czmy0xOUMPyq5w9spDtTEC+7OWzt/q/MxlySj+BuyjRI5eCrXhlIwFOQeKkNd6xP+kdVO6URf3TmRTuJExDUfIjIoaqR7bGigg66dSaPTvjjkugIrUFbs60QVg82U+oKGlGZU3/TTKSd33YA18CKdZWvjutChGcfIX5a5sqXhmS1S3Bio4EZdqxVHUp1I1AE41TYfG2mtFMfwRNNzUGByft1kYjbyuisXgzKD0bda4ng/4vZftuEvAnEUsIaqSCFZsb7jzGuWm39CkhoxOailk5cTC8wcmjoj1wzIqNJ712je1oh207t6554mqj11dx+hgyVHNfscWqGKpXay9sdzEeOX7XaBitVTh4SqMUYymmzMqyNdNtK14V7w97vd6MeYJ0bsO78XcVntx24yKHpDKIzijncXPuFbOsDlQ0QJ1E36mpEw2GSfYAxWa08xQfi2BimTUjjDZhNWd22XhDwEqGolwCFjRbsg6CpGyJsuXUfpYlDIDQEabItzzA+et2FS5n/WGToU5iIsTTGmzd7w8R5RNsoxbBLF42R2vid7bSXAc7a/9/pAw13Yva7ma6gzunyTbQmSsaHfpuIhGL1kIu/LvZtmBs45UtJAFM/DT7qhrXufRvrUaL6UPTaoxOdUOaLfneF8Bb4J+jIa9XT13DD3nkPuWOpDxtTvHzs9dLHiteXRaDrAPxzl0XoEU/izxVJH1UEmy55DsY0TB3w0RFRHEx3fcMatgP3PSReawlWshYGH3wzl46eO7f/8+bDT2LLC3qs+jdBR3hrpTG8Cd2WSyz+yze/fveZkne4b1PPB+Fh4cBB9PBSt8T6vOTh3XgD3PMmHATjrqpS8BqNAa4sEe097GQrIfSTaMhn3sdmSOBhHm9CnY9+bgVIktm49KBnlGKkGRLOGFMcExzjr+V1e+Jrbm0d+DQVJepsnr/iPIDSXByLtH19v5JfqhqK6+70GRJ25fNsg2SlDbXmo9kMEFW8IBE2Ymo0RQ9npQ2SD5BhShr2DC6GmiEkONnYWgPKf6YEDwgL3HSgKZvPNSTZ5tY9UTspRSOwfp9yzNXcqaqdySgB9bDxvnOUtR9aCByhVVeap1cPCVgarhQObgA+Cgf8jpvkTiq79FZDZYzwmWAGrKbkGAxvoDYASfmjfqooAZM1G60sUh/+BDkZywYFtbfCtpZOWJjLYy4wP+C5Xs6vsfOP3Rrgk1iLaI5hN+GvVQ8DEkL4PGVQutVPxgT2DZUE7j0R+i9PDsAg98n9zfKENSvqEM9KjrE2vRHWry1RnQ6Dx4bKAzABPZNPXcC5uWeye9DNdnCTAPSmVvVb+HtFNt4uF8jQof64Mz+D9V0Qjemp38Oi/E7yGbi09SuhKebT7PChLiRSplp3e8QYGKbXv0ta9sv/9P/+9FloKlAd3dvumd79ve9i1/2iPcVz9GE08/+dj2H/87P7z92z/+vTeCFQZS/A//269t/83f/cXt0en5aPjGi66305e/un3mt355Ozt9eeo/s43+pue/fXv7+757N/tjOfjXzRdkpFJ/EwrZGqjww9AVcQgXF9yubHHSjcY5c/AXR/fQt4HKbKmLCEVvHvVvLzXFEs19oBBFc6NykLaCDo44OaPqVrUHhjRqKDquvA/OuN6LwDSuaVxDV19z0Mwnxq7SsEtDNyl+GfSjMiGI7JAC2Rp4NaMiRJT/gvRcRLHlN8VZqUhjKjxTI1+OzAXdr5zfyJLA3iqSBn1INBjuO5dGfrv2NW1N99pYKurFl74i3tzKFZ4ecMFLqoJYS0j5GIOm6gGUz+nBFxmA9VCzZ5hi5T9ct4ptJA3qsGSEnpfDgsMdytd+GZOymdNdmY0VY+roIJwO9XNVgJkcxJ7q46Y5H7d2VsbLSppzXatwZjLS3g/nSZTCLBIlwYoKPNHQ4doDdGrngFJxSJVF4zsoKvYjkAzZNCVyUjwyXenyfBFw88p2fShtbnWCVP46DGia75tFB1l6tKXuOtjIOdeauuPAWhlYnYQk8iTFaI5WQIDeWymeCGEkOhLL8G8aZG44MRV7lM+9U3VGiywzwqidBGJaZlg5UhoApYngTmkavzF7QH/7ylUgq5xZka7cv7hEZ0ImpaYrsLfukRsB0xJnpa9FuUFKvfaunpMwlsY1nDkC2/CtkcZvIvAwOscjtrl17fwv2Zl1fivboYt6PXh8vHDP2KzPamQVAYe9e+P6Ur7qprG13+faj/7jEajAWNqm3OKJdPLfPIJwCtjTVnV6u9IVI8e07zkIZFoMbcJGOJ86ctYcI4rRdJQOKA+5VtTeaZDO3oRC9U6CdIfYbX52FiT4ooDMTHO4zRtaheCAO9emOW8egA41Lq9MWrI4bsioqCu2ZO1u3HHPZP1w5s11KzkH0uEI/dSDIBZlSZbyabGW/fX9Pk55u5wB+r7JhAj9Gb/sASSqJ270H7bELlkWT0tsMZz6s0ja+Vm0JqyFiGiyFMLRT34OJ1yYcHQ+deUI61kXAGIF8WIxK+CZ4Emvb4Au0qmMDH3Uk+fC47+yTgGKlGtaMFOCIksWmZ3npancqYo67OjxgJ8I4rC5LGSKO7JYO17ZP4hgz0C/hlbo5LT7DASRreljcF2ZLy+0UumszslL7hSbsaFxq7YQ2Ugo0Vx9DHkWKSMwX+16OmWygx7MeHDQggFzcLoiWrzp88Dv7flmX9l1BgR4T4eTY2b2s0nvVYItTudmzxVnuDItcilwpsY5r3II9FlcHxloIhLBQrpOy4bA+BufqWSY1jOrDiATRkGcrr+zmbOBSGbXAFhBeVXfey9FheA7d3bzM7u+KXuGEYVe4NUFGBCpJtcXBrawH4BAAn2nyP+gJ867luQRwCbakH0r37DTiOkRXuoM0e4qL5W9M0a53duG+ht2NErdSdZpvLLtbLwqYSZndTSkx2Qy24Y2Uy0T5ddahH/JLhj4X7IgAm3bcmVytgv0NJqVDaym4z5uAxLlzwngM09Ez4DiuYY1LaWy2ScEzcxRokpZFF6+6/pqs2wrWzOcD7CRUZFEID3OQfSbAk+qCoXZlPC5EMzhme50wcwN9ydSiIDH52fCCqjwq+2woK5m96vHqZ6k0mheCtr3nllfE7stylw54Aw5rvNMNGHj9PJeDKTvfTL9OVv1fIFwQZ81MGAydenTCgL2/RZoEv4HW7QMWI0qJAQo7BkOZh9nksAbFqiwjvRf/v3f2f7oDz7BXhXjqptgf+u7P7A9+573b3eMMRY/RmwGVvwn/96PbT/1575zO7FmThMCtp4U/+Bjn9j+y7/989tLr5wuMylsY09feoGZFK9MFTYTem959l3bOz/w/STAWxoPy9l8I34R1hKEBKM7VkDFX3juEZDPoncpamMGVPjhqobGAYYwPX9ivKr2ptJvgWBS8ePvrScVbr0o7eTpkzhEXdhF1L4GLAc8v9kxDMM91jWVXt9S6GQaqT0HKiBa5jRWUd7mEt8C7J0Mah0MONDaCGtThOAQG7VJR12pCTVOTq93m+iyC0pvWtmW49HhA+NgYSquvXyM3sHBOaT60+ldXC0zEe6fYWwWeZENne12Lx9UjHUpcnNQCkp+RvsywrwYrtoTTbWB0Cbz1OHlzl6tIQ/IHAMNSPJgRCJFvUXUCFWzNPHcysGlWIR2P9ul+7qAinA4LyU3VVvtXIPylZvCggYooD+ZRdBEMFIp8vUkcFHf3isJ+V1VegpQ4aVmx/ILDVBhEVyl5wlSW6Gzm1Km2r8ZETpbj8ITYLQOG2l5v3Lp8LTKX4XWXiugwuYHIC/7/qzXVaNrZUprcBVTrTHEAHaDcXk/b4w7Ol4KSiqfu9JKw7yWo6pnRH3Mil/88wJU1Ojrdhg8FeqW9TwfSi+mJ0PLL1MKc9wjV0mew7wrI4w6Ighqahx+ZUBDxOgaRphRqwo2VP7J9fyXB1SANIqhtRA1a1/tzVlGjfyogKVosa28NWHHdCpQ4JGmF4MlMKEz00XBTmmETCtNf3FEnq1E7/B5OT2D1WTQzDIqRONtLW8ZSlimVZtoUS8z+ryHExwjU8l4S6BiOeWF2jEuheLu1hmVMpi9hIpHEsNQH/vhpVNMs27fB0me4qEKDfJ9MrNrVbcGKlbrp6zQUi4LgOXtbBns+cGEBnG+Jv3xe3ekzm5QWRfnlJUEbFhu7902pv4pzgHF0K8v8dryLLtjnyt4RU5SZWert4Ycq1MaXyzgTTsxABbTda1n6KhHILsmb4ysnsWYvFyLZ57KmYlM6PmPomm7HWdEu73XsryN7mSP+XrNauiv3uD1/m+gvxWwwNsg6aogl66NC5BxOMuu1cLVTArc4/0Ra8FSMnlkz3hAQik9W7iiXXqtYZa8lMyvEds+zqpGWnNrjxyGw0nZPFop161oT63oTOVqzYloTbVdRh/dcf0PoEc5NzgAlbERmKWSURcX55vV4Fe5INjjsL2wyNJzuH6M/g8/whWy7mHuwaHuOrV9TtvL1yNsBOwqgCCrqgB+RWkr0y3R9FtrGH97lLHtHZzTAHzQO1GOSeiCcNS6DDCn5vHdaGIsueAyxeSjVWZgg3JFq8MG5/qlQgtHsTutW57yjB4Ga1VnbWTlkNoEVFgGho3R7A85273nAoOnbL09O2qzUlwn6AdiTb/DdgIoIYDL1skyawyAsh8rWXV2gXWp0kMBDD4u8jECm66284vz7fiEAJCVULNeE9bI2gJJ2W/y7PS0aRjtmRBs9O7OU7O9bQyMSPelK7a7Sj9VmxoOX1vPzFATLaiUFh5DvictCqgQ4KGMGqdb9itRltBjjz/ugIPoUvfa2p+ePYqm7QALwNO2LrZHNmdbL1tT1wia4IZRtgVwxOwOPwfYh8amoJJGcrLXktRWusx7gXZz9Zk7oAa6U4URuwyBqknvKrUlP4/2GWXFtMaWMZI9QwSoRflRAsLuyGfwm9GBABvNWkCF9kdZAOiN0mUR8ab+XIwVLHaX7k2wElehFDzAp2rX6pkgjQx884wlX8u0zwTQGt1aFZboNUR9ogKpseEc5AyoCBmlcnkLXVlrK8DMxuwl1gnI4tl9f0ZlM6kXzBgU8oYFKsAIl9sLn/vU9qXf/adUBkdtw4TL0+/85u3t3/ZnMgp+5FsnrPv3Tra/8u/+6PaX/vyfcTQvFC4eVj/3f/2z7a//d//79sqjea8JnJVX2+X5+fb7v/EL2+mjl6ZOVdvsx97y7Pbu7/ohR9sXWvRklK/Xj5IBDwEqfvq5R1A6vcQSmwn3nrXiuIEvigpFoKWsqjZx6sqMtHeYwFTtvBRGLtLK2WlRE0yFZY29EEjNdVLopaR2KaQCaVwmtb0klE1REbJ0xmEogzG6B1Tg9MV9Er57BmToOxo7TzpG6ijaD0KZNfEGoMKPohK9W5RQt2X6skXtOsupKDS7d3KHEnBrNkAtRB0GriRQmePKdvjMzGrBaHBgFKCCG+NGJDMqbC8REYG6oXpHu4cZpVydrss6i9WZ1tF0c6iGwzvrt8Zy0YGpg9UiXRQBhGigbkyN93NcdLAknWgB1rXXff1ARXVWzcwh0TgO0HmIRFHmqdjHEtKfX4FRrcMMqNgnPY6FBoJGuwIqcF7IvZHN2StQoeilm0m+Wpjkq4aM27XrxWnz/H/BQIXRjEWToRYqMkm0Cmt/gb7RGmPEi6HCd1JBajmLCBZovikbK5e2yiuUTdR+lZLZRK41snmi+BZ+lVHk1Fp6cISsrsdO5fPJOYasxDwbfM54sHNjKy9lxOssrgZVeWnnXGr2oxo/A1CxS1ED+cKY6h2IdRwjr98OCiF93Mw47RW39Jhed2fgTa+LiM8CUuie1asbEK8uy563VpFtAdStR+aOEBq+1anT31ENoNGQW8tmp9PGmZ7nvjItIQCombnRvE9PcuA4TzJ4YHvNgIrZXPa19AbsKrzaRi3nc2HIZs1w+x3Gdl+qdh9wht7YysbctySQSlsAK26i1PL9wovruk33aulHazmez23p6RbjOQCoGJ7m8+1GZc7u5gzu78rrD2G72QzsvhVQIUeZMn4jGEhlfNwpit4a9gNwa/6zcqyst7k/+XSethTbnorJt3UUcmb1WZazJ9l9VkLSy4Yog6iULZrPbgJYujOZ9ckJ9kSEudc+P5yeUAZoDn71Nlg8VbXmZV8JbAtGy2wdnFJ0evIAACAASURBVHMK64GmU4/z1Cm0B/jfnLzLkF8OJHYxArBmPJ96gu8glJC0C5uDB0/0skIs1aRoepNPYb+XYAj0YphTJmwtK9V0D9HY12j4rCApD4UrAIO9XTZ/AHORhQBHscrU2ET60pzO5XyeehAGndjoTc4aQMF+NZJBiuxW1YbqcA7HO5+NEjKpvyHQKSsyeMT4CYAZ+zFHnzmjvWQyHebKJEYWAEtXeYAZMkkwt5LpT3p357iBG3bfcVsBIuwNBiVgDnqG3UeHqALAuGVxBosq+L1DzqV3DmhH+jezvVkqWWCA99tkpDoyIjKzBBHi1pMCvSGRGXHZnUWuuaKfiGVn8OxB3xSC+d5wGKXFjKYAIAFIcCCFGTyR9cEyWAYSGNhlY1VWhvsaGh8J5UBkA1zTP0T9udB5gFYTnV0+DIERimzX2Gxe1kjZaELZE3aPAQBml6OPCUAcPMvKhiPYOsqhWRkk9t1w0Ih7445v9k3lA5pzQ2MToOAOdQOfrCE4+8n0QIXKwNlq2ThODQwicKMxxjKUyim2XKYnCAwLc5fXBNBKmrWxZZnRtvcvaBF052cm+cPGbRH8IYO6BvE2ZpW4rT09JZdnJ8USqMBkYV/WXrJe4pl0y96i4tUaCBRnIolOAFAGa+AgAr1DrvbN2TXeJqhn4R9KcAT0q55GQwlcPhQAKxhCwUrKfjMfKNYeOomDlHyv+pqA51CNI0qD2eM+9Jf+xiE64eGn9uvsSlvYr3zmk9uXP/3by8wKgBXfsr39fd+zWwbKpm7ZFD/1575j+/M/8IHt297zNifGT3/+he3nP/o729//pY9vD097BLhdsEcvvbB99rd/ZTt7+LXFSh5tb3n2+e2dH/i+7e7xvdfZar/a4co5QscmDdFVRsVH3vYQ9Q4JItgeW8RBG7ndGn2hQEXka0Vm23ELqHCG8+wZ1Hr19Fg2oBqAimtESCCSQq1lgOzHT6N90vlGBDLRUh6MjSINARya48wpxZc0X02V8bIuHYiy64OZCHd5wbIkAZ7tQskPjWyoDeFmtT+Lg6Faw8o8kXAvLS6q4LWnNiW+KDT9P05+zz8zp1ApVwIrMiVRUnnYjolRK8NShy+MUCc4pBEXpc4FtqUeF+fJ3Dihss0oAleqp4BSWlKriO1QGHboR+vjCoEUZKXkMnscygLSmMP5mZuE0TEKbZb5UvfgtQMqUkHOOTTxZuQf8lJDCHV3W6ZxXYflfRoaq7UsD1jPIgQSIAx6nWdUNPMIo501aRmFEqWfqECu977KIWka7U70vDHjI/+seL+1171na06j3RtmQCplgkdZXYDgBFTsny6tR6x3ICTw1O0vHxrOosqP5YW9qy/XOR0iiqZKnmjPoOGU0ddLoEK0Op9bs9fdM7RPrUzHc2SYN04OdKWMn/4siL8nh0TjriuOmDpfGHyHq6I4JfrrEVntU71V6ac15RwyokoxSwNlIQOur6aH8K5XO3Z7cevApz1x7jMKa5PzJkVQ7hz+AVQwpX0GVgQtcsxjxkXK5+C1UpsbQ667oaAFGURdmTY35HZ2T9mHcjLiUJ6vzGruC2/9UtzvDid5r+GLzpNf5ZSXQKFDap9Ox0jtwsnR16wc0VhtCImB578RgIr+HNvVTW+g9+XXzUYWvTQO3tIkeqJzVfl0IKtOhzIFKpy+x8AXlDqBIwBmEssjlhKE85fcdpHmQqXaUfnEtmzq8KaVk3pxHugoqkDDrmPI86W4YGXv7Fd3nLiTDo2lQfe3OYnwQAfYJku4kgXam0ZBjkAfexAoRs/E01tQMZzkkf3RjmDom8F1VmS/O9A5ZtX+x5/VBsw//faYJ+VVT/ccgt6tYArvF3FuZXdSxsb4w56f0SDq6Juzzffp7h2WkxJN5TrFDhSnpb1DJXPsd0Upe+ZZ9F/gOjd9fNEgHCAangE7HyWI0N9BTjmUVpHjDz3jMBc5dR0gUfnP0qRatmplAXeae7ksOFrN8Xx+dhZZCXJai34VKZ46HfwQymTxMVuvdC9hA53RcwjN/D7KfmPBGgwKRNyWJoL7ZV8GvSigR47jYmP79R1QYfvnZXS2zed0cu8e/CbesNqyb0587eTMdACoZP6ghA1LZDFwsz2GqRPTo52miCuFnp1ufG5OfDlzle0hB7Y50m1N7RrfV9t/ytPw8ZA75fcB2/Cctf9Z7qxpHl16QGBdFQyYWRY9wGWPtSygs7PTYI67xydR0tzW2CPWt82d/wIj7G/XD7zPiwU0gCajV4zJuivreXKx3X9wPwIO5dw2oKL+VPmq3wWMI4sIgV3iGa1t9tNAaUrLWHAaDL9WUJ0YBgGPkSvFfWOFFNFfBRV0vfMbS1u5NcGeFQ7Ylp+a2WTjtXJRAnNUiEVbCRkMcFMAscbg6wmhOAiufaAiJbsABvlBNA5VbfG/J9l9Pj+e7f4/S1OhogX8kd4vyDKAPOPqCllo5Vmym32sJZik6lY4I9Cfw2Wp0Q37fMyktcpONzq8jwl+UslE0Bky2kBHrC7DbEmATcVyfKMDFXAebNsLn//d7Uuf+o0FWAEmf+q592zveP/3MTVprXqaULCDsDpDjEBAhLPtxWeX52fbp3/zF7fTV16ch2dsR9uDJ9+yvedDP7pZE+0/+ZkUvRA7EKh49mGkTKFOO70XjZ1b9s+9GzyEo86vUuY7BTciYNIIMH5S8yYcVn5q5UYfGYp8h4fN0XZ894Qp24bmq9ZmhKpQYFO1HjTdkYDgKLDr29r2MYDOW5zG7owW2wIt1Vm1R7uNcCvpjSYM1QjLgRqBOjjZm3VyRXNR+kkqNd0ZcWg4csuBZY3+LryJW7HnoIeeseJpCFJcI2NGjrIEBuLuWWA+tSmtYRzyJqz13iLI1aMiFP1KTn5wgA4EAjn6TqUa4+yc8DghOIfOGVuivTXPqZQqAk31NnNNWO/XS5qhNiyU8DZqOx1WTDnHTuJ1GpYiKhbfNdfymkZx4eChbJC3sVoRxZBGnN7OBm9T+TyjizLmWiqlhOLJoNCcZcj0ikC71i1PgLfnQEUe/Fw+yh6lpEpJldI4GOvNi8vEfWo3ReLOj6jefeFjhK7ZZi/sZWdpXAugwks/Wc8hlc5jGbR9/m5HNmX18mHyMst7kI4jw6m7djrvoEMYuaBRnCdVERa/xmlXSjZj/cLqjahxATQt47QBlM16TCYMZ3HVSVI+RJPDUUyXjS/RjNWJMYtwHfiq5amVwj+VQ1WF7bJU8swbeXaVUZFL095ziMNqRierMc9lah8Bj6t2DZ1mmEVoLl5Mmz2+rZm+s1sUpYatT+NiNS/Rshs17A3mcyiNDiUH1u8uDhEOOMm+K/1E+eQGVDG8/N3iM2ezHWWb5SUUkevrvQIqFhNfPX6lJ60thjXFrFRWlBNh01gulBvgvVFLXbSYfOVl+rR826nFeTGuAZvfLqPizmobeC74g/leZVTMIsGr8duv2HLNFzrdir96OZ7jkOyuy7fTo6IDXluWPYwSgrPrnhZnqjsBu/nJ+MeZwoa1pXntkiN2WGVGnakPa5SUE3N3/cKe7amrBDnsCNFwsJegHHMar85/6E8NJ5HkaDcpgpz8owbjt5HjK6BCzxjPGGS7CKhwVmj2oNIWOA/nV70Iv/fN0+u442r/JalbjiJ3iLk9gSj1MEVCJ8e+VoqFrUFdgS9LfuL1fijAwa8ocHOceiAaXxT0vQMM2TVWZkcZDB7JTnseTjfoIOGstsezd4TOApVOivOpnBOaS4WZYi4sryMHvaK6UY6I0eMMTkRGNZuPu7pez03Wxy8ZTTgbcc4r21bVBgRUeOAeHa/mNLcVV1ldB6hZSgpbADtUc0ZZp6A+dyAraMmD4K4tu8AyL/IaPSftBIVkJkV5FHro83yB/m7KF3uFru2ogH8CBW0OBjY4UHECX4jbKp4hCH3IAYk6v5Itabq/l3CySHinqUrx9kcF5lFRw9UBLxWHcq5eRozyUZkB9jfAoXZtj+9Y2ShmcTAz4+zs3LMWIjuHO47zET0h1PulglzwAbLfHBdSJcEls51TyV/2v3pIqGQZ5Fz2KAkwh2CPO5RZkgzA3rnvhfupPHJ/24695NbmmTr3uAdaRQA3tb9J1Q/IbyVrz+6TrenyiOCSwCYAUHejmX3st/tEW2ll4kH7IS6y67H+GQisDJh+rXQGYJ7yN4GW/Fqv5qHfN9CRlc9kxYwAH0OuiUfnZ/aql5H2uT9DSh4av0r9XWOTDqcKG6HTdUPw9TW+YV8K+YDu3jHgKhul29wt+6bvUSH1y2ltD6gI25Xl+6zU3SqIoMglZa34/nlJLZW1wkSiNGFjG+N4EHAR0ulNoAIHuC3qi1/49PaHv/ubFFa95oZD4C3PvWt7+/u+dzu+d/+1AwqsJ8XDl7bPfeIfbqcvfWVupB5t2xNPv317/oMf3o5P7t+Y0tkzyOv7b+5FSQmDA3TeTNt6VEjguE7kQt0YuupqYlNXhXx5hPTiGyloC6OCt8ORCNTRU8guSrqZn45YeatR6VCCC0mkaHozLOfKTmbxoMXhqgiUhSWRfsBxzNXBhVMwyABn3Wxua6DC19znrcnbWZBGq6m8ERfLA9nWxxQKE1Q4v/XO+u7ye5dkEQNWmVTOA4e/GeamcFFpljLDAykni99eLVChQ7iWe0pjRusFTcD/cvuxbH5hPgwVDbYgwFnzlBE7OuAAVMD4wpKJHklPIhnWS/VDiop73ermYKS2VldeiavRXErdyjtPau9cR7rkOVF2pOA6D3kmyMV27/79aGTmB6FHXFRQohhiHFB1islw+LoyKhg5pPWDzxdKXnVU4B08PKdslo2u20wAeyBuwL4hTRUyIQ0mdypzUypV6FUYi+SRr2LDp7NYPacLjrt34BidWlSFPVZGooy0lYOmMYBFb81adLLC17FegO8RUZn8Vmm3Mai/LqDCokNMdiJd2yV49GeZybRxnIPoW4EU2FzuJxyDrRAtzF00AvGLIlhS7kERh0E5f5ToodJtjdbC9nD3Sc+teKesaERsty6kV7wrB5KGMwy6ED2t0IgDS3RPJsCTwuPRZWFU4BESme9GxA7O4dn50K6x/spa+ZMAkD7a/cicK7PntPVS6xU+NwJLK5BPexFjWtQ2nztScQ7UddB7ErjRelBG+J/92aJ1nJ85MbZh/Sm7yqrjCSkfs66y3jtZw66nhZfcZECCgASBCPOd1KdpBIOeKVPcQC28UmikASoUHAQixL+owZ2/Q0YZfeOZ8Olkw8n9MZZvJ/TkO7FW1Q5+NJSIFrBK1Qn6o/1kVKMCbRa8sqzV1A62l4s5l6QVz6i4xUyWXVgmAQnRo2Kmm1ZPavf+1bnW11kPXoBhkDRCfQ0OR3GBznfwV9wSHKgzr9WDEfEfmnBIuhjyAjxJLmgn14BPBagYRFxppq7zXo40Gf/hsOl4/lYb6jSewROpG3KdBtqgDLuBaKruIJuKHNroR9oHzdH5ZKeHzgqoQMAA9CiXFrRZXPbcgr69x5zKx/X3ySkfD0x5HkBusVvCo1qFNvWqLAGKc1Uc2cubABtCfqbsxrXqm4DyJwI4Gx5SaSZpB5GBVgI3iq7nTy3lcNW4GpkUF3TqXrLRMJz6sRI7QIXKQqmUjN1kos8yM6BPKkgPq+F7SaDC/jZbxDISFG0ejvwiPwEytTqQ3Yu+BigFJBAAvUzQ10DOU7PjU66ojBVlg/evsAOmOkjNiYqSpeeeFZeBLDYnB928FQKzUNiHCHXfL92J38r+dPgKWnD7NBr2quQVPnO70/wRCloOvBO6iMubrj8F7Es4RhHEUmyi6sgUQOMD5LnKxQkdgEF06p8nG8V1edK10QxKSlECUN4oe+CVV17ZHn/iCbdBd4EKAmbXm+2h+YAAzghsktPcezTcvYsSY15iCtUuzs/OM5uG/UBk3xloZmvla+3Eh7X1ADU2Qre/zfEPH4LRkvTtWqoXJXHwiNR5xFPyP1hmhTnWkSFhvg+7QbyMkkrKHlKQHMpCIXsEwIyn1sTa2h6cWNCX901hzx8CCJKJo0hL2qrj1lpKjlTb03nx8tJ7YRg/eqAZMzEK50VsSdq02v9sqq1sApRcZyk3Bm6oRwXAEulPKBVsS6vm6gbePLj/AJlw7D2Dtddo8swPuUi6lWuEVuH0pKhnSX+Bys3hcwWtMXPMS6FhTAI+R/9gPhH7jd4xIYMIbiqjxvq6mPwTUKlzM6yGHaACviz2feVBY6XvRl8aBuDvYEkna1xvsk32rsnAvpye6JW77DqW99cgsKE5veFLP1UiMqHz4hd/b/vip36TjrdRs7INeuq5925v//bv3SwF63YqzYSmva7c6fbZj39se/i1L09BCnvnvcef3t7zXT+0ndx78AYDKVxci46zxuUOUPGTz3yNkdNI70wOzt8ro+ESpma64IDzC2pQqfNYDXhPc0NNYBN2+n0qtQomIMEeqHFPYjjx/DHCA+aAAsVco1GzEZUMFpeoEtblwoi2r+uR7x2daHIgtLNLJ2QKd3cGM+IfkSj1nhYEqU5MzdkVqAZDgfIkoZ6jhAA1xQ018DZPa7N1ndUdDSGuqE+V62HKYnX2SunAW5n2JoqoQEvsHctQ8CX+sTUGJ+30a+B1HI9Qx9XHX6NUZH6UXgioQwijwp3Qnn7XKtd5mOVapW2E3wz4ODm557LNlOfj45NILxbAghnzTtY85TKkclppttnfskvqs1CCWwQSVGWMLUwGYu7HHmwR3qUy/+KfwzyMa+FkUGRFpR8wV6HLMgeL6Llg9AZqKOJipR/3/C0acQU7cYvgXdGVHNygjTSLtNYDADIIkvEsgiLZRcFRcAXQQ1lmj1Na5vBo57d5ZLcMG/Bk0rmDxNVhOgxvJIzWDZ3uq6wYU3mdDqNJ2PIMLPLm4hX07SY5Al/1Xbi4Gvyr5pzDeshg080N4NHWkh5kYScbZ/tSP1Mafc8bVQdpJGyAnORqn7IIpDbfbOW3eKX2WFn5mFYOwnSuFebs+a6csqPSL87imDmAWht1jGbq95TnKLPNEEk1Mn7ue0uzMEiKE6DZwPZaATZ37nZ0X8ftznHyEJ0z7tD3gAs6b0r1gBU94GjQe7S+Kh/QNaoTXZP5RL92V6SIFwcTHIQIpuh/mj2KbVWx3Zuolz5hLfaqCHzjdcsxrFilOkyqrjMaUjm+KZAwioO4YdkYvBNXdVea1Zgyz4ROaAHb5WqoeHXV1lm+aZVX824AxXr0QWGj4zP17JWntgWxoBeq5EMFY+s4vbqZHLb8Atg812DoVwPH3vBzg4O/yng5CqRz6FmtI6h1SkjutUBglV9N2EdIr6mTvwOZmrks5uEu18m0VzIW4hQ36Gzec5DEGnRQp+sRdJTV2fLJN5HcfvZXLnxzyFKt4thnvImgH4whZdxwhFRazh1pgY3pDOhwb/TdcuECbVydg7cBeuwZyBzKp82CUXK/6FzeyRqZTdEdnLKTwXCMd5hXdjAaMqem/W+2gYKPzOnqNdpL5HQ4Swtghfn050b7t/otmHPUa+jL69fY6bnrQeMNa9RnTs6pbu9SB8/SXhXgvnty7BHH6mkpIGBF+H5GWsQ8+wKhrAmy7nO9K4iMprs+F225RG2UPYJzXP0GLLAvnLkciOr/y/ntjv6TY9cdbC3NDnZHOR3tcHADXPCo+trvwhoaX6GvEfYbGSKZfd3r+yoRxb0J0rUKEdas+cyd/OY0tTH42I8sEt7qzadtAVBMJaFGCBsBnMyquLz0Z1rUv41RPhM4l7PCgYNZpDzfBwYMyqGtfQwHLfuWIohI2ZqLAIPYt9a3Uv041VkP2qHkJNgRAXilP0rNsujHBzrBM8Rndn0AKAUo9n1nzwxlodh9tg/37z/YHj16iOoGXvf/7nZ2fr7dv6dSR6x4ECCjBRrae0DHFpmvaH0AhJNePxw8xgk55eDHyYnzlJX2Qk8U/KgvBIKMsx9plYVyqLt/x3wV9OsAaGkDNGZnY71O571AMQFJ0lUE0nppJM/SZ5moIuhBRwhCjCwB+gv78wiqOXR87RfmjdJmDjCxt236nLLp+0zmNFUuyrg0dvvfspNcFpQAYfkGfA14n/M4gdEYn0pIlvJaPi/VwSJzaS09M8rWi5k4VoI5wVYC1gIzfEFcw2iCGKtcFxAHfyFoSBlBvkamor6ZUdGShkW+v/Tlz2+f/+Q/cjR+pjma4Hn8re/Ynv/A92/HVmPvVvEX9X3X2/npo+1zv/Or2ysv/uH0XfboB08+s737O35gO3nw+NfxrtWx+3r4PA0oRN2opMw8o+Inn/kqlTI6Oxi9Gs1R2VgqFEE1PlIPCdcqigLktrhqYqZogtOY9RJZt3JlVJhzWY2aTHGwiHQJzRhHOIhd2pVIgVEZq2PPHTwMqOiNN8rWDhCwZ41N26o+KaFcD1Y3mCSaagha+MiK86FfZwMFSpmbfFf28gjHLr/0uqV2QPKwVVaMIgp66tbbzWnvkQ4sGyOhLGFc5zYLfU4jCohSdRAoMa7xJ1WnXJTIMDTcDq/u/lD4S8QXhbeNGwffYmZclwo2iGJNAbHD2A8+b0bGhkWdfVGdnTWawN+oQ6vyR2jhRZHROBzs4FhLdojsk9ZvOHFMxXxEnnlNHwUFY11pnawly9RjcNT83uY7UwirMiTnwayUFqd1Z6ezqErCRa1WLmLR8zGx9oNmc+VL6ndcNA/+7deOf5eGkzj0V7Jk/nk4NgvAF0pGb50HuIa0//aka01xKE+KGqa07aK4PML+JqAipkk6W3gS2gjNioTO432bRtplIpJtWnM47ticpblOZ09++FoBFaDX+tOWAOllpADhirGCDHFeCIyTIyPPFvUBKJlyMyLsP3Mlt60Le5MDYxmGrsOJ+3oIUDFzmLiBcbePBMcq7gEViKROJ0+dB9hJz+B1C7mcz0igQplPclrVZy0d7X1Ftsnatx8dIeuxN0LYPDEyOjVuX+cZT6xcdKXsxo1jKRkCt+lWC2y3MNLiRc0QZ/UXOzSye8zSWTiRmavVqNu/V3lqmIHrTdBz3KHiTUX7kjUHLPBqaRaO1/Sg4ca6Bi0gnA9WvWI5tYxWrda1avz3Q/Djn2cPgkhIBwugQobtgaIGl0XjAkZVR4BOSstGRysO1sNWdZkXsrx9RSMrWbc6mZdARQFDDgUqlu9YNDzPrLV2mklOclxytjeASZp7XRs5jVbz7D9fruthG8mr/viBCh3izfxKllEzHTaVbvU8nj0LlIQ7E2e89IA94AsZOMxUbbK504mkqgHVqQ0W7wwJMGYzDZMpp2en2/179+G6cickGyRLTlQxTVNcez68Y0f3HuimlKtpvmNVhOoUVibSlKTM6chGxeask+MOOi3LYsnRHKV+iu1RCBjljrLpsz3DHPNeAaJmfdBZq2Ajcwx6Rjud4dUp6jZxKZVkc3CQw2w+OumvCGLVnh+wQxH5DztPduleyfLUf7xChPeftChqs+VtLVAmC/Xw4VNAU+51MARs1HR4JyiWa4seHIgmz9I4nvcSvTRm+w+dC+csSsgiGM0AmzkblaAyOlHTwZyNmTNrAhk1DixcXPg7DGwxIOeuG3IYo+8JmwtXGkM2Ks4auyqrKjAoQIEtBVxG9gd6UtjauaP+8pqZRI+QJXJupX8suwLX6EeggP2NDAesix0HPX+vfCrSHGQrCvCyrBgDKkR7fjKH3ofG9CWFgvpHa8v24IjWFqDqRYAYzRqWzBa73kATNU335usEXG2uAvdCphHoisHwwQ7YFODP/kYJugKjk+dB/9moXetmY/GMDy9ZnL1UBfCsVLRlUCr1NYEiqjIgUAV6JOUOH+4Br8wkhE2EEia1lJP2MWR6ASqknxpXKJDTVCk/w83OKP5ZvJo6bLUvYkistFEzsjz4GKBXBB69CVTMNRvbjK9+8fe3L37q17fLC2t+PapGtplPPvv89o5v/7OvugzU+enD7Quf/CfbS1/5/Byk8J4UT2/v+o5/dbv32BNvUJDC2UWy8MCMCgMqsswLbi5CcgeoyJr/qcjKxQm0nlGWJB3ViDM54ErA4sebKhHJVLSuC8fOedhEs4duszIvuoQRCUqvE521GSv5Zip8dbnpOb0y1QIVmpqyTGp5Iykh9hmcd56jEnqq7BfMLw/dVpE1cKZPKc/rdXg0ThwXaDhctXeZdjyum5RJi0SwA9xODFfyujr30xXvQICQCgugItarnBXYFzZm8igJAyosgqSTMeppwYfYep6coC6/HxaK2gh6k2NUI28dNVLMpAQ5R7CJUXPId878qpTl/neO0XrwDPSvlAoqaXVhu2bpUs6aR1SgApjQQmhjPvWAw4oy8qbMyxW5WrqgAoT+HWSH+tv4gb9jgN8WqPBokgp8lIgHyapmTxj02k98BVRQ2vFRJYJ7Zx7ZVrF9Sw9U5LcqnVGu3wUq4ARr11GEQ6OI+5CccFugYkEcvQZY+bhBXtdyNmk/FdPsV9MCFQkU9GvZcVrzugPe7aIwrxt+a77LknFyUDhd0PCHLK1ARZBLShQaVvpgyntL//Uk+kqKrD+wm+9SS+egbwFUcGp4i4xLRev0yxxpi1PpA1NASQNcvArsNO/os9zKPHXaKuPLJRMb30Ge54roLJsJOhvuoY46nHUQmpLjtYGeyhtIvmmMEI3DQi0ELxpyzn8yXR97Uq77FwFUNIOohN6NbkFrK6BiJft7Cu9X7FCgQsNJeaLw4WsvATL9OZQIlruGL1KHueHC8rUDFWow6lGR0KHUvLV/Us29Az/eAFTctvmHkzhmAv4i+NgDV2Vgu724pkvxjQlUiK8qUDHwWpnPUn36OoGKeOeBQEVd4ll525mT8SYKvR1L/PECFU2QTUOXbaZFM2dNkJsoPWOVKZugPk6XBCrmkdHI4sooZsg9i9Dn9XTEexT6HStnY02kkfGVQAJGjFtHGWyfm33Wy9RwSBbZ7L+6P7v2HPC3MJGI3QAAIABJREFU57JMlJIVENM7WuPcszI9KtFEGYJMbIKe3YlbgRU5c90pbef5sQW/3dkenZ66fWnfnz56FHXxA6gLfQa2oJpxy0nv68RocpusnPUYF8ozyensZbGst0IBZ2Xn2hxtbObQt9JB9+5ZFZBte/jokdW28rI/Vn7K5u/PsObNJydNQJqrEHxvy7eQuN6DwEvrIMvESyKxTLRVSBAwYFdbf84o1VxKCPqOEsww57zpKXKon52fZTPeALeTGcJGDdnPiOwA/UEvxnMOQLmjGqCMg3IEN4bm87xLZWXFG9VZHnoVm1Z7lpBlqzK7xd5sZZA9o4VjFwhm36nvhOjf7U5VWGBDbL0PS4SG1LJh/cwlPehcNfo8fXTqPSHk0DcXcvg4wvbHenh2h2IQyWsXnolj1ULA+3JQr3Qh8BKvY8aMBUZ6NgdLPEEGqWSY+iJgHxvdq/bAUSbN9bYZHXgkP8GY6pvQ+LRG8TfBCK0/7PoMCMkyvCzZFa7GcpoQJNZ6KNrf/UySxarkQV5FSbArlLwjHRqfWD8Qu8VKMYHXLLvlajs9RUbS9IcysV0jAB2oHAs93/v4hKxuXUpaK5eB0QcE/XG8tB1Lldn7q43g5QkVwM2MGc+IsqAvOPms6D3LimnxXGLEv+g3kUZQ4Tn4Rf1ZKgnnumRmv/nnb2ZUzEgDNcJeefFLnu1wcX42ARJw8D/21LPb8x/8ge3k/oNbAQmXF2fbZ3/7V7dXXvjCInX2aDt58MT23u/6we3ksbfsOsrm1P0n6dOQHgcDFSlQpdTsABVRT5YR7C5wU5F1hJLR2k3EGQU8Dj82xVosu0UphIAl8+sAwHFflC+c2rfOqAiDl6g8Di6UIEr7QcqjBAkGXJ1Z1RHTHkxq1j2r663SWSX7xCONVfO3zvFmoKLdv1Izu1undESlgHVhfVT7YbSbooNDtRlNQbG0OaXWDsbc4ByU4sPnHghUYJ2VIgxgywGsohBwN/hgHuxXlkJ75UolBDpqTTbjLJEakPitG1NmvJwMdonN2xW2wSmF1yt1FmdhLRKOZ7c2qU6hXGscjnWU3X3urednK3FVvh8M0coypSSUBucjchrMh0caLg9GfaMMGVcAWZcRNWGRfeKRIAtL+DZAhb3Plb/eQb7jVHF/8WJ9Vsa571fJgnBu3wMqFg+6LVARfDsU0JYyGlZ2hzpJtnCZtW+3yqhYrVJG9EKy5q7HPnR0eJPTo/JEzahYgRQzfhn5Z//MjusX8qhnytoPqAErCiv3DbX7McE3f7ua9BAetwQqlLnUL0EYpvjikIwKfz03sDrwXJ71JHIroIL9pfzhcv7wLCBIMTpJJPNSfsBYK0CFBsy5IhJq8iPcYZ9MSAZ8gh+/Br6yrjDvFRgSToOmv9MBL6iXlFJ29eMZyI1zZa0qLzm4MuTiov4cW4Gvq9ndFqiYOcRW41dpwIQ5iwyKrKYsbwEjsO3N0azt6jBaHgjzWRdSPmjTnXbp1LP1VinKLOcxPsb1LW55OGvqOCf9ZJaDmYFMzhfScKDnoyx8OrP6590eqDB9vIRPipB1nHXtUPYWc7lFS7B2vamNPdJF/C5EyHRoq/JmN2dUBEfzuXMOiEjL9oCZ6J4519uCFTed2e3E/7iBCjJEOKEwuupw26OhDGhjiY7JxVZLPKQMbUrXb5d9lFQfELZaq/uhSa6tcZTgYekcDjz2P2hyAlRYFLmc4/Z89eIbM23iAI855P5W4GKkN79OLoMG+GCPSLu9AnN35GxHLwGU0ymOsvo8zxKAzSYQwJzNshWkZ8lxiz0tsqgDYrz0kvVOUCkjvtcCZNUsWs5Vu6b22tDChE4kx7xH9FuWCiLk05GPcZjdZ+Vt77BPgI3fsxOslLXZwecXcbooE6L2YOl9CRalDvsZzmrPymB5YwOQT6xvIX0k907uY93cYZo+DpyPZrQDoHHasIx/u4/loLCvjBpRX5PqxpDKIzuH2Ulpk+CcsDU3YMWyVmw9410q+9PxUrWdBDIYDSvbIfiWEfZyhAvYmGWRyRZrSiEVtUjnpbL77R3SZb0KwzEjGNho2jbM5mTPtUbfdm0FCWoMbQ3M1FgdsDhCn1V7hoFXVvpJTmr5AlCGus+WBl2hETlAGsgO9hswIEzsHL1NWqACLJYcXrOJoHPAZq6yq9qzM6DCn2l05pk3bQky+0576b49lSQre9+AyWr4zhLczkfMsrASasgMQ/+WyndeHongmIAKWwwvERblzJQptCPxq9zgOmHPUN5PfpzIRqj6CeWPr5H6zJRzWPSk9ZRElZ9Myls9DyoocsfoxA0a7qHbL9kDzH1VcmKQsOWfqNkmcFuVklkR0PImULGnCzjzvfTlz2xf+NRvbBenjyZgBRb2sW96+/bOb/ve7d5jT/beu/H57Enxhf/v17eXvvzZpilZKhVH270nnt6e/8CHt/uPv9FBikZLOAio+Klnv0YFWA7l1qkgZJeqYRPHi0ONjhkpOwQS0ukBhkTZp/3a77Gnqu/JZlwmHF3ZkYOmKy3TnL+dcr8kWp8mhC4UWVNKQKN+0DHiQPdDENPAoyIbhy69CU3zWPVc6KLTU2FCdEKCDBY5jnekEyEdO1rrnA9KP2m64/eM0ml0Uyitqv1tgk8O+Ll7N5uCwVkP5Rz1QMcD2LendxSLRnR4TICKmJMMBDmKieb7mhBJ9qgKKkktQKO9sygKoMyaWzrg63q3JYQq2cDAQKNrZR5YlE3UD21SzkETofBT+cTY2OgJmhPo6iD/MPhKPIf/53Q5o29FvfTfxXq5E2E0VYXUJx9WmVApj2OjRqeD1ZtyOU+1zY8rX+9FzqL0UwVJW2dpv99T/9PS+5WpztiwMv+SPizH6NIBSg6drXuNPmm/n2dUDPMpN4XiV+VRDDusDNId69jeAqhwhGnyU6miFR3YU+11Nf5X5TnC9aXIJ1d4lcqesnZYKxoa9fNcq4Gqp/NoeG0FVpQJNtlT9Xo2yXbJ7AZ7pvZXNpLR7Z8degbFyCfx5vVQ62ZYJE75pkyGC/+qgQqchpN1nfO1LoSRn80DzZLujSIp8JCZowwSRA/2VJ1wgKgqW4i9zWbSa9qop/Y4HUnUoBUffgJN/lwa+YqIsidGzyyeU0todDa9RbD5WreZ1+IvR8I4sSUTdzI8jpj1obQCJFb6wooZ5ztdxtNdAH88LbWGyqUTSRYx7V1p80tpcIOwO+C+3pdf6W4KxIhGVfZA5QwWEfk+41qiiJk0ja90RA+nttZa0SjOOJYrAdvKqYWFCH3GmWO2e90ZyvUDC1X9pVvYGallfM6ESRe0uVMDfBolUYHN8vsyIGEJhExVJ6zZYpn6SaX8XvFdlqXFvYtFC/mzJt4Dh5QPmDZr/gYAKnhWaD5VHu+xbpXx2KP5itQyunXNV9dD14M9pJr4+lvvMTLz6HkvS8Nsivp+DgXvGPcYEdx3/V5z9rojugDzMRO/nc+oZs0w1UmfgxhPXiywAPYs7Rg5wjwzxEoUwcFqJWuyTLRkhxqYZ/a+l8ixCG82u1aWg91hTmLPVLDSP94cVrXvySllnXD2MoCN62HrLqBC/CwHvvpYSFYHv8tpbc3GmSWiuvh2j9l+3kzYxvTg/mYjemSZFRyv6YIOOFg5pchbQQQ8wObc0/AplJryFxdYC7/es2bgG7F9hpujACiwikJbsh3xd5huyshtG5eN5cGD+/48gRbu32BgxaWdOyITyUCeRRW8zpQB2Pyy6RCBrrJmE64jCdu7UT0DcszmaZ9FBLs7ZgvwRn0O4B42u9oXcL4DNNGP5mRXV4d81S9tH62hdpQXukSzd/RkhB/j4cNH24MHFjiNclDenPj8zJegL/8E5zXW1n6UCeJlotmDQLxv16qfwEw+eblXrYFlGBlwxSoHrDbNTCsF0PqTcc4kssi/U2KJz6KXAcfR6yoByJWz0NbGSz+VBukOKqgPivFoySIIiSX+jHEBoFW2j8bs5c6ur4K/VdVDDnf7P4KCKCtQ2g0ZSO6PMVDp3omXz5z9SFXJMxZXKRumgjDqKSKASWskUMbuO3aQFb33QA9ZQs6+rxkVdTyyDV3esEcP/G5WzgpMGPaS0z9G7H614vqBvU2dl7yozB1fr2gWn+V038yomJJGfmgLb02u/+C3PrpdTTMrcO49ePKt23s/9MP7DbYp5D77yX+4vfSlP5grGIZq3j3Z3vvdP7I9eOLpm4GPG8b/J+PrkBoHARUfefalxiEAQYt0P4m/FHJuhjSHha7p9T+kyOGwMkVLqYmO2pZ0vamwsRHpAObrgOxbI2iOq/plqkLWe5zLdYX/fRp+2LHElJQzOCf6cj3qpMBD1B+Ep3kKpBt5VAjifWms1ejFqjD5U2K85pQ18KIRdziIIrq7fps9KnLKbf+GihrIee0osR08li7rzayQBjfzGbm6xetrvc9+z5bOjBhYZnmMPSpAU73TFuh+CyyYEFf6Z7t22C8DMBQpofqhaVAUsMBXuYwpUr2xryb8Xck5P0dvDjugzhG1I/7AGtRa66z36Y72zMpJ5axFKVRrsa4lyIiw2aJuU91rjSGfQbMscIiGMcJ3AeMCtSGx7llbPpm7jKx9TOF/0JF+FJEhh/2Ut3csZwAVzMjA8ubzG2dzywfNGk6dnwQl9YwKNPk70pwVULHndVhFH/flYcS7WKNu4g1gNxqpzlON7CLNdv5jOaO9ItrkZ8w+o8zZqYujkaYoo6LEL6A7FRm5MP71HGXYAQxGNA1+kl5jrQIMbve49f2v979fghRBuceFgOPXVUZFBZ/hdBffg2wi+qmcCaueHfMdmoEC++kAvRJe15Jiyf87HKgAo+E8lEFcK7HmXuVW9zTLMnt+VrGsnMoaqnxfOEZ3hIBeJfqEeALdsG8GlvpwoGK17qMuYd6C5NQGqLDMTk5e55IMjWH9G4HUnejzctNBVwJn4rxu+gd0MxnFBi5YyOt6dwvurDPgVmf7MrNwJQs41tWQe194AhXNqFmTGpFkJANk9HrQxuLph6zTikjK5xWoWL5r8pzqtPAACCtHscj7E1AB+crtLDQ5SXOaAxVanH48ETWcgKKfZ1GTPm9I2Tbn16XTdw+onX33mgMV4ya4rG506YzIX+7lipYX4mteDqXNVq63rqXgCFSE6lLGVNe/OugOIOXlJX7GDd/+cQMV7YkX8171qBjEZAqAm4GKKizW/QZsP0yPlsNT8gg6NQ4xfeZRwV6GZa6kwUYYhZRnLFhE+NGd7bHHH9teefnlcCTWzACJfNG4pk9rtTD0ShBWAEcOM0YeK6udDm3LLlDZOoH2Knmis0eguwcoHpvT/9IdlCgHw5JCrIdvczQAwGwrc25bA+OGHwni5L5JF8U4HVS4BMhh9wk0UraHAAzvPXB56T0tvFqDR7XD8e7lhAWkHB97+Sl3sB+feONdAyps+raH3ribkd+114V0AOiIhL1IBxDltFEZ7GJAhTVqBviE38/Pz6Ksi5qOu83rNQ3bvTPt7NJCFUvwoJX7wXPMoYtgO9kkDtx4KWU8KvwQAiqYURS+GQoB9OU493GZQ9/eZ2tYgzUqu/n+MmvE3uXOaqtawR4Z9j8yatBI3INFWQbLgRprLH1mtrbtK5pDa1+xthhYrdph1+lzgSJ2jfUhOLtgCSRvko0m7DZH75viYAUc8+bAvn8fGSznZyo1dBJZOUYf6tUJOgew4HLAelwwu8Lul6NbQMZ4BFuWADKR7J02FtsGLzflemaxfVUW3D8qxh/XAeZraZ7OMkrekJrrYmsqMEB8EllJBagw+91BQ9tvBgur+bvKtrku05/h5cAIp7/vd/Ky0b9lrdk41IhbgKSerRJG3vDafC8ECQCMoncL5kQf4uQUq3pkPcnsvfZ8639ic3SZxUoEBuAJNPGtjebzKC1mtGHLbQCJ8SOqwpDja88IbVvTezazW8Az6Ini2R3qq+PlAWHoWJ8aAJV4WLXJVBIf76/NtBG8C356M6PiIP3HwYoX/3D73Cf/0Xb+6JVltM+DJ7/JG2xbFsTskL48P/XsDOt/MfWiWj27x9/imRSPveWtB43tjXERWUhKHDzwQAWvLrbrS0Nvz7eri9Pt8vzR9hPf9GLWCDy647X9velSCJ+29wKQP0TaS1Gw/+1vHH5yPtWD9YaatZ1Dzpq0+080t0W0QY16bc/tsXyPlDcXzNr44pCEo5qCgIennNSDMXgEoEJ9JqSIAtFMt97oTJsrhjMjFTEYmSGRtCoHG/6XgurI9xVQZQkznp90BqL+pw7O/jqsT9JKwxtrfTYu2zO0/V0FhIGuKau7fbiv7KTMTs0KCGGdnk+MozHaMqOiyhO81pRSKGreeM0RbY0S/9e9E12012jqNJp6I7Y+YGGot++Y9XKgV86nhr4PlbemNr5OtDIfXbcywDMCpa3Nr3q4vt6FwZoDv37uCngtc8U1YsM1L7+lSBWm/6JxnRoPZ+SMDtlKh04DU1oskc6sDCVeNGfmbtpKQ+ghGApdTy9oPlwBFYoGqU4DAWWD+X8jUNEZr1wHlPqE3HGFyw0uA/BErY0wnQP8TjNljxu5OPdzwsnDd3RABegFsgmZTFBIZYj0q9xzn2QT/h/3pN+RnleTf0nPRBAELPj42J8nNzrXqT8foIhnNL8bmqVevOqIrp2VFbRMw7q/Po3v4piiCBBwHgBCWYSIvl+Sai9jbW/6DLj+TM576KroHFY9I2peSRPjcA44SA6cg0vxVVPfhbydO91aOd6CZQxS0JnKMzJ1m9kMcXJ7cAfHATnQgnHiTgCQoytQANh8ORbrWKPv6aWSATN9zvhavwyO9Ky5Ho4MOjVuloh5xaosjvvC8bJ0RE0SzTAg9lHIGlD+MYw51PYOXmr2fj7BKo9rwEadlxuRXE/NId/BK/eSW3ZocOUcmq0r2lcOEi96QNn4sVco+5HRvO09Wuvp3q3OVK79aI/RMC9718v2+p55Vf89Kmr1jebKBVhwSIG9vJXZIt0QJH+rjuyONJWyWfWiWI2Jkb9CsOXsqeVDjLgRIWr7lxHE/eqsHOq3AcjE23pWOCfJ74gUBb01QMdAywUUduFQ9DZn1jnfLcQNpto4t1R2hHRQHam0Y2fPcvk+2SPpWtJz3XlrDn/vc2flg7qALoc5eeoxSMmcU6lHsy44ndreb6I4R1PPGPk2zJ4oLZxz15zggKJTmY4ynDk3SV4oC64rwKvV9JODXWWOYesXWeqtlcfK+VvpCucBGkXr7BNPqERWtdlUys5pSWdGrZ5QF4HTdwc8Sy6B9pgV4eCPU2QIXR37oNXZoqh/WM3mZFmkKO2c13hAm/WbODtjtgHKA3uDXTp6fUysOOBBEfbmu3CyI/OCvSUYhGF+E3dyK8NkwP6lUyKgTvq09cFwx7Ca4kb1AEOnIes9C9lkvoLr+GxLipaTV/Sq6PcZ5Xh2jvpC1CbRO3Kot/OrHRO+laJvy8lsvSa8jI+VVzpHTwH4SuoesmxSlD/CHkUwUylHhf0Axwg8sd8BVMF5rMA7BwiurKzT6XbijejxnTeUJo2qxBBKPl1Hs3Wnc5Yp0hpKRoo27BqBEL4GbNAteatm0xkI2GdyoZSTdDX5zXzuptsw2BGligBkEecKOa0ASFsRA8/M7nIAhr8rkGclQZp17rJSZveonJTOCZUYMxABfgNkRmEvcp9DhrKM1d6ZgLVnRhL3CedxylvXsy1DgfLR9/X8AsG29FqgHB14x368ZB7BUmWOYs0NfILcsR8DVhwgZGN2o6ETNZB3mQFAcyWYa2BYriEygbJyi71W59yRNwu/ukKmyN1jmwNoYHGkzreTIlFZZG9mVNx0bupoub7aHn3the0zH/9/0LNisuq2Mfcee4tnQxyf3G82/+ryYvvip35ze/Hzv7soD7Btd0/ub+/+zn9te/ypZ1+FY+rAibwuL6MoOBCo+MizL7vz1ojcm/zdReqhgwRQYZMv6fR1gRxAhRl4tR4eDHToGlIqDmiux0thSCLlEmOQQ6RDURt9BUqAdJhUcVpndo2chlXK26L8Uza9aRQiAhWK2kulTgpst065Ao3CFU6RKV1ZRsUoxqVU23I4qkzFxZUod/JjmbO5pBwPbtKGsleNp1Q+xoihVjm+UVMeZ1JKE9cDeAVUQMWmsaSnFcUWpKgasLiAPhn8keQeQFmjXHEKnmpZbpaiyQ+b/1pluF+DA4yy1wCokIPSBqZDeWak9gZtvWZq1Er5KzsXBpPc16ldYImL/O7XNguVjbQC4yYNYXtWGIoEYeiXnSoA/t10LTEKH5f789OpHA0FbyW7c+yHUPxePffe4JNCdDugInkiphHrAAbzhn/WyE/rUBukBh8tMX7yjoSuJH3DUoNJKDrxOcVCkSJYy9jrcaoB5GBXjqvrkruRGXXw801s17hrhF1lB7x18+yPMpSgaRrIIM1CEywRiKi7UQmfCkEeLsquaPg0FlJ3JlDhhgDPVxiCAN7qyuH2Xg5J0I3GvH0ylLYYEMB8A102BwEV+2y2z023+RarvmfmjCO5Gago62rL7GWfkhewF9jzuYMQ9WXFrXd43uo0a7mq8NaslM4yOnhnlSAE81yDMFjrw4vlk2PKzxoFdlSmPFSWkt9ml6NnQTkLSqbIfDlQChNnPxtYhk5b+PMQoEK1nsUaXZZK6E8Cfuo6dcu/MiBXDuRw3hFoaZx5k4UajV1SEXVsBTA4WB1RsBPaFy1M3jFXTyQ/WtkHSSPDOfnAyWy8FLLrhmNnJi97h1hc85oAFTeXnJ3rSgtdb8FHciTqfJQDF0AFslfD0aKz5NAu8ofyYHed6K0BMN25ppIWKfFCvi6Ait4mA218nUAFyc7LtFKvCJuP8n6gp6i5v8h4IJCCngYCJVjbXO4sXqM5+7UOLgO0Nedf9C4IHZjR92o0zEa4HrnOKPEWYOgDoHhyi6YbOkobxyPyG7C73/xWgcA5xwhb6R0ELdwGDLk2niUroAJ6kzKuYe+7vFGT2A60DKCrk7E+0kZ5yTXwevh0nNtlXnaHABBIkNbBQGL9PFqgQqsVZYtIz7VEkO2X9xZgz4zIEmDmpGcf2Fp62T6rXpAZp+gvgEbNKINsZY0Q3Gn6noM85mButs01XWRbeL9DOFEN4LB3Qw9m5o1XPEDktQAT49dQ++xi24dt8znYnx7Rz6CwKFHckY1d++D+fZZhgvPUHfy1p2K5xwASe2ZmRAfHI/i1827Yt/as07NH2x33I8mJD98NgmWp73f6DhzN2SdBIGR15isKXiWZ3LlLoEJgHACbBCLtd8sCAjlZhDxksDdNZwNru6YJrvKm4fwpslBAp+RgRMR7WXK6yVkiW3tQaa61ATJA0+We9UZjBYskHPijLMjIM5NYPs7Ko9mPnO+qACEwBvswh/JrWSO/jqB8HecgbRA1FYHDITOKPmbyymnQeIG0rzWs8nx6dPJDVJlAQJLWM3pfsqm7Z0pZXxFlrpncZYUI3qyN8/8BLqHnrdNXU50EczLZ783Mj4+9qfrFmdEGwB/3E3kmlQUDVn/feCD7OdXrK04PRpPwk0I5gl9T19Lio56laJh966i+XYFr4Ud7s5n2uDnLT66vt0cvv+gNtk8ffm0RdXHkWRHvssyKJ59GetLFxfbF3/uN7auf//Qigs4aZz+2Pf/+D2+PPf3sOt37FkP9k3Upuf5AoOInnn5hO7l3D+vICAwdEliXPkIZTZ8D3W46ztfIKBzMeMQ+UNGwpAtYAhV+tqhR1z5QMXNOuw7d9HwoQ4rohFLyotGIy6h8aS5ZESrFb+/QvjkChstRlTCt8cQNE1CRKVXnEJSKUgdQIcO/BSpwJuf4E+wwRUGOO1J9q/MGKywNxx1m6ZVSKHsd689qLItMKtJU6LeWCttDmgWMtE5GHR7VSDjyck4ZjdU5AqtTuOJtO3N3B0Ndc9n95WSu9FEjkvKx2jMe07whDrTJ2eWP5zvy+bhwxXWiDf0PZciAMiH9GTHnh70rbi0/YGOF9WkDc9KuQLKBoEUpKPXdohZcMW6MF65ANz+8c3Zg01Fu72dfGTgVoQUvqmbt7F7llZtPgxVQMVtXPG2mnuGd8yixSagxNxcKDgCfphTZCqgo02kc/Mh6rwJputJt9EgSWlXkRZ/GT1LmdJ7cFBYYa8ajRsPdVdMKf1Ya8Y8Lk0VkdOkzEY2rG/nY3ofHFDW7AUrhHNmX9XavZLP2WXQwmdmdDNUOnlSztTCASp2pbq24iaClSdShjeT2QEXXTDuEez0wZkxc+Wdf2b7Nt4PDo7xmMA703eKwqNxY6RgMyehJX+Na8mQmF5AdkQYHdCW8VrKwnSXoZpQHUwPuBodv8f1nHED1HtwsykIGyVnhsp7ngM9rsUkG6hz6g+UgT6jPjSKBGfDSPo3rSgebotzNcRMgaKffYFVXq8izivWC4VvN1HmfL4HzCiykOkIeXk54XSKm0UFjCVbAF6qOjj98v8pCWAgKQbTV+bJeievNxM3qHZIl7ffFyUsHrwNak7FKhbZoX5XNd5IkXep3zTP99KvmLYuZrACMGFTeV50fcb4U3cr2vzpskp8PpXBex6bkHknrDUeRW4KhMlo4SmdAh1ny/RIRu+WYSrnC1PfgoMqMCgZ68NHjmCaln+LaPZ5bfFfLZdB5I1kzgBSdQ7M+cSX3NU+POi6OQ/UgAPifk1U2QkTq0gGcEdEKJEAktcsg6sXm4Er6kcOcXDTjj8m++kecmGgFnrqVjK1nsCQApJ/KomgujTowES51DQNsaBx66XyDjp2gX70edN7qPOH8LAeVRq4ysa7Hak0JHsDRXM5QHpl4/ignzMFfAZfktyxhre/rOFWOyp3ZdAJ7pDszSnRO2GZbeRg/Mxj1bc9xp3gpZYSSl/MGypKrKpPlAaEOMFhGBTI7jAjM/+U6tEX5X6hUkcn70qOTS2Pb6SWDytkFp/uE7xTJ+f/rAAAgAElEQVTM6CXLLOL8rmc5WLaDP25CaxYe4BBYKXspmpTsCF4q2Q+w9ZBhAsc1xhNnqzKU2bsU5aHgBMb8AcporQQ8CCwLwMAyKrycGDImotQa3yUQwzJhfO/E8rSf0MhatTihW7jTX2Acm1LXtaklk0Ke+ljlKoMDOvV4zl2gq3iEfQ9s2WXDCJQxPSfEhPqd2HWBnVFH455VQE6ZXrP9rLQvfqjnXvUH1FMm7IoCAMl5r3LsXpqdfWTrPvfPmR9rvdzQ3zg7LZDalu/07BQ0y9JgsMOU4cR198xm7rfKTDlARqCVeojb0TyTLzkoAyYqvXsfGgFo1wADvbTZKrObdBd+JTckEegBEB6AFNRqjNvGf0zQ0QANyYnpKb9ShdIRA15+E6i4vZL08KUXts/+9q9s56cvz8EKZla864Mf9iyJFz73qe2PPvOJUPKaNx4Zsdzf3vn+f2V74pnn3wQp9qj5QKDip575GqN9TBBCubb0RTtIVQKDJxm1KesdgJPS09SYjq/ooXRopqPntkAFlHomkIfR/OqAip5+8m95WYm+x0FbFKGwpojylpTk1HSrQ6vfkF6yQBlJJaxVOOvV0FvwbBNmSK9DGi8+27zmn1zFanxmSooL9g4gCASXh2gesu0YW4f0jjNipnBzrFL8q2EUK9MryzU4mwqYrq0OICjJ2LO5vK7KbY7b18nQcVd+CoodDiW8tHG5weOZZL8Se00twnSTVJ2vLlP7+bz0U+r0GRUiXljZLa3jlONeuPilrEj5k7GB2tiZ1h+f1wUfyKFY2t3gPEuLjebU0M5AtnQ0SWssi9s9/1CgIsp2gOr/2IAKKdvi2TQCZxRL59PEsewULs+Olkfr61FbppSj5rErzlS+Bkru17PQtStTIX6SZlp52fLAaB7jajgZkJp9G6CiASk63t+RPMWANwppDdeex5y31W+pegQaR+cIVOSyI6Jb0X3Ja/Q6LmSDrmtlYLuCsaUlqtavJwAXj44LCx1NeXHSa4YnxNyJK3k4MB6MzP4d/kGdQ0aMzp1Gu7u48oFz2u298tvMOOm2QAWkRE0KKu+qzbSLiJrPxOjezmD7l80nEqjIUlItG4+zWNgglGhzIvOaxnQYp+G1I/hX55jS6d2jC8cHnLuvDVChgzQzJxVRhujSjvWxO76clgaP761xqak7KOFYzudCRXtARQ3QcCoWAchwLY7rukxVM9jdo5VjWU6/zjm66mOz0m2cZt3YhviDg8hmMi+05Pw73e9XB1TUvbPH3gRUVP6qS629rlIEv7/WQIW4nGdUWYteXoQjrNRA58G24pj551eQp3YGonQOHCRNnyMcmH4/mu7e7ufWd/gLBK6nziHHaDrV+N0U7qP0c3nAfYqGwTvjX/JE1c+LHhSv4apQRalzbtZrkYXmuquXnZHthOxTdwxVPiSJeNZcqXuuCgMqIYOmwAIk2GPGbTHYZdlUG3JpWaJQ50msC85T9DmME4IR4ZPo3Mn9BQPwwDUvE8RIc3uu64dRQnk8xXqgAuTZUqVoxJ3gdO6Bj/E8Oe56oMJ1zArGlecqc8/Wz7IKVMoGJbqwjs6X0jgau29QTBDhX8Dn6iwOW0YOc9K4PUUNylEfHyWgwLNwduo5bmlzLW2v3KbxMtrWz9AyKMxpjnGb818O4OQOjPnk5F7Qpt2vckxwtuNq78/p5yIC6pT1EGcy98jsf6NrjzI/tzr6+NsAjuGHZaKsRr/Nye8Lv8Jcu1Hde/FMZDYSEGtUQU8+QRlai/5XaST1t9Df1e60MXr9fwMcjpGVJNBCsnPIqCC4YYCG3Wf+EDXZtns8y9x7YyDbxd5fFU2sKjIx/N3GHuyFKV392BtBo++J7weB1ZnzPzIUSvaR8wTLXtVslZBjRqdFflagAvO5imPdaYEZXMcnoAUHXAmK+XdWbokA+CHnic1LWUDqVVn5RbSj+atMlvbOZYSP49IDZ22MAoFnB1rOex5MIl0lQGrqtLb8tn/WIN726/T0zH+3z9ToXj7LCAxgJpqv/2alm6xEepYiBg+DBiD34Ycx+vMSYAykFCDtYF0pR+aybuGIcW1MMkZglftVWNLdzyXa1JZBQxqB3IDs9j58DmYsdnK1wZyT79GbQMXtlCq/+vp6O334koMVp6+8sPAyGqGcbHdP7m3nD19eREYdbccn97yvxRNvfcdNIY2vYqB/Um6pSh4jLHd6VPzFtz90pm8j6VqlCUoJfgwdvGt14Gvqec1OiCvL4efNoNY/zTHpVhiQeDgnilI7i+rGUbKM+I638jFSfdLwopNKUXZUWHoFAwpXlRIaV/7fyq+FROkd82VZIgm7GavV50PEgJV+MgHmkQMmyCjgXKGJfgZK57MJ5cvcUOd6+pp23vQm82TlEa9beDBQoQhT0WWnFPmfWUCoj7TXuCraD7pIGm3Co7oofAAVVtIsHUn2GRwkZe/qPsyACloEmjYuSUU6DttmXK3S/+qBChvroTVrMRFw6PxHh6l/r7IyAhyLAVIVjHhoA+tkeml9F+iLJasaxbvxMUugZATKQBqrWeBCRG7AER30YbLj1qK8ypibb95rpq06kRHNw7UYDr7qBR7Au1q7WsKA/xvbm/Hiqaj2fzbWkiRsZF7xCGGNuHZuefFLEuYgh1v//XJh9AqTMabwKVouDLvuzlamly/rkbF7YFS+XVF5ygf1p4Ayzs93gIr21YherjIm13FNaS2gARmXnEk+iDF4HE86UQRUxNZThjaoZ79AKltY5Vqw2FKngkI8yuRDgIrcR7t/Vld1f29u861k/mzFl0r9HsXGdvSjyNJlko/rFBqjJ5u3OQbsajNrKvgjuqnvgCw/9Gfv6hpVXyOR17bMfMVh8KeRBeOaDrTFJt0mowJnRxskkPK7coVWBWUwbRhytnn2GJuqg4mLzmd/LpyWsc4k86DZUJML33VOujZoQ+84dOfyOjnsqg4zc3pUKdHLIERyjpuxUtVWQIWv3NQIbk7w7vV91hAzUhYaxrrzwmrtsuTacMXCYF/JjhHTxUbHGdU9T/tQo1JDnizZdP6F1xT34K0EKtBPBSez6aD2PvQAXDs81nQwd/TsUqQPtT17EqatJQcZTbpqph0vkR6CMwszm//sLd9Mr8dIgzHjwY0MDGczz7YDHTqRMdVFmyv4yQUgo2UtSE9lVpS1avsoMEOR17aXyroAzXD0zcTHVejPK9kiOm9CTjAjp1/dvL8ECvAid9oSqLD5WCZAysCF/C8O2ZDLvKmCeCh/wt4MxWaDPVFkRAV9u1f223V6ehq91tw5yP4NsRaFwlYyEHtIWozSmQBwpatFBoCNzWrel14kNq97bltDrqlprYAKux5bgUMk+2uYXQkdXLRh4/YAwinxYzHkFFa5GdszAUx4DvrXQGbAd+LBMjE+OFetpJE9y5uDM7Ic5bpGfnQT44qAAEubuXOZz59xsHpBudyiv8eCz3w8zMjqM6BsXTOAAsGs3hibTlm7t2YqOTChDIri5PV16vo4KFLdghbQ4DhLY2nSNh416sbaNS2oi3MYdFwDJaBjIsLdS5CZg9tLDEF3Ua8hAX8Co5FVJZRJ2WqsOkLdROsLuYczOPjYr8mgE++nrIBSAhUAbLYIDhbQ4mMg/Tl4wSDV2kOn7i2Og8xAcr+SVzzIhuQpLyDPplkk9gwH6VD2CqXy2Ky9vLCxxhcHguRH78dxPiC92bwkbx89egTAj5k0tlYO8FjmxAVK+EFuQSzIVhZvN7oyA7JkB3mGiPMZSnNFpjHBDve9KfCtYxp/J5i1WQGUFfQvIGPYZxKAuMBzAE4go3Ed42ycrKGtsfsImRn8JlAxk2aHfOZgxde2z33iV7dHL63ACmzkyoizbIu3f9v3bk8/9543QYrdNU9FLw7wHaDiI898jc5KRIJAQPbAQjLe1ZXVhzNeRSqim4tizNLXojqBZVi2CjMtx1lpJq93rjp1yfiD4RjrcANQweHn/UXJDgGCg0VNedolZv3QRvzgDyCzRVlv7L1OqkTE+moDY6CK5+eFjNSyOpVsVMyXx4szhY+GGaOJ5KBHkyZFD6Dmc6ZxpqKH584U2jrLNrOhci0iAOgoj7Jd1cAqBenDiMpaKm1uA+4LJL9xRtT6rz6ziGyqphMOq9Lcl8ofFEH9dG9153JZA9lmntqvRp7mIJfM6qNP895qlBwEVNQx0cmdCtse4+c7gx0XioGihRRtpbTEBrvRqxriBr036zZZJ0W0KOrDj967FvVjzarask9Rnicc+v2uLIwr+tl959lDwNe6kBcO9xHGqmZ7LhHeM39bu+6otz7uhUc2KSLDIjTopHBFt7+hASf6t3qsRxl46b/DSBrPemOqraJDJI8KCWVUECMJw3Dby6ioTvwytGHKBeiQg9YNN0b3mPE1kyU6L+LRAfj1u7Gg90QbSq2UObE34Iyn9EukFn7pZV7IJcnjjuoXxmCwTLk/HZJJifCzplKLmqwdUMHpVIemDOkVjcoI6anYT7uBxPoP2r+9Ln2z/Pi+dZKQZ9gMc/QZ7XPTzbxW5CjePiWIhZjbEZaZTZknALgHhhmemOnaOp9GyQGgwj5HTW+kdiPyGKNPgBzrV2uu7clzfIcnz3+Q+YBvnU54Pq6u78/W+lQ3ghkB63KFtbRXAnEFVCz3oigJ2tUqm3tauLy68OaCdo0CNWy8XrfbS7klb2qhVhC15KN0VTkewknJ9XM+0XrOgmKW2ZxtQE1d1/b873lo3NcKEKKXOOepyE+Oy7jTe6p4Rs/kRxkxk69GoGJfFsByT11McmBFT73kuInKyT2d/UeCmR/WK19BvKqVRaAMOX9aukdkI4JZ2NDYm5qi2e90aRfOcYvEdb3SfaGoUw9HnTm+M8rZHSx08GT50fZNGHFhGgUY3ALkhESrEf7qgyDQK0saBWAz1NZH7x4aDGV9YTOUWKhhqVayoJbGSOCwcG/Zc/BqNrte8Vb7eaodqt9uDi8Poqh7J8cv7SI49ywq+x6jlOXszjJZaGSfUbbhUOQZGLI44kAwGby2XZH6kfNSayB0UbXJowDVuLtxD+jlguVDvLSQOzaLrdtlC2o0PV/Y33CEnvuZIEe47IXwKxRAIpz60sfVt7Jz2mkVNBsr43L/vjkdcX76HpQskKqVt3X0kzdqiSkElTBbSb3SyPuap8kn09OtjAxsK5R1sZJImgcyLDKW5+z8wrP6VGLIaMAzHdikOcoTqtxbY1+KOuGMth88B9kY3nzZh025QzAI34Pe0OOhPZ9s5OZQNyDAecSa/560sqbyhe/lvROnbWVk2/f2jNmPdArn83JBPb9BhaRsAn3KArHPDaCwdRawEPzCXEAv/UXgwQEj2xM50idAhclUyVM5kgX6CjQyx3DNphDPC3SU7S/ndLWH4WxHCSibt80l9AUBKcqW4D4BuEjAQPxSZX7L+uxtRn0LhFaACil9TstqMG5rg+wAyyZRzw+VsEZ5ZgBayjCptoO2r+qLWD/ovAqwm9GB5hF+GJ2l7F9rPGTv9HUs/dyqfhV+nIlCiYbhEH9pUkK7EL+4Qz8ACPh+IAchm50fLy3D4x763pQ+RQJwbL5+D/V8aDQWXIeMLmThMNOIPXutLJ1KSdlLPZNnYbhIHlS7wbPcrpHl5mBfsbvt2d4nx4Flli7zLZ9nVNT1nDMs1+TNjIrp8hz24fX1dnb6yvaZ3/rl7eyVr65TWyZPs8Y8z3/g+7Ynn333m+WeblxtHily6sK7wUZGF9u1pyueb1cXp9vl+aPtp599OYSUnEy1/iAOYIASiAxbdNHrHJi9QgmhWU1TGvbhF5fTIxHccObszpnRWHy0BEII5uIAap0+QsFxo+5T05y+wVRvQMoYs+sUPe2OWB5sNULL5qGoXCh7o8PXxwsoN5V/JkUYKCRJ7qto6L7Xy8Qsx8i/lKQVRLLlNxDKFBNzRki4IwIsm7khJc1FrKPH0VOApIU0u4zGsudGRo4ZafZspQRzX/yA9N/pZLCIyQ1RXEOZG2qIuBzRHEFebrQwqiM+9CO6c6Il0eThzNWCp7AAG1K3eM80Kh/jznYrWuPFqcVHVaVbI3LFR5FO1SncmzJRX1gAU+UfPM3pkqnKUJphbHmUyjC00nRalLMY/hSr6miNLrJYaNGaj6kAkIPCVN655zyzB9foTI/zbWp6jiAEFMIWrWjM/VhCDMIid6tToOUlPadCnL3NXu5QinBR3P0l7JHg7yNtx8ipmPQiTusfJgKxxOp4j3tKRYbmOW6YptWfzj0tEXjSnxkvrOVeeuIocmUgrrqp1ZRpjXMp/TOR7ndxHPXNVUEe71vznwyRnFopw1FkspxYkgKADHpHUTu2Og+AxKSnRe32kNTtxOoWzpZk/plkafftniLr44W3Mei98oUMBPGuO9pjrLM1Nvlfn7DaURnXLFlY9hglIyRFlJ3VBkpUORQis75KDhFuT+XfueOaY5acGBgvqUB7xkVjJCCOYhleSiVvN7I2MixrJ5JSqS8BC2QROVnqkECb/KSTm7Hf7hgV/fFM6LeMdbfDUVfLaiwA2pRVCawFrxSARA0qg3bYX0WRk25ULpy7S7+rjz9rNRv9KlKzcTbm6dOB6Iexk2hEdBNOuznJ7z50SW9NtO8O2kHeiPmVwIw+QCCcnlXUxu8Cy6Dv+UqyVjhEfd7Ul86bTRAlRpcSe/KFPC2H7QF2uvJdjs+XjupfRK26ECsnWzm72tMm368yJuF4ojNUjhroYxkw4+vFZsmS9XE+0abCdtmnrI9dSpLVmQP4BDiQdpCU96QH9Oazzxmk4L+3zL+qj61G0D1vzHklAWfotHl2yaHeklXNnMV8NS6sWtEE6W3y966UyKrXFmc3zvluymwyq8wA6QIaJ/4fhB37HJJ2HEDuyyK29yDueqSetdyqEdFVP1zz94o2xZ+V1u1aOa/gSFVJPvXWAQihhsfm9BLQ3pnZsUPVKelyLqI2Rj6VIx48QV3A67Tf3R4+euQBR3a/BcyYA9Ua3AKguwt60tkWAA4bFjNoCf1DUKLL9zR4xyK15yvlYyo9lMxp64CiSqBaI/RoWo/G1BB+1PAtWt7W6c6Rz+GxBw82y+gwR+Xpo9PtwYMH7gsxG6o6w618jNvcDmiipJAACtm15mBXiTB/Bp3uXnoo5AT4zkGRiwuvtW/AgtniKAMFfnfggg3vbc4I8Lq7Pf7EE5tFk1+cX2yPP/G4X4dm5OZsPcnIfwc+YKNbgJj6BaIPIdYjmoDTWa336HMBt2nn0xZ3fQvzs7VEzw7wmUr9ipp6u08ZMQ4s8B7PL+D+wAfBNTjHekRJtiJP3Cnu5aLQ5yPKL/Vngu0ZX2RjUXki+WtWp5MtEcorGV3e8XlK77F3af9UHggkNqdZ2Oel/FqhR5QnspJhbGru8712xzUyUBiEV0ScgFcBPy2YTWC6Ox81TwcmOp5XnwSBFv2aSB+K/j42NoL60YMpX+C/eY8SNoS3+3z9KH/Fk8pGsX3x+U/WLwNHymlUltk+jRJbJfNlthee9eK+rDzryJiIJZKKw75o9SiIt3ufE/aWqjpdzY4Bs4c2Y7/YGggMsdutXJYDslR84iQSEFbLgjHgqfYJtXs9GLBUkqg0+GZGxYqzD/78ejt7+Mr2hf/3H2+vvPilA8AKlIR67n0f2p5+x7dketXB73sjXkhOPhCo+AvPvBRORTkXrc6fagsqOkgHgqfCdalPEqhY7cMtvHqQtSACFd+VojtsKyLvJETCsS2HAoVL7/DWUPVuqZs1TVi17kxRmP1YZIatl6OlSkVjIWFFX5ji44a2R5P3pUSqSTA38MJQiqauACpc8exBj275c13tC6urapEySEXDmPEc3+dSlxNjNeUMdTQV0SHFFamqBBFkSTISLRzWzIYQIh3O6+Js9jJfg4FQofXDgYoWCMuFiBqBjAAAjbbAhs4XUJ7Ak7LjvtCTJm9xybzGcjg+eF2sjYpN6/OOuOI81oEYZb7qhXno2l54M6hy4PcOhgQS+gjQSoPk4hkb3wKoaEbZ83F59h5Qgb4ZpI4D77Hov4j2HeQHteNqOHgjvpK9QNqAJJOjv9TLjZCPnOE4h0LRbuepkVZQV7vbXYgGfR9hN8MhSeUnnDLc+/+fve8A07So0j0z3T3dPXl68gw5DlGUJEhOknN2lWVXXddNYlh3zSgrgoigkkGSCCiSk2QQBAQREMnRQJI8qdPM3OeEt+pUfVV/96B3dy+Xfx+X6f//QoVTp0697wkACYpq13+ZRwnZukP7PBOYtC57RpDX8vdi9clP0GXRsmwQVvasSCSmpE98g4+eyrVwRVANTPF7kxrqYSEG8jiAr2h2gyzxEV9YH651dpAHeFK3OjCH7goYzktjqiwtUZHY+SnwBZPaj0EAmUIXy3t6DXv2KwNgc8NjVCQE0QgRwEttiRTrWow1kCqXWM8sRHTqBXWiAuh/vlnWJ8HrcRy65CDb0DFYl3hWPnZZ3YcqGB3b0iL2z6I3MqIi208x4wCqBATJ5K5qtQV9p2sTchLKqhhJoiCNUXxuzwoEQI2RqKB3KoNppAh08lDra6mWUtCfBq6h4HbpIa2Qxsb+HdNZhr5gP4nbUOEtNhPh0Np6PxawD/ogrHMDzg1o4S6q12Ka5iofz/J6aUEyFW19r/uHPxO1ofXrLllr3rvYvELrKdrM+cmAGgVhVb6UZEtB55AaA1FSXl0HZwMF25BqpRUwnwAnub7APGN9pOq5MYCVbEABpBzuiAMo8mk9gnw0HoKVrxLj3UNg0QSRHgZRIU9zm4c/3xSXHUeRh+t97TaQ5TAkbAFwlJuQPiWiwtvpcWN8u0RFyaapgpaVydH1q6svFkbWdYR0MyFK1WRVHQjbVSeD4fCkdvKuWKNESGPUBbIUSMVmBcBObR/ocfYOVqC7Q/ZXBttDeiJ5UBxftQBR/yPWtBTvc4sKETKQpymQZeLhVmwSiPl4jrHC15wWBnWVmEwIud9jW5TkWCLAPmMY/YMD1NXZJVEjo0Z1CgHA53g577N/nuEcDL6jUHBuU/CwM0nDY8Af9fo25yY7r/E1midfneuEhLA5E5BWIio09ROcHDWCEHUUNCWP1LJgwNMcIdUDHnuDrgmkSYRzqfZFx5LPgp1dXaF+BhO2fb29SRFqbQ9SexmeYk6u8pfNkeAGkioIup5rb5i3fyU6wwPTmFzuFwB50SzBnuKIHq0vwUSURFwMaNSJECmc7tZS52HtqA6JDiTQWAKAO9wE706jc1Jxk8g4I9DgcIo1ze1hUgoyhrRCNb2LvUWmyhHqbNMhioHb7iP6EOGH8eBnyHv4nDFyhIx1f1+/4k3RczJf8QlBxz+iz97zH/2M3jBpT6T9tqZCZJWkKNJ6tlECoIMtAsRFayTklxEKcrURlTUyODmXRaGRf4GwCQQ09p3KRECPKrHmLB0kR8gKoIsu9tS1IyawfiGzAaNwtrL8Zm1RUkF1Hu4J5CkG0O2HuqxSDFTfEe0U1gesI3gtSGopX3/13YiK2nJcmu+X0EB/L/3xodupf8HcOllhymXGSuvR+BkrvBtJMewhXjqiYvuxr4nik41GPAGsEn2b1kMAkycbgVl+wZZ2QEYKiOeNLRgeGajwlxIVcLvKyQgPjqNVcUNsKmU2TGCkyHUBhLdrC7iDFJDl8DcUerTCUgglx2bHkUHqqZXnG2ZDo0xSeKUYlFwAYcpEhT9wRFJJDxis4HSj17nlj6Z6sAJiiJyRa7V2HgwKda6x/LsWlqo5KUeaBwobYQBqEEGhhznvRZGCVktBVJhhJGkP4mQaoItvmmCgHnbDDSFs2hv4+qux5TWiIohLE9aJ3n71hZrKeLwu6Utj6djakYvydWRjbQcVhCsDNPI4QnqgiqC170l6eCz3I/VY9tuxIz88+FYiG91Lh0VUDPN6bs1IzhMvgGaLYjBuKQsZ4guSyrvcYRbD74E9A9GcRCWDlQM+okccuRtskmDo5/KEyB2DAUQ1+GtMxv1bc55MbvUpqsKpRu6SSBJb/9Eg9jIW3xft6+y9gVHxXpA29vL2GA/j5a+5emz1JbLSfH9NIkvfA/xIdGZWoyK0yTtBCrjh+pnIXrmdYX5zz5pig1P9pK/zHvh1/RF+qRAVOns15Fd/wxpHYcR4eIraJRwc9HSlmtHGIdrTgKisVcXXQuZUfp0Klpt8btrm8zHWcTxaEhUNkgKLPGsY2uH6Fse1Pn58OQ4QIX3D2yUqUrUZ56QC/CL9T75uFN+KgKvMf+Q0G4Lk+zAcoiLXBgB7hOgw0N0TEbA7goe1A7iqclkRdwDUcHKArVICBk1ShrFwsksyRxYdv0jiLP0DC3fke6EDU4rPz8UVF9VYQexLBryLLrGIFvWW1zzdIWIgzJsTwvCMSmHuisKuE5V1W7Y2phWtlcxHg6iAwHvl0cK5CXOroJ6m9tBc61l+/YL9orKNMYsbRmxTawkPZ6bwDH59oZqHbAgGEjbFtYYnDcPpL31YiagIIGtdczSKnid9yGq21eYa4jTctSaJUuxMFTxiba2qDDoBFYcijY6Qsx/ahIhU+SW3pQROL9jXpRgL7ZU/z2gL4jNrREUxJRq3K6xdPSspua9t15onCmT6FCRCaFiKkAgYR9srH/u478f9XCIiDDgvzVUoCm56XO2HxXJe5O6ingTSQOvApGlLeDrgFY8ULXwGRToZfYeL9K4rlTAmCp7GcxE8luFoh0UiqdeMCGGPZhRrFiB48WJJOSUe3+1MNvSrh77UIrBzsWEgTGZgnXPfcT88wRWsjl7xOHtwmhj+dIwaJaA7qybuO6IskJZZPKQljVQkTZU0iGmcWC64jSGaQwgXZEEAqBnrKUgWDO88wMvCUtOC7AjkDPd5kCNjLO2Spb1EyuEknU8g0JEmW+sm8EcIHdSb8Hao2SkSLeCAapEBS2kla8hsMm43X9fX3yfz125VmYcAACAASURBVNnZaemOuLi4plgSUbMi04h8KKULt5EJbRPcw0VFlOQe5DWiZrRtOtYsL6O4YDdpoWd+Psid6t6GLBpIhW0XYg1ALiXd2sBgmFec5yV6xaIOuP0coZCn60qXjY+cjroJ6xnkBGpTIFK1tLkEgsZqusg8M85V2JvwFUcM9LN8hmtiQXCMlRAN5jUWIp/yAWzY6BZh6+ZQbFojHrTGQ9lhlH8TwgrRXraf6/k/S+ph6eCaZo9tzgU7EW0omUpiDXkiwt7tz5+2qYQRSOwFOFNYgfAojzFS0Fsf70ZU1FbiUn+/hAb7++nFx++l+W+8lDCz+ihV0lNWWJsmzlzxXZJiqcbXRHyYERW7TVkQmD5sbLKR8abp0vuoh70ymXpQT2sEDJeoyAmJBMDCgSljE4fqvoa3FxCl0unHDgEIK8Sil43PUujEQ3wE25ODitdGprv04KObFo+d5J5D2iznDSTvEZJAQ/7wt76zFmLvQrVtwxSj10CJBOxFEWPrZxL9smSEhLeO6uySzY6jQTjkFXPNhlBg9q0Q1cBAX/DY4Xt4XSLVCd/X39cnxikbeRJGaIW3GsRTwKwyVd4oUq7rP3hDedA4AHEBPTZtkR883BYJzyAHtgUyJciHk2Vgu8Fl1KTP0pw0Dkb2c42oqAErgXyHcLc4YOslpcO/FfNznlThAJqED6bjA4MwlRv1khmqOcMlKhpnQTw47vWFuUtXOsKUF7uDew3QxJ1CVGQy40Frv95lVAWwz9OPKUEJD65ER+iCzdSNjm8JqpDxkgNFrsWcJ2wBoGw4ytiBHORamIfgVpXrDj3IJnljwrVoa56jOqZa0T77NhvMCcIk/JjJVtKXvNB3U5Pr+miad55YrMMFpisKG0Scc1dwMicqTAJ1/q0NwyAqchkS0N/2y9ZtDatL3xwyiynh3PjU0bvqa4YiKmILsggb0bn6QkhSMJY9DpTtZbHNlc3Wxrg5x/AQ0ieoHKTyl8tglagIICIGFS4VBdFKOlU4brUAhAPYYw3DISmdN+iCdK4b42Q6LcxXba6TQQDIZO9gIMbaG9IvqZt3GPVcVv2BKteLBQkMcIOsUnM44KayltVnRdICe3bcu+t6sfSuVNtEz+kQDWDRqLUpajWExb7BzgwpeSLxM1T7qms1s3P8GEHNtQRo805kNnGtXf6Z0i0A3kj95ActGB+pnVT3Mi0ppxaRFrntNIzBrIG7YRW5zYivBZgUFCn/w3tKZu+ErEtPzJMTpgiABPwmt7p0MeFRyT5hnuBhflqQxBXbToG1stSWHDi0neXBHGr88rv8XKsHtkXjFl8QI3Vh53pyJzh6ZERFWWqMmM/OeK3bzy4P3hlCAfGYBit9k9ptVuMwtEnPs7LnFjbbpSUq/ETkc1WaU+iBsh7CHijCKR2VegPsPW5R+kJUWIpJAb2NvOFrJZ2Z1VYqTZ/2mc+cFj0PwbcUM0V+XMBlS1kD5zNrC7cSZwXNkY+/lVCKpqHVfDLgOQKkIx3QGiE5kYEhiAoA1TirS9NCVFlcHOhvyVDiseV2c9olPvPy/Qx+I5UPp9QKaYcYi+JULZxmidM+MXlh8yOpV2xs2NET6XhkvzIA26fWwdwLaMrNhs0YIvUNdA1rQ4FIBaX1rIdUN6zPkPrFp7/h8zn3XdIwhbSuOgr8HI08iQUBuM/cv96FC4UE8ftI0BFO5+B3EEywL3gs+XopQp3NYbxHHwRdLA6cIQsA1rDKvpI6I0MxZemTkTnad8VOtF6DpmgK8uOINbnGCmGjJgkTKvxvmfsWC5LfMTDQL+SSRBNwDRhz5OXfhNzKCoEXH5elfsJ+ExxYpV6JphsTMipLNQVQn2WeZYtljT8oqF0ab4WH4niDnBc9L7geyCUlDLw+932QvTaTO2m37aPYK3GPHp+U0AG+xb8h5SLLPush2M4gFmq2hzuOqWow2UK7Ii5nESOVvRZjHWxeyCjWQ8gsoGky1X7y52fdf3BmQ3+9DV3bw3h98bwq+ahp3MVuD/ZnQe2BZOQXWjvE7rZU7CA3efx4nFHnRs6i70ZUlNf12/tWWdwXn9A0UIsG+kyJjaT2zm6asuwaNH76cu+SFEs9uLarLAVRwYA1K2Eo3bChWi7BsDEYCO7P+k2gqY645KBtOPj7gzWMjgBeDD0ADaJiqFsspQA8WWTTs/B4eIvw3xKuGQ58ESSIIKF54NkhHmytKF17hw/HRDEg2XQXaeErOerbxqzNbp5ESkArAAfbMWKPWbfa8+RQgfQ55gXJCrKvr19u6+waRd3do8VjgZUmIkn4fg5n5X5waKsoVs5LaXk1pbCYeEZw4Vz2omi3zXMkDS7mjciBpjauoc5FaW4aIuMO0Egl4zZeVRT6oBSScT8k1nccUw+ARnsqBZIZvG7Og29k3mCxlqtSl2zqfkePu128twQi5ARNuDpLX+VTG9ghI20UZNiPXGy3n7cabzIsosK/1A2LGic5p1gfN1kNLijAt6l4IFNzvkFUFEUOAEOL1E/yfuMkInnZgqjAxfZCrycCeBi6ayCeGCyFMTCwJyeA1ZMsHpCQjiyJCgkypgedsFL8ACYp19LUOyIdWTuDbrIUaCpBsd0KV7p1K/+M0VK+h65FIcd3eY6GUuR+vWeS7vaRuDa1EC9O0woJCKYRI16cZex7F5dcU+MAQADQXls7pbUoPWBjub5tNgdBZGY4Y+PVit4AL1PMnu7BzZfDvzQnq4KXJTSv3apiljcKz3X60S1cJQlNOpPnxHb796sTZQYLYRIz5RB6lXfNGy8lv7AKUILDpfSE9z70tnG9rWuno9OZQoeH54Ur9xZIQbUJIlERIhucDoLuaDgNBNvKF9ptylNYHygsbnWd5MBkqS4xI/5MB/IC3ykwUpbXWkQd7pU9yQEurSLwWu3BpbeHKA0DgfiaWg2AguSFRyJSyet7H2mSsD1YJpXxaAzVEERFmCOfugDmi9igsSgsxEjt3lxXm2d3YaBqqqaav///IlGRnBkMcPN5p2tt8l6jsKe95gN4F/Z5l2LHgzgyaiac2AkABFdVcsVwAXjdcDoQGSk/LY0GiJPlgZ7Sei/JPwBEvD9Gz+dXK5Dlz3oYE91PQPCZHWFATM2y8+cZP971Hc0RFW6fiMBQU8mHNRnSvsRzEesJP7wczR6j+4a3r+b7XbLeS2vIOQ6VNG2Ua516IbEM8EYKYU01qGlpuFYEjAaNUBi0PjVHPQDDIVVMJC1qrnG5k07UcdEJQL2jSZzywl7TcCzTtEPIw8/Cwv3QVEhh8w4yJGfXymbBIDE8sgWvsNoUDAJi3SOLgURGmNc2QGzGm/g6Xisc5cCgH1IKSaYB3k8HObKhTdINyXOtGDQDgwz+S557B+wq3hiLaosVzM8dHJRzNY8NQFWe9/7+PjkvgxRA/QIFL2NqGAVWm2nKADhr6huuP6H1S6R9HGnAHvecGqhfMR3uh6oTSbQp7w5gu0Xy8jMlsiZsC0qCaOFfc2ZCai6r5aNkgs6f9k8jTSS7BBZXgTgGQBvPAD7y3ZwfxBl2sThV8jjiXeIxL8BtjN5H7SH9PgLL4lRhbROCZsQIGtXZqWSKyWsNWA5Wq9UH4fn2URMAvUEueNC5qGeR8sfqsEgqJRR25ropVrNA01qp57/2W8kzLRIenQh9avZcf6JPCuqjHqp3pDJcyxrK1wfwvJBXEHrfE2RCDLkUciZgoetwZkYtEBDhGHv+G4WkEd1S2ysk3sqfDbJ9ETVuAplSUd9hnfGzfMQEiAqHN4p9ZLYF2uUJEb8z1/YvL1tK3MTaoawLhbQVQeZoDjubuQcH0s21CxE4THxwf3gd861CCJkqlbl5JxEVPPmju0ZR16iOkBdxeFu0XtXbP0DzF8QNIr+Xnz9hbLcM4twFvdQ/EBeav5YHvG/Bm9TfO48WcxGjzm7qHjOOurrHitJj5evz2A3Vxva2kTR+bJdshgt6B2hhX79MJv89afzot9VXFpq58/uoj/Pk/a//mLQPk6iQYtpcnGjESN1kOIWR/Q1jRRVTLNAXoilCugVsqGXQI6D9NnZQPGDOA9ysp4CECR7WcMuGXlZ1JQMSCkI2Vuu3EBXm4ST9RYi8GFasWDQPnLTQeVJET1qfZ9PGwQx4ZVI5ZDEqJFY6YMbFw0MUZtlshHGCsYhzYX32h04f2u8OuXgHNlyEmYpBY8Yjnsv/ZWNHrkUqsHY1rtRI04MU9DlvoupJQVLmmscK4aJa36IAAFTwU930fL901BUHc4XGw2CozOh97t9+4ymieuGpdr/NLSI8Godtgah005Qih/Gj66RyTM1RS7sORS4j4aLv9+CJClv6pnQ96I9CMJEW4ELedBimpeu9HMVh9B5quTd9fEpOVCSHiqyvOchZBnJrJopNKUTBdyQBofMeomive25i6UTLBxKgJrzvs81vSK3ictEHZLU5JsE4CW1OG58QF0FmyzozeOW5PO0sDOrNYvVS7L/akoLucMW0Q5QJxiIUjPcABHIZJ4OdDrD9Zasl/FWSA5AnYSZsvwh5UbHywoHMKQU8ubV4tCQIIwiOAxV79vjDjHr8tSIqcu/IpDk2lnHNqRLyQFGyejNQHoub993Sp3aQUiO2eEv1yyQ0GPLDBRA5tUSFqEiXnOknn2c1zBG86/PX+9GKRRNtZVsXVP7jGTNdD2WMLz63pmPcqTtrlK36bK8IF1XkTe7C4cUaiwNrScfG6ckfqL/IboL9WcSmGgvjFY3dG5/pwU49mNvT7RIFcbG3eRvDp40YjjDF6/XwGj3q/Tt8ezxAVlsTrYgKtln4/zRdRPQmLZt6KVE6nNVRIirQ/tL9tbYGINvrfR8xE9a9i9KryFkCoKIRLfe7omuLS40SyWoUrF3Ceebd2sW/a/qmVQ7p8jgNZ/TjNbDtqne5Re5BMF0MCnzCSaiWRkJk0XLXiw1r61nk0nkv+jXp13cADnDmkYnyNWparN/M/girLWNpvUgUV2Qrh/MUeQ/gTs1TFZ61taiEkk7T4fbetwZaxwDo6P1purKyscnXkfwYSl6UqIDe4asjppYvJP4bkSpxb1FHNNZb2V5r202r6JZS68Kad3ocZ8bqvl3pJpzVdHzTvQ0gN2orqE5Vmx8pfFGo1Xu5+1dBDysoqec3XFuN4XeyGexkSZWmKZ/UQUajVGIEX9xrdHzUrub/AUhEH5GfH3+HNlbqU8icGyGAdFjq8T4gZ1XYD5JauUAyyqhayjcAzCH1DoPB4iHvC1+j1zjaoYh5tE80ykXnQ2pNWHou31dusxbLVp3LY9cxSotzo0Cx2hVRvhG5qI74avOntqzZIs7W1PGOa0oLabcJdiHAsV0LLYW0UnwfxkPma4kVkkaKZweyi3xbW7kv6okPT3Ytpq1OO7BD0ghZANcgRJloQuoxxVyMUEENFcvggaLZ0BcybygGj1SKzokCcx0HDUW5Y2otP0f5ssT6RdFsrEkmupjgSgpQW7RByb6BjsDzwjVIVWR1MEBE+vfJuue9zWqGQFZl3Dn1k6UVC1gQ7FPbOLD21M6MQDZ/r5EplsLbMDCtOdLcdbyO9r8LdpbVxGxgIBKpxDVGOsQpHboMe69tAjr8OU5ik6L7E3RiPPdIu0y3AL/SVGJlwyoQFWGcrHYJUjIz8eaicrDKAQP53d2Pkp/3fPzwt6Q8sznj8UCKOczLyMwJF+s4pGbGOR97amY36F4a69G8o4gKVrB/t8fG9NE9309tWXFkv3Bz0YVw3Hzvk/SFH1wV8vmlGyPR1Ilj6cKjPkLdnaPoexfcRudfe18Vy9N7I0jR0d5GZ3zlAFp1ual05Jk30JW3PVysCp8rmFEdbbT7lmvTvx20Bb3yxnw67DuX0nMvvCbv7exop1tO/+dGX4fCQbhVff2D9NnvXk53P/TcUBbV/4Lfoaks9Eul3gR5UIDnxYsGaPFgHy0a6KXdpi4IBo9fdFDkUEahoJQw7WreaBFmSzHivPTSQdBiPJhhVZC6YUSiQjSV6Rg9zHFbGMjv49RCQ+YBjEQFP5e9CNiAkeJD0kZoNNcybHAWRiibiiirtECmJzVgVHnjSjFqnES9oYmiQjpO3I5FKBzmjE2v3HIdGw5NPgzMuiD3VfLxNdhg120eXTXYYz9F0QejQ70PVPmzMazeMsETwUJheVOFTygrXvFw4QJYS9QThI0QuW8RanLACNG/1ZhUuQhhxEJqqLELDzidEz1s41ClHg5KYqqHi27cLGdSYM7aj3ZLwW4L7YvpzLyXgckeDq3sYWV5R20XDR4j+DvZZDG+NoGQGR9+GS4Jm26meexP3YAD4qF+6oiKcaGcSTtscakRGR6khdb9PMtNICQ8gIUDaJlMxgHMy7/2Lf00gByMh+vqcPkcz9BowXgvxCno6cwYi6ioGCuuxYHAlGGIew/GNZkH7XhRjeBL0R+YHzd/+ZipE0Vek8CNnDJhhZQQLrQEGelcDnhia8d/5M8sosKrP3deL3Fp+p0f2SjB/pfonRijkuLYRlA2LpEIauNAoW8BiGf3JI3KU2fF+c3wmUTTeZtCf4D3p3dSj+PKemVwkPWX5sJV3dzsQ24Ml4sqZ4ujxZ/ioQ/Q2nXIHxJwOw4/OmJD12FpSWgYeBfm2Y25BydRhLl0kPHtEtDQ7e2qjrDPRL1k012vp1Edq9K6joAC1i7mrAy/2/UA9Bvvcne58ZD9SBwZojlRmh+0IbY0b3PWKlvvXp9W73A/JA4YweRTDYQCi7mubZ7hTNeUB8o7KAbbLIytAwhMPUrXIwmpLdTtPNqMQW5t3CvnSvlVPRUhQ+ZpXBXooSz5glA5tZ+MZ6JFvK6p6Pjk5Jq9J/+toaaN2AyH1TIdUpmiMsEVHD1sD/D9ka2znmK0tPTEXnQetljT1YgKBlnM6QlAioD+FolUekfoX12hx9sKgo1ZqrVJJL1wwA8PdbYTNAquT9a5Awuwb+EZxRoEGZVenUeshzxSy9tzweJujqBuVUM93Q2hAxPjt7U15HWs85jGWnSmiTwLabN8M4Nt7OYhXypZ++OeiBSd0YnNqwGkcoo2ixEVpqxVBvW9UucBylYMawN3fVkyn9u/MqYM/bbaW/1ZGvZzlfBzdkZq6cb5DDUZWAaCZ7aeayI43EydmA5xdKJAt2oSU1RbMp6RgMCzQ3Fs+cIchYxcFe99PvPzWdJAex5/T1SoyPi2lVuFsxvfH52z9LyKfTkROUQ+OE9xvi54wvvUa7LPxOiztD2oo6G1QvABJiJtGTFCClVruhvk5I+2LHRuAGudRz3OqRqJqPul2nmKHehZ2Tk2hLHKx0nXr+IzStwH/RuICh1rHQNOma17ttoM+h7V1SOkL3zGltoiljKIr+f75OwtnuIDArwqxmM4h4wRZ4zQdFj8fT7fGENZi+zIKaQTR8woiQx9LRgRinibDgme5TzWVtQ5ePxHoYwaVbJMKEAPUFvVZV1fiiMpYxwW3QA8DOOJOcdYAkPhdmg9GSUZMB+Yd/wd9iNH0ECOFevQtnkSQ9L9cKF1c2xCOji0CesoCKjDuHAN2otni7jZDYHUdqmW0W6+RmpltLVJpBH3DcXdkaoKcwC8D/1RUlVTPkEmmHjl4u58Dz9P03IpLqQRVxw11i7pyUGO42whWBOf1WQ8uD4ME3I1ZyntXKPwt8dKsn1ISDA4K5tzA2ye0sk8v93/rbiArl3FPNWZNNFT2QNqe7nIrK9T4c5/CUbzToqoYIXwsb3eT5/YZ9NghEqolyO3MtwrObjcfO8T9B/fu5IGrbCNH2sWqF03W5O++g87EpMOf3jpdTrgP86h+Qs5332radXfOke109mHH0SrrzCdjjj9Orrk5t9qGFqLD79z/+3Xo389cHPiqIp/OfoSuufh34f7+Jl3nf2pEIIIRZD3sdT/voFF9KljLqG7f/vOIyo4oiIJrzeYrKNdi2vjwwpDAGIu0mTXBKLC4rMAMqfThHlTYiIqeGXvPSCGf0vRJ970OfemA3C88ZcsdKtRoYqAPRa0eBWMmXCt1w/+kOoNVhAbdlPpnQCI/AahCt8dajWTpfXRpYoI1zUPBcMhKtAe2VRaERVekO2d0cM5A7g8iG9GIBsNbLrwJiRkgBn4ICR6+3rVE1ktK1PERCOsKLt8a5EnmEdm1nlD0ugSDcFkg0Y2HCsyzoaPvFvyvmukAG9uvDlj3Fk2ENqpu5B6imqu1jTfIssDkybanlh8SEN94aImaErE+ANRYfcJ4M+hrQhXzkA3OyOGSBs3tQ3AW4ernO7H1hXkCHPdiqjgRwHQ8WC6HBYdUeEP1R5MQrSTElWtiQoxfHFIMu8brK1Irgwt1+lGHv8qA2k6VMlTG4d327Rkc+GWlD3US9uH1t2OBwF/qFV5i2/Gv+JBN4LFYvQWAKsETMbBGURFUIDDICoMfJL2IXTVt63R5UKNCjcAPiioDBaWlCWEVx8UxoMLFCfjpL9oCrV07ho6090nV5uBkOpdNwfhn/YON+ZpP2qgS2rjGJIqBqB6vehhRvMVs4eOa39BFlTNpv1vYaZUfsqKrVtxzbC2MhIj6BQXAq9Dl9lIw7C1IrmZwm4cmo7PcIgK2Y+y9kiCoBDAks9HqwiCWsNr67qw8FQCC1iSgW5yS0lGygIV9Wz8HQeQ5qR6S2CId9jNtR6op6Vd5B5VBNbtOt0btf9uSdWczRTEy0hWM4mCTst1RM2O18KpCpIIoBTSlVhebjfmrUiKCKTFkYkEb00+amt+6Vdkvq95MEklJ5mM+gtaNBXrVXRdRvwMt8Viizcmw49DvmbUel+aj4AHyFNteZL5/tqZTB1G1JNX+mZElQKq5Y+tSv3R9sXku2E2uBX4NMxHhMsSUtg5Ksj8F4ZwqJio5JZWQIl5SAY5MyWq4Gkt+g6KBCsfe295TVRJpuIgRcsHQDQu07dER7RE4YRFlNpQtTny3/v9XyWWbTTb8xOWQiMi4eEfnTx8dKhvf5ZLNEtto+IXi1l7gsAPTX2ufTpD1YPyzKLziT6xjm00hSzBK7h4W/JZunXtrbNAyg2xSJpnBDGgg/2HND1eX6AuQh6h5HUo6hAJbl1xnPXzgogSyf5ghYZ1vfizgKkT0ykYHRAV6GpIG2UpWeQ8aWSWjks8HyASBQ6cbCPyWZI/AG75+lpkl49w8jKuGEyakk96EyIt0yLlrmduxlQe5B1qnCTyh+LpciZuaxcbV87Sds7Opz5EnJhzqc6pOgxKZEjHKMGI+EzPqcd0DDTFjabdimB2TAOkpCFkQQgMcw4F8C5ND+rM7f9GPAVHWSOIxBmS7Q7fgWCD2Hq2wtuaJqdOnPAjUNyasQ/GFBhL4nciG4XXU7zXaURPBKJDkXnb72A7BOwGKawKaw299XKC6AXcr46aWixdCnpXjLFwJkWqcwPKeZz5N8mQ4aLZMd9qv5lWt8gf9IHn2kdzcFuktilHm3SMUnvf5g97v7ZDcR7GckJ0gRGI3D+kvwIxAqKon4mwNk1fJiSWEWLcBn4Wt1P6Y/NWW3cgKvIhL2lMyJHYHyAXbI3oealuQekeHSWx5T6Ls26uxStqXPQfSNea6ue5fqcSFbff/zR9+cRraGAwBaogcIniMCEcWLRYIg1KHyYKfvD5fej96yxPC/sYMB5Bnzn2MvrlA88OKzJiaYkKlosdN12D/vPQbeX5Xzv553TbfU8l7wJRwe39rzOup2vueKTsIes65Pvf2z9YjB4ZYl//H/jZpHwpUj/5EHi/yMCCo8hUYBWdYtSQa8u1pj50jT5j3eIQK5upecOrcRHvl9ZbyB+z9sK0tvAA0/bGUG5ezKzAEIZYTKUThsgxp8HLRpsfgdfyFIaaC1Aq1u3UMI1kjB6y9dcmoeMN6fR9NWBPN6fhH8z1nWljHd4ra9TnwEOoHvLpgWDSRyiQx03Q6BUunKQb+gguquXACoR5poafpSsaOZI6hIzivzkXY5xHTpOl4YhqrKFI14g2HUNuhm5csTC55qJUMoL7CwOW62hwW7mP4u0iHn9cBC56gUCk1UjmiArLh8rdlc1J3wWgvkFKyaEcxmGcw9IsyaZfTEqfAUbes8EdzuIatUOQA8lFXuT1LiQ7pGjTcdPDREzXpvYxHzbKOySAFJn5UAB+MY0IfXAH0YZIDsPrWxRClscc4CyG0j03Aem8p5GZSAmINIQGRhfMrjfvDfVcCGOUAdR6aLZjXla4LdEdpsuCxJowiC6Q24NJF0BE/m1xUj/COuCJCj07GYhuEWhLSVQkOBt0lwfMPIEQ+poPpp9s/XecG667YGPkbhsOUZHLtwecI4kHALcmezXdiHmzRumi1WgsyQWrIJuAa7JHDY+o8ETn0m/6kahQYKSgpwNY5QfTR/ClOeYTIMWtkbxtNaIiB42kVbUDkT3UR8lpyj94KJa04NITFfV17fVWnHc/krHftnvA0GhMlnuWR9INvBIZz3VT4xlLT1RAZdsiSp4YSYRkIblNJrZZ9ZgCJ7kMVM2FHCT3Syezb/SlJdBEfwE5If+2e3m4xCt/mCSF77wXuVbEhq7S4dtD/I5W9SjQhqhvLBIxE+UiYZR0oKINmuZYa/6g0vnymrT5Kco49tnyXl9qLYiKIIcgy6sAiXmCOg9WfYblPc9eohZ8mhYrjGvlHQ2M1p5ZJSpqzJou6OIkeWBUbaC4opaGqEhGergCjUL17LDjwPMILKVNTrrXqq8YpwpZ5UxJr2zCXSWigu1GNWdSmYp7C7RGZS20mjsbd0+F6Gui7RvxXftOvMdTG0181a194Tgpl3smODREZaLFONZWj7cNVbRim2q9XxqiIlEtRaJi+OtaxyQ+cSix0aNY7sykejeAklKoNwXrdB3pWQsAtQL9OB/HQtHqgFdfjwDhQWbIuxqFlLVbQRe4dQuwT86vumGpQ+FiTakDp69on8doD34PagXgPOxBWwWz2yX18ZB7ix/3QGLltWbgKwAAIABJREFUc2fnBDvr49eo45rX6zJ0ZJnTqyM4PZXVZ/DFv/P5gkRoyhpL77RksTgtsqxKlIxEVnSElNgoJM54AUgJgLz8Ls3IoKmysLZQy4NrdfLZPRZ1Tm2XFFOJtgfwKE2B5qIEbc3hvkCCCcmuxYyl3okRTPm6lHgsWwySdhKku13I4wIiAesb/WfAHSSCRBjYuSKMKb6rEM4BL4FXv7x7kaTI0iwWkeRpRVAEvePWYiAKrf4qHAcCQeEGIkbyGDjuslTwb9wevo/rsEjtF6vlIjhNVjwc+6ZEh7Bzqj0Lqc8wXsAbEVEh11stFnFytugW7MtCJBkegfmo6uVWyi37DdrH2yCBZHL6qWprmN5HO8urNOqnXNtVm+rOIKmJ6fY61sXvVKLi1vueos8dd3m1jkRr8yL9lYVpleWm0IXfOoTemreQfnL9A5JiiomBr55y7bDA/qUhKljxbbPBKnTkv+wqDfnG6dfRVbc/0ngPiAoWnq+efA1dcdvDS9Ot/4eutWWxFESFLCjxfotoVwCLJGxO61bwd1DuaiDAcw6GaOmwiNMqsFMLizSiAiSFmowKagrDamGDYFqRtxET4QkVBrP5LfD6b+cURAPMxGqBrHCPO8gCOA/kC4iKeLH8KyEsMjwEbUgAFNM6OqLs2aBGmB427OE+ZYu9Rb029ALft1zw/Aa0NAfz0FZpn4Z56jsNuLdDJG/4mhOS51pD8Jbw3GNT14GmxQP83UiJXulduFDYdGH+29ukoLZIhoDmarQK6GfkgYa2agoopE0BzGm2o4wXj5sCXvqr/JtzpBqrrEy6Igd4PoxhvZ7Djflg7o1n7W8cj1Rm0WbuMwxXgNbKV5hh7iMwxGHAPEYLIFa+Ecl41ECVAjCkJFcUvhJREcgGExiPUaRrRUdYCru7gqgqd2U1lwBMGVHRkFW4VKC9wWjUZze6B3Ac69RdbxwVlEu6ji0dltcbMq+tAKtK/2wlRAIx5DNW/RZfDDmMeWO5uZgfr8sS3YGeG8j1FxEVnFrHKh3jcKgsXMEcSsiwhjmUzHcrnRP1khuKMC6QTTdWcv41YCfjqVoRFan0mUZA2jOHesae5GvXP6EGWkLHRl0ciArzGAsh20JauGdmhFU6ZrX3lddU0lLLsR4BKfyqAgMCVMUohhL7Z8gchT0//uLBxdL4Ri8+r4FTUkJ1YmuiQg424rUW97A4ZWW7oA6plH/5HycqDB4LoIyMee0YgtEuyUWl5wXdrzrTxjQVmhaCVfG6roCTydfW3LDnFNskklp8f9iHsnRP5abXn+N8Kv0CHGIxLd0arBNvbq81PQe9JfYMdB90v0v7N/Rqx3YW8303xrr0kNrmXKxtgjQeYqxlT4M93Jy/2h6AVKGw5bi9IZVHccg1HSeDErpWrJBxC6KiZCOJ7Fci6WtERQ1clt7WEIAhSKAwLgAKWF8XxL/ie5IQHNDh8l/nQJLoct9WH8mRkX0lMQldHAp1rgiqgnT5j352ChMug9H8fmlTjNXWjp6lmtOn6jcqKHALKqdq1cV2xfRPwTQVJzt9hjoxxegGsdHhfFS01StEeyPfuBvMopzFc1+1/5W5XFIiKpZGBUrfow4eSmT00sWhhCA0mY6bpg/yz8A5C57yALBxDmQvfKQQkoK+loaoejQCQGznsHh2Bzifp05q7s+wYwR0t/1bgGdJqaMgthLx6WywfPD7AEjj3eg79gd4i9dsG4gAng8pMgkvqii9NiXOtB95Cj/YzEoIJ/sbn2lcTQv0RQo4F4ooyxvD+V8JC1VZmrFA6oVIZAKTBLrWxAHOzt2qwmKKachALgsDg/3iWMrOjkxYKN6gEXzYa1X/MgaVR5zoHAVCORMcYAM8qHCeRAoybgdkrqHtJPMCpzpSR2zUjvD98VgNt89Hn/Bv2Ps0ZZZle0D60Eah9NgCeMzr+GoKbX6e1D9BRgi73Gc8SfaPjCjEb56oUKJGa38pFhbJF77eExU+zRXjauII7MYvlx8vd8l5D/2wGqh8naZo9zVwjfS09FfAJVGfBrVPWSLEMdai32ukQE2ntvpetw5v+Ko8sjMlY1ueSK3ZkLAZNNK8qZT5m0B2ZY1pRVTgUm/PeHJcTuHvZKKCazDkERVvZ5K5FsQR/7Qz7bDJ6vTNM26ge373e/rREX8jj9rv82fRC39+a8ioiuESFaw8N1xzWfr6P+5E40Z30vHn30Y/u/HBYj/eJSp4A2jWqODUT56o8AtM0u2wEh5cFApsSxqdsIZRXNgA6QJIiE0MbvDqrWqscHbgi/tMJCyUjefCU5rKSTdLLHz9LzxDJHefta2vvy8Uq9ZtPpzAbXdzjKYdppooql4qi18AwtT88CGqOVkh3iIj9FCr0RfRUPaQUAoiuwNyptzKJMbwrVJ9j6bi0M09qjwNLdSIBvECkH1L81IuWsyHTRSzVAKCPSnkCMyFyEeOlDoiwvab4T+4WFM3oRAUvwk1Jdg45fnkv5lQ4nkFWKZGDrdDN2f9HxtdWpyb3yltbRshZIqGG2o6KfbWgJeM5HI0o4mN0PZ2Zea585prPI6zjqsCaXrQsagJJmzaOBenPgttQqqYRKbMI8bnHtQ1BflJNWkroqIGxg1FVPDLvPGspmPu2RTnHHMKryZdVzXzOl0HIj8yvnHcbGGGtZUAWV6WFclyS93WsNudIdVDERUAZiOQgP5V1kXl65hbGjLgySzfVp11yZVphV5BTkSSJJ6N07lEYQkjNtTSSGQPMtUyogJERSB27QCzlESFn+scoPLtjkaQI/dy8iaITWQl0L08bdfwiAocuKKu8oeyVP/HSU1VZk03amPjFqIyDB3EkVw4HCCFSZDllkSFX+PD18toC/K3e8MXukm2J/fu0ipNiAqIlge5G8ay2wiUCbG9DmOe7kU44KeazC338C5XayrJrZyPSQXo0d2p9JqUNEyu8NfH96gOzD8GzODw3/jd3ZHrLZsszIWOef6GvJ8lWajo2cqGUSUqTJfmWk/Lo7v3gjyvRaZCDYX9CnaVS2eXdMPGsDBLwpk6MtsPTxxO/7DanhN2AfeW6I1ZFJAawlW+uEWEkJP9VkSF95xbapk1+zOPmqwOR0WntCAqsGun3QeAVVgZFcAe+yMAJAAztRQtcM5BAVlZ0ZYOqjIVKfDvUlYygFj6VImK2guK41S7ONWBARBF6oWlJSrwGlsMNbvQt0b3T9tzUUx9GESF3RYfNRT6nA3B2yEqEDkp6jF3BssalKmalhMQ9kLhE/TOFAjHGU73HHW8UQexRJTFsIeqZg9h3e5gr/OTBSwzAo4bFQrW1gjCYlrB5objd7na0h4OoeMJGexqfw2iIh3T2MKS2CgRV+oFA7WDNLJNaxXmNowSQYolCMhtaXQULOfUNbBvNDq+psaRnx8OiXo2Y6dGBtvNGc0kqpW9EtL4OBARjm7xPNhcQiwK3pMezwne3NJPTnc0UE1flaxxN5TBsTGczXN5Tw/u2r/hERWBCDegHKl2QMbVwFY521sKbj5jD/QjBZLiMHzmhi0kDqVWMBmAPuYdnvNSc8CBy4IbdLDzoaaC9oXePdGCd7CzrAhHADEy9ZGZDGHthTo0FuFbS59jj0MtBqTO4n2O0xuJfvM1TW2RcP9kTNvaNA0UTnZGYPhaEmErqKWyN9wDfWUyQVJt+fMxap7y+BuBVptDP0KBUDASAKnbcYaVlFWOXAIGw89AKjfUk8B3XGtCUm5zlIWRDjWPR9STCMSO6QWRJavroTiZObcK1qNzpo4Rmi0jpiGPNTyQzq11HaDCdlNQdAyDABPFfiYyaOMmWKB7lMfmcpzur0pUuL0U9oGXcRXQd3DqJ46o+GsRFSvN7qHTvnygLNy9PvND4voOn//bbWi/7dejs6+4h753/m3FuhZehIZDVDBY9L45y9APPr+3FPc56/Jf0Sk/u7NKtrxLVLQmKqCEcfhgBYQiWAEADXulL3Joizas3CYgAc3tDRbUxYj8Qep6i8fppspkReqx7q0Z1jUapqgeEXwvt3/UqM70MGpNgzEVijMjv0flwC5jYx43AIR0v0z7Go10CSYVT37xW3f57VSRBvWXAlCZ0vSAiFeAOVHT0tq3H/WeCEgFY9feyUaEbCDIG2hFihBBwI/BRtc2kg1DNhL14R6s5Z4vkjBRDYHkDRdpuLRAV5vlLNbCUNwsKVrlDgkwh9WDQDcuNmLkICG1KPTgId4t4QCzRAgL8RCwNELY0PiaEFZoRcP5HXIYkVBFNTC5LciZyS/gtrIBzu8XciYUuUqNxnjoSQEYkBUN6Eo8lMter7VzkWBi8Kx1RB0/GzLli/pKWzOiAsA+PwshreoMo6sNNUxyefJiqcaNEToBEDOQMxsWPKfAU0SyIoBo2oZkBHFAz36QI2UonuXStyVeEFkvijiPmpRNogK4NW7KKQc99QrZE6LKyjUqwvrQwVdD4i9I/SSeRr5GhZye6hEVZXDQ1m1hTLCWTSAsN7QIiRFhNq6egUiKt+qBHwfF4RMVmS51fwbi1Ml9nN144V9CVOBwEYgKI2xV19hu5F6gIEcJTB2ONm5ek5CMrmZQICkyz1oRJbc+GkQFlOhwmvNXICrk/bInxqKMcf/KV7Y2rgbc/G8kKnyBQBl3A1+RCi8d5kphCSyq2pxUEMzhEBUiifb/cAbWtWy6eSlTHYUZKrQJ67vUDRRMxW9lEC7dJ8vDEddW5GOGWm/Dr03UalmUonAF1MmAIewK2D1Lz6w5HvjnqSey+Y3XF0WxyeXLkzCw7D6kYWnemduzYQ7Na1XzjuueFyNYm82SNA3i9KIetrArtdBs4ZOlNMD+LnbG0kZUVNfW0mqb6BEsSwv2BtJaFB5Xi6hoSG1hP0mandSMMVYddROqZFz6lmAK/XcQFVajAvqnFVnRAodOh8C1GxEV+dSGLIlCOqiTWiAqZBsymxI1e8zxSZFx7FV6HcByBtMkUlwKuartXxTZFrtXAIbdHlzrg1xSnaP03RFEN43zl0ZUyMsRXa+9RFNKbWpFVIj9InpBz1oageDq1Mj50cDGzNse74LTVG0dBZ1jxhp0JjuWwMEO22Ar4NYX7AVZJZEdQT/FPRNTKEVsxeZXZzpgDBppoNfD4Q+1zUpyg/N1vi+kRAWimqIDDcQtSkQpEgfnsDSiQkFWokVLtDaFjpWelxlcrn009Y7iLvxvJiakJgh7xLe3a1FlybTA53MmIfq1tqSB+QCPtV6o1nyDHuXx1s2BiUN1DkSdOP6Nny9ZFwyYlrO52eQ5EI59K/Hs95FNwXy3SHhrL9J45f3neqzsCIkIBvkdKX6tTR6bQaoiT9BIFgYj5/B8RFnwsxdnafZxDaIevJOhrKc2deDk3+Uau6EVMB+iD3hshWSPWgjnDcFQzIkAZyDs2TxsnpgDceHbIcRB20iZd58SqxgahLO+Fc3m50mdCS5E39+vzq4WdRFrmqhjs0aPsIzof+EMw+QQywWcVqs1Kmo6NmG+3YkOmIg4B8D5hvEnk+HKooEM4OeIGaU3yFhjf8qe1Xo7MN2fRfGCxBFRfTeioqrTTJlpQevP/+22dMVtv6NvnHadAIErzZ5M5x7xN/Tya/Po40dcKP9t9RmKqGB5n7PCdDrqX3elZaZPpLOuuIdO+ukdLSNC3iUq6kSFn4vgJeUOqAG8ysJaRdnBx6J2DsgAFuSng9LTs3UE7vmBCDVnRc+EAyst5A1XZa/GQlDqgSGOEReSwojzRZpHFkLw+HVMbEnIooOaAD5E4zZD8TyLXyAp1ECK9yCUUz3X00N3uDagC0jb4aPE3LOc5wfGK5kz/GG3qNENA1RnKJIJwZRzj0COUDV+AmMt0W7migTAA/0B68ygt4UnKqHAG4ca+CGVmDQh5iAWT5R2Lnyth/+wMQZEQlNDKSKuzQy5CDlSxUDfWLw6Atc4JEhBZd0NJNIDm4I+Rx86UggXNdpQv0JlSg0oGNp8rebPLDjQCiirxctCKKn1Q3I5Wj7PxGPZgEGVP5u0TNxy/ajAbxpFmAAlvjC9PMsGTl7CDdfx101QI0tCfRkNx2hZC8bOdq4BKfCu7fWdwOqC8axXBLWCNZHfEjpu8FyWJi0ha0rAXqKH3MPDWsvWqaUF84ZhNCAcsOIeBfAkrO2w7uI6S9dnAezO9CV0hK5WkCesaHTuTE2G0GsRUrb11ckk/QR1kxd5dqao1cFQWgFgSHNXVrnDgR8ki0U7QZ5w8M9kAASQ14t6UInvAYEKQB4GdA6ahf2iQRDEiQmHB0ujB/Beu4c8ygZq5F21w5zqAgUOlVTyalJ74g8pKtOI/oppYfR9XvenHnC+f7rf6bWqKm33YN1kuhseiQ0wMfBjcQ+R9lgIvR72sn40p9mWb+yt1rGB16nqBm4jIiJVbiCtypVhvOKyjB7wbmQwYrVWFL/H/Afg2+XMDfKVsWIiuzmdFIRvCIXrPN25Qf7AhgbKoaSQT1v2CfHwjDWQPBHVquMeYPEmh3csiHsjCHbnZWgerQ2C0gABTbkID1duSSqj0NK612mdKF0/Jp9YR0ZGNvri84FzJKRpfX9/uo/V5yGnsqC96uOnz2roqwaoaMCkXQvZSubVrd9ARmde+bWWe3UMUsc0uI2G2guaO1tTPIR6LgL64sk1miOOQKr6Y4viesHSxvzxq/M883aN35/tFXh+iCBE7a9KpEMYQyPyTHgisR/2YWf3WASvyJmzhxLAN5l0S1WB3PeyyFXfalCvG20TmtrxJP1e5ULHTiOLBcTOUjSBpNY15m0MJ6E+GCkT3GpbQhSxegDle6FuSWWpwz7hwbJg/4ZViDWt8oc9V21ibx/GwQ6mRACxda8Tj2eze8O7LYI8X59qr9sgiF6NUdO+bpy/LwWacZpycu8G0dvRUd94PeD0grvPOxsMWmpajJ9El1uRXsiEC8vQtetsgWjHxIhCv0pTGy2dQyVArdajaQixALm2nkWuy/ywrnCOVkHXuQLUsu/beYmjZuGZHnWcjpYAqbJhRwMy6lvYm/G/6B+ukWF0mytS6sDm4utGWq0kgARIZyNn/EUMei/W2jSwwXkcTEwCBmAEsQcAA3k5gsQhjsdFndZGUBuTUrYueX59ZSQ0F+MjERmMEzDxEIBJeG9rHUb+IMUO7kdNDC0graA9j6fUWZB7JM+S2TnQESaZSaS9ji8734nDFGo7Si5/rauIlEtI1ww9rM0tG/5yNDD7AzqDp1nT9bTLGMsZ3DCUqKNVDGUuGUxWdwy17dxIYhwAoPNlvI5Rr0O0lJ0nBdQ2EoixG45+4e5y6iGJhBEAmpTYtvRbPK7ALxin8c5xQbc7pyHINvAg1ELgdoZ0YzZaAQfIziFe93inVADfqJ/h8RAlgHRFIGME2sLv1XerjCjBoESd1GoaZCIjAu54royp2AOxHiTfi4gDnYqYUovbwL/zOHEbUNdBxtCcL0MqLSYBuDC4kVSwUTWahck3kycYaJzCyupMQdfgbOTXo6TgNuxHyMoCCRPsCEsxL2nFBnn9sUOopsdSsnOkEZ2aLh3jL8/Hucz0rnc+DVFNNpFIXYV2p/tJnG3gQSB15HpLzSXr0RqOc4/WRC2nc1KiMk2fL/MO5Y8t0GQXESyjLGsM9DvSqclZUxydtbL5IjVIdIdwJIcce1zN0XeJitwCyf4e2z2KzvjqgbTa8tPok0deRHf/9jmZJP7+uM/tReutPpsOO+ZSuuP+Z1qmf2pFVPAcr7bcNDrhP/ahCWO76Pq7H6OvnfJzISmqTBQRvUtU1ImKBPwY6vQli00XCwzpmhJQ8cjRHic00F4eFEjrezUkDgpRFLILVWuKpgLSunm1CTnBHgEgMFTRJtuT/eE3f3fws18B+CuolNUOSA4t8dnJ4SKcz8x4zmpTlK4NBV6hoMJ4WVtDM7VN7PWguSdNqQGMN8MrzEtoogc03QSMVAY+HvxxHYB/GLJDKIagWDUNFitizkcpJIH9XwrYuza4ScJ4RxBRARp/mIozVpC75EyZpfLKfmvyB15Y0n+HLP0utBljFrwIk36wZGJDiwcbGJgYTQ9USS7ZIDtDj7eeRCHSZoKIOPhDSOlQNZxn6zV6QHUfA3udGQANENoSvaVqshONP/Xi99WMdZ+uAYTNludz5qXD1p+Awlb0ofGAmjI0QjT2LoxH0Is2MjJG1eTVTkc4vRCJCp+6Sy+Aocj6hw09MVQt5NwtZ7+y47+dDPIxBB8QimIGiW5XE6l4ELLQ/cFFA3IwkVRubLglZyaVKxhoNtM6WrJG0nHl79hQZp3FHjZ8+AwkZBDhWGcmkh3upBy4FtX5fCjiw5DUVrLDZHtbh3pKVQrZWQNLwxjanhMMMld43yBC49uI38VRWBIJBsPUQtBSsgFyaGNj+pbTB/D/EPLMh7qO9lF6EPb7ZTLuSnDJwWZggAb6+2UMxIivhZpXljvkgw+z0Ls8N1yLiPsmh6xABuOwbQ8L5KLbP11qOhzm0v23rncAmLOnG8sdPBd5fPl/QuIkQI/pJ3l9hCfi4b62rvMoSX9dDgpAB6btZvuC9zcef26rHOLb200eWPYq77bv+ZAEj88QDWERbHzQVbngNafFBVUm2Psv1nJKFqM812R00SDxGEoI/khdbzy/TNhHb1JdZyx36AP3XNIa8Prhd4kXaaUOhpEb7F3JsqeHLz6081zxuxjIQei8ES2FqRcZaQAxTY1UlRo7bKdaDCCrggZ8oJbCp5JCBKSKknMsUwo2cGSoji8AmNI2kUhKcOhhqbQc0JZeRmRZZITHt19yHvNI4j0SxSxDGyjk1DshB6qTmjWYa02Vyp6sYv+O5DSbWCusm8vplGS1uHHD36pvYWsaPVk9bKlVsGiAC4D2K1Bj4JfIgIylpkJFL3WVltdXE5g3WV48KPpNQS0dv/b2USJjuY3T+nwCYkJJOY0A5n2D/2eEL3ZElgtZB7wGsHag31Ndl2qHmr6JfYaO4/7w3GlO7jbi6GVepyATamk1sG9rPnSLZpExjo49/EzVH/0hilh0aMeomM7S5zf3NonJrewtvLfa3PpCtXUNrr+IRAuh1C7e3KxDoL9TSjnTqTglFEXE9k/3m+KHqj/0ndFuBMDmLUGWz0WL7EzrIudBVIiuMFsCtfX8uUUBR9VtPF/qSR2J3dCbzEbC93AegszwuW0xy/dAHy1a3K+6kwH5xUuofZR6IId7LOoopkVOibZFAwPUN9DHzICBjmooKUCsaXWFUMAgIbWpObuFfomzoO4x3n6BGmDHM6Ri0i13iZEI0Q70s6oA3iJZvyxLooNRfM2Icb5ezvhMrLdrJLH0PXjgL6ERbeYtzoB2u+pr1rkM0rLO0/OhpfyxdQygUdeceu/jXIH00XBgU8Q4khW5jAvgLzaZ2uORJlUfozDHZokg3Q50lEYAab/YXsC/1bZX4Fll1qLulDVLHDDyNuG1oQ/B0Q/RLrq3BRLLxtPrTZ0fI44iPGoRONDX8ZzuMYLo1GES7VJ7iR5wZzqNtkhTeiNVEuvaUOsB9pGB5/ocXcWSHtA5j8raN7CZ5xNrPgHXhdhaug/6hbvwft4zeDyh3xhcl4wkBrxDHwVCmElO21v8uhNig4tNa+cajQMJKb8YSSLyY/Ya9gn9jovSK+Ek0QaSMUOLwbP+RjQN4xNCYEkES3QAUJKP5N7wmwfIQw0fl93AnLwAwIeTJI+DyJvaWFjDIKTaAymsERYgMdnmlPm1c5MnSUAe4uwoNoTZLiAMAnnRAhhGpDTfL8+3bCxwDNN9i/9fdHwFIZZPEOt9Hk+WacgaR+XhzKY7oE2v/Zev5bkQ0sai+TRVCWcf0Rol/OEaLqKr4VRgjmPY4X1b3iUqhljXO206h77xyZ3pyT+8Qod85cfUL6GTyjbuvx1HWmxDv3zwWfrUMZe0LNxdIyp48cyeNoGO/9xetPzMHrr69ofpyDNvpAW9mj+u1eddoqJMVOw2ZUEctqHP5Ql4JYrascrV4/8QiEQA/8W7ohwKK8DcIgbg2VBTwwEbXPkgEgsKMlGhBhY8imLxtFRtuKFwnZF3Iyc/jPe3S1SEXc7+UUjpUyM2ctIgpiSJD+V7+wc0jE5MNFfvITlwhq7agVHmyHVagHH2JtNNVXW1vyaq3KEBJxx0FZjg3QD5KpNzd3i9l6TmgRZEhW4iPmdlGnKAp8TMNFUJTbqeYwHeMNe5SZ8DUAMGE//N/9aNOBGkMOoRrE3JgmjwJVuP+bZk0hpOYCXNB5DbQQCNg1L53Y0NuOUERwBD7kveAQM0PrFGVKgHt9Z/8CC5eFa58VbvvJiKbSi931zfKcmg3utLT1SU1qj39MLv4llWkJnmGKOl6mGmHmWpDIi8G2jEYDu8bN4OUYGDNp6pYHROVKStlNihxYtpqx02pa2231S9s/5Kn9dfe53OOu0C+uNzL1J312gFZxyh4EFm23IcCG1jZ55iM2ZPpQM+sjv19EyUw9atN95BF51/BY0ZPY66Orv1MDsEYKy6JfsYKYo54PHi8Vj7PavSLntvS12dnXII+PnVN9GN195BY7rHUccoBpIVSI8kUGxvWC5yMGAPpkW04kqzaafdt6KpUyfLhX/84wt03lkX07y3eiWdodSOQusyooIPSWutuwrtvMfW0p6/1mdhby9dcO4l9LsHnqDu7jECQvD/dMmrjtGDSUC3QiSQXPM2iQoQQVtsswFtsc2G8s7e3l46/0eX0m/v17YwWC+2QEaA5akqWjmyYJxKJJL+NjRRoQfGQdpljy1o403eIzL26iuv0WknX0AvvfA6dXePpQ4hVgr7kCMqcJiLbdJ1t/f+29J73jtHRnnBggX043Mupd8+8BSN7h4rh50AZvq2mmfjWuusTLvuuQV1d3dLTamf/fQauvuOB2n0aL63MxII1ofd996SNtx4bXnXiy++TKeecAHNm9dPnaO6bP2UiAoFQrbZfgP+ixF7AAAgAElEQVTafKv1gzfj9T//BV171S+1/x3ov4Jt3gPNy2qNqKjPRLw77PvhK/WUV6JnkHomj6VNNl2XVl11OZrUM5G6uhg01bv494ULF9ILz79Mv7r7Qbr3Vw8xjWD9NqImsYOaKyzuuE2iQuqtLRqgQz+6K6262vIiV7976Ak65aQLGbalLtF9HZre0vYNEIXYIZI3JkSF6qN137MK7bH35tRp+ujqq26j6665i7pHjyP23hsp9YzKtlCDqPC7sSd/4HXZ6P4S6pk0ng780PY0a/Y0+fW1V1+n00+7iJ59hnV7Kqt+nyzpqpSo0HWw/ArTaf+Dt6NJkybILc888wf63rHn0sgRnSLLMR1LtPnLa189zkEObPT+NWnd9VajZZadTqNHdyuAaWu/r6+fXn/9TXrskWfollvuoef/+CqN6uyijo5OI180dWhO8A9H54BI3G6H9Wnb7TeSdcM67pyzLqP7fv247Ye2vlvaYupdi1pzuk8JdS0pefY9YGvaZJN1pUevv/YGnXLKhfTsMy9Rd/c4ISKFQHROaGE+uF+cOmbRInrf+qvRvvtvS11dS7+3cNvmz19ATz31e7r2mjvokYefpe7R0N/qgVySS2+rxPHEuYX3Fmtg0mAlfEFUyBVwcskFTYB7i5wx734Qieu+Z2V6//vXpuWWm04TJ46jzs6oK3hQenv7RC6eeuoPdOddD9J99z0uMsH/A8EZbNoK0RLTt+j4szx+/fC/pVmzpkpLH3zwMTrim6fTqI5u6uoeLcSyOvFoFBHmjEkoTaUyUlKpsKh8+lP70ZprrlRaWtXvGDxbsKCXXnrpFXrssWfouuvvphdffF1lPRDj3mlNdSvSB8OLOOqSXNeop/aeu29Ku+36AbfOlqqZxYtfefU1OvbYc+mxx5+njk7bq0jBPnzEpjBBAiDJ8x0AcotoCB7bTJJUmibnvMWLqKuzS+aDgUmRNeRFzsgKpCvWOeQ1xbU91JES9h9/j8LkqM/IQGnUL6aVKspFQNKgufQfateA6Ile3qG2h8kSXysAr10fTCp7V+pkpG/JSWZNkwWsXd+r6bKWSJ0LnJdFRsWWjTQlHFBD+kCJsjBbwx6a4z0AjlEYXCNHLBrG0rchCkYbrPIXMiAMU+wiARPlWf41coT0izuiDgdtMv9cJxW1OjEHfL3UnLCoAyngbucunqNaOio4ksCRBc9jQoTrYmBMAhHLsmhOGPxOIRlt2xcgXxxGBwMRJvNjaa34GUijzrqAiQrMEduOfK4AQQJ7Wew1+x/qeSJdmgmgRuJJRAUyeKgDFZ7h/ys6xCIUfJ8gn2of6lwKSWT4IMsPn4vDOdlIsJxkCrrAiEq8g5+FlH+exEiwzmyPDHumFTtHTRa0Rfsfz0aQHn6mpE+zKBu0uZ3nYvEScSpiXS61WySSQ8dOxsD920dayKveqamfbvvN0/T5468YVjFtzUPWVNtMBBz3mT1pgzWXpS+fdA39/M5HI446gmjS+NF08TGH0piuUfQP//VTuu/RP1bVQ4moYKnkNE/f/tRuNGfF6RKV8ZWTrqFX3+Ri0ENrGhAVPM1fO+VauvqOR4a8SQ43xroP5x1DPvC/5QIbDADgYOCFxW0W0w5ERcAXbCGUvD/tGvVssM3PeVuVjz5ldljXbgQ1QFZgEfqhigosRkmwcggAsUUM4B69Xv/H/1QPFfWcEOUh3grhaujRxux40MJITrvWjOS3EVGBTb0BvgbQXZvhf5f8jTKPUeFpPlAL4Xd94fuE4eewTlesyHsVpB2FwY8xs185VZAY7cyCm8EfvI18qBnA7qZwe8MK4w7wERtCcu4K4gDDENCXlyxfU8DLkM8LHmUuP8L483kJbA69aAgzxonfWQBpXIEq9b60nKzwFklfbPU94jMx6zrWifTLHw0V5weupJxCAIa/0wxL+crPG74vK9IqqOtbZu2RMQ3hzbF4OxacB3GkFdZZEBWRUNReS9fyufgfJio4dUFJTjxREX4HQFsBhqLOiuteyRM3F9J/FIRUPYA8oQjZxbnIlIdrnjOqncz4wz9frOneECzH/3IhrK4zbIRtuf0mtM0HN//rHjBfeYVOPO40euFPr9KEcROpkw+Zto5EEtQqTeQ2B/7ZEuf2bf3BTWirbZlI0Xn6wx/+SMcc+X0a6F1M48f1COiYA6RhaNwYNVVA1BgKzCswu8Y6K9Oe++5AXV1dYlxe/NPL6edX3kKTe6YJOQLS2Mt7LtRswHP+0+kzemj3vbejWbNnSNtfevnPdPrJ59BzzzxPPROn0OjuMXpwQDuTg7CGiK+x1oq0+97bS3v+Wh8Gxk8/5Vx65MEnacKEHiF80C/4rjbXaRzBv4So4DndfOv30dbbbSLvXLBwIZ160ln00ANP0aSJk4WskMOK5NuOH1lD2SS2tOOydE/pzUMTFWxjjJ/QTX9z6O40ffoUaQi3/dKLr6YrL7+FJk+aRqNHM8lTAOSMfSsCxSbXa6y1Au2573Y0evRokb5bb/4lnX7KBSZn4yXaBYBEVAAKXvb399Lff2JvWmXVFeTe2269k04/+XzqmTSNxozhezs1Okv60EV/c+hu0gc+vF579U103rmXSfvHjsV7UvCH3yeAwcjF9NFP7EXLLDtT5fell+m7x5xKr74ynyZOmCxAfAQkLWKuIKTeKWO4MowZCkVyzQtcQdYBWnGlWbTVthvQiisuM2zd9dZbc+mOX9xDDPa3jeiQ9vM4o6aVgLtQTZnsKUjKuZvNGhVbeREx6H3ox3ah1ecogMjjdvNNd9BZP7yYJk2cIjoDgCN2hXzfTKTceayyPlprnRVp7323ETCZwcuf/uQquvrKX1DPJAbgx1J7e2br4WHelgdxZqAXQIEATFSoDpZflvn1N1iNdt1DiTGWt7vvuo+OO/YsmjSR5Y37NyqmhimAXaFJ3klhyWLJg/7hQ3eiddZdVVowb948OuP08+neux+hnklThAxjD3TYEWxg+Nzc+txIXPEWs9XW76ONN1mXJkwYWyVwvAzyGD/11HN06cU30JOP/0n0j5J9kYRLZRYpN9Nv41ajY7bNdu+l7T+oOo7JshN+cDbdf98Ttm5Yx3HaltopCzacRmIAvGN5kwiewUHad/+t6AObvU8a8corr9J3v3Ma/f4Pr9KE8ZNFn8f0EaUVp218z3tXpgMP+uBfvLfwGN5912/ovPOuot6Fi6mzs5s6OnRfzu3N3FZRHZ472cQ2qypNwVI5B9hZuNS7xeaYpcTVAG299Xq01Vbr0/TpPcOSCcjVyy+/SldfcxtdfdUd1CVywfukkgcp6RYlXEHzeO4eGOilb3z972mZZabLRffe+wB96cvH0YQJU2nsuEmydnCew1yL93zIi686hdf+pw/bn9ZZm9fK2//wXD3++DN08SU30H33PUGdnawDmQSwVJBWX5DbxWtLUiBZiqpyDn0lY3bbbRPac/cthq2Lh9ODl//8Cn3zyJPo6af/TF2jx1NHO6/LzKFGHB015W8AtC3yVkgMS4WjkUlqU9XM95Ae2PAQAZIZXDfQEm3G3iRElIDk6ojDUYf8bNRvEEBzBEcatdHggBLrqsuAZ3ibqhwZJ/U2XKYBzAGPuXisWxoibgPsIXWq0xTbwVtdigZ7R7f8MNbURQJgW/GYkM7QUpsByJb6JaHWno4MwF54zQvhylkhrD6DjKsRKDmZ6kFyvl8cBW0exFEMKYMMEwPW5IFoL1tVOLFmPFraK9Th4PawkwB7wYumMgcqrFnTXmG9gnyINn1sgZcb0Y0GUuNZwLVACmgdD64bwYD7gFwf5hwpmZgoEILTpRgU50pN4cTvlHRoTCxZZAiiG9hhifd0jmZEDY6giyy6H1EwnoTRNGEa6QfiSvZhS8GO+poA+UU2Fy+iASYdjGgDkM995PbIWjJSin8DQeEJDh+FUdzVjLCS7ACLF4sjR4nU8HuSn0cvuyqXutfLecRS12MOA45pDRHihucqpOqzaDEhOlVP8KcUhe2JCo7K9e17xxIVL7zyFt354LPiNZ5/AFKK+C4hevCJF+iq23+X5ZkmWm5GD511+EE0d34vffTrF9Kf35iXXMOD/S8HbkaH7LYRXX7rQ/T1064rEh78/pyouOyWh2j82C468T/2oTVWnCGTcsJPbqcfXnb3sMgVPPOusz8l3mzPv/wmvT53YdjsIwwIxavjwIvq53c+Rudd8+tqW4ezef73XmNzOFyiYmqMqEjAc6+UkwO8OzIhpzaubent0xwFT074f0NZ5gYrL37kQQR7ngPw8Z4Y8qeeQpFBZ6LCA1WlZjeM5bwqbGFSa8B3lZTQHavsrJli8y6MOYbexnzd0eiVw7ERCkgNI8qUXwVPzmSZV4gKOzwiHBfGkunipPBYipnrwz0RxPfyxshMtScq1PBIPTKaEQuBvQgjDjCnqaysYwE01ysK3dU2ZuRBaqz4tDuYKDia+DHTu9QwRJ5fX+AZFccdYBxSX9QOndn7xDix1mV9a/QvjlKaRVxOb/G51uphq6YSWeHB9DDfiVcz5s4Z12E2UpKmaQOGDoemeu/LockTP7b+3z6iQmWPiYGhF6EfqhToCe0SNNZdZzpYco6+HaIiiD4eCjBCa6aguKkaPO69rg0J4ZkoOiX8opHJREWMfJLc9UHk8F728uinLbbdmLbbaSsreLdEQJWQN3/YEhUv5KczcHLi906nV19+kyZNmCxepLnHU+6llcuMtGHEYvroPx9Myy43O7yAPZvOOfPHdOuNd9HUyTMa5EGir1oRFYkI6Frn/WjO2ivSXvvvRN1MVAwM0I/OvYCuufxGmj1jORo/bkIAgZv7jI2rRVJMmDSW9j14Z5ptJMXLL/+Zvn30cfT4I0/T9GmzaPKkqUJUcIqDUkQFzyjr2DlrrkB77PtBaQ/PL3vnIgXW25geuYXn+IxTz6XHH36WJvdoO8TzGykJpCvZOne64G0TFUv4sNRPm239Ptp2B/W+nL9gPh1/7En00INP0vSpswU8F9IkIypQIwX6ubzG8xGp6Y3yyEUdqLLw/g+sQzvstJkcDvF57NHH6atf+jZNmjidJoyfJKBcMZLAp3QIRBTrFH32ggXz6OP/tD+tPmcVefSLL75Ixxx1Ir35Wi9NmjRV1gyKW4aXG/nQ17eQ3v+BtWmX3beRtr304kt0zNEn0huvLbR7xwhAwoAFX7fDTh+Q61577XU66sjv0jNPvUDTpy1D48dNNHnOyXpt4/s2XI123m0LOaiz7F338xvpu8ecQjNmLEdTJk8PpBKI0Joez7000R8A5jU5FjsnpB7TNDVtbSNox102oQ02XDuZFzyDQSL2jGYZ0pQ06Yf78cLzL9KF519JTzz+B9EfPIfw5BPXgtT0gOaUNeH1Fts8vb0L6O8+vhvNWWPl8CIG3M8680L69a8epokTeX0x4K6EZHoqy20GHSnVBzoHa669PO27/3ZKnA4M0Lnn/oSuvOxWmYNxY1kfVSLKjCzDeglj3YLAKI0Vt2H+vLl08Ed2pE02fW8gFM764YV0910PU0/PNOruZP3BAKLq0aH2R/Rto03m0C67abSIkGjX3EDf+fbJIpuTWbePGW8EtwHZjgA0SEzkktu4+pxlabc9tqBp0zlyrWmL9fX1CmjR1cUgfvN39oa89ZY76acXXk/t7V3UJQAuA6Na8yEu4Sr0JcPH7eF9dZtt30sf3El1HBPD3znmRLr/N0/StCmzpV+SC79qR2CPLhEViwRY2mf/rWmLLTaQd7788sv0zf86nv70p9dpyuRZNHr0uOAY0Fh7KggyZuu+Z0U66OCdqKs77i1ax6aVLatSwvrEry/u99NPP0fHH3c2zX1rgEYzsCyRCLFAsY6PT1Tp7UK332TrD6CRvtmkqwA0AvRk+4nPOu3tI+nQQ3eiddddxXRplHDoCdzD7WSHiuZZcQk9+eQzdN6Pr6LHH3+eukdzJF2Ui/hEbZfmp9e+8Dv6+hbQN77xMVp2WXVWuOuue+hz/34kTZ22HE2YMEXID6zRWMhXwXGpyWi1k1h+P3PY/rTuuqvL9azb2RbAmDQUnelOJjjhbOWvYVDwjl/eSz884zJaIOTSaJlPjepQvct2BoOmcAqU9GnZuOv6G6Ddd9uY9tpz68SO1JqFQ8tSqe383Z///AoddfTJ9Mxzr9G4cZNlrBpEBTv5Afi2PutCdCnDbA8R73cGfyXCrflBii/2bOd+iQOR1RnA1bH/FjHj6n0p2Ir0dVzfcZFzRFIgVlWYOz8OMTxNu1gdNZm0VHLCalFaijJup0R6GMAq5wk+mzNegHeFhyLtGC84n48/OhMFR+Zwb0yvp0Wy9fm8D/VbMW+MUUJUWPFolSsQQHE/VFwhRoKDYOE0R2wHc4dY5zDe41M78n2Yp9KcttbWwWsKIiNDNCgyH6MjxMnZalJofxVMRu0NlnEA4r7v+tCwUwW7AvVPfH99ZIgQO0w28LuYaGOiy1JaaoRHLLCppKlGgjCpkNrwOlcAx4Wksxqd3H6eLwbz+/o5JZ1GMqhsLQnrOBBdgjm5tF6SHk1TBYc6qLbmeN6RZUPWkRXnDo69tpniXbwouI1q38VC40LUSPpDJTJAWkFfNubb2s39lD44jDHXW/7enLjAORrXoCauEI1ZajMsC24ry6oQZrb/cGQfF3FBJIV8nzmN+/Ura/f/F6ICBXtKeHM0shW4v+zWh+hrJ1+b1JhgGfrXA7egQ3bbkC69+bd0xOnXN2pQ8DWrLz+NTvnifvTmvF7626+dT6+96dIOOSnIiYpbf/0UHfHJnWmjtZeTSAqO2ujoaKP//N6VdMOvHl+qiArOhxY3kNRBJe8/b/rnXXsfffdHtxAX2/p/47N0RMXuRlQke594IcWCMZ6dF0jPBkoWKw4CLUzVVoq/RFZUMLcQ7iSKlll55LDEuwOIy7/EjQCeuY22+zZnHmQy1zhpvA27KfG6zw85blGBJS5bQfYtQpZdflBVjPZ7aJ+B5ZZnVphnzgsdvKVdYZ+wCKSjhYMYikTH2UDxZXl3KBqUmpXsFaxD5/NOagPZIGNvNzWkjUiSWm5GbsAqkgJvsmPrDA1z/O3qOJRuTrWXGK/mA/03Hmv3hEu4PSE41PgUTwCkquEQUPHs0LyMXpZiGzLv33DQKhukbKhmXEWix8ryg3GNLU8HMx2HVqn7S88v85P53Ok7FEbxpJR9b03AOvDGgX6nyzA1DOqOhTDx0vaqPvCfSIjBZ6igpSrEa+h38kA3b4i0MuBR5GIIEherCHySkicmOpEy0HGQ9aP5TMUQcx55Xm3Zym6shzghlh4BhYmXaD511S0gdOL64/f0D/TR5ttuTDvsrAfM+fPn0Rf/88t09VXXCnit3saR5HCd0H9Kt7yM86GhnUZ3jaGJE3toSs80AffziAq51cmCnO2Tfuuh7r0brUk776lpmHDo5TG777776fAvHkWzZixLEydMUg9YJ/BBvoZLVHB7RpDkol19rRVp7wN3DkTFWWeeS1dfdgMtM2sFmjShR96lz09lHsPB7Z7QM5b23G8HWm6F2XJQf+311+nE759Ct9x0O02fOoumTplBE8ZPDM8qHeYZzhnsH6BV11ye9tpvR/F84jSAJ55wEp3w/ZMVYEWan2HqVG4j75/d3aNpwrhJNG3qTJo4fpKAcnwYUnnE2sYUo5JsfMlfQlT09/fRB7Z6L22/o0bxzJ8/Xwic3z34tMwng+cc/l4mKgzGjUxqWFVFnZlpiaGv0XXKstbf1xeiFhAaz2thwYL5dNrJ59Cvf/UITZ06k8aMHmvh9OkkeLsq1Ycq2wt7FwiJsPue22uO4cFBuvD8n9GVl90sQO1YiYyIBImuc3XS4DHs6h5JH/3E/jRr9kzRHRdeeIncO43JHgZ429ot8mIvi7wg+sVtd9CXvvBfNGvm8kIKMdDNY53XqNB39NPBh+xIa6+zmrz6rbfeom8deSzdf9+jcr+QKZ1jQioHtf2WQhCxfxRVtdkYBpq2sZfjokU0ceJo2mPvLWmVVTnNkl7D4/zCCy/S9dfdKETKI488HvKvT5s2lbbaejPaaqvN6D3rrSPrDZ+5c+fSpRdfS7fd8huROU3TxKC/12nNHO7+EKtExXw69GO70Rprpp7ODB6fdMLZ9IfnXhUv+s4uBtmYlPR1mvLxAlGh2oSJiTXXWp72O9AivAYG6Kwzz6PLL7uZZs9cicaPZ92nEQf5x9uigSCB0s02e+lTcXGwrC6mhQvmU8+Ubvr4Jw6g6TM0BdQTTzxJxx5zGg0OdEg7Oju6tVBk0f60h5sdyOM2YeJo+tBHdgzROn/605/oi1/4Br304ps0c/qy4nHebWOmoo/5RkN1b2OQ9AObr0vb7bAxjR7D0Un66e1dSL+570G68spr6KYbb6PeXvUa5c+GG76XtttuS9p8iw/Q9OnT3LOX0G9/+widc9YlNPfNfgH8eQ/UtIgx9VQrPcJt4n2ViYodd4467qhvHUcP3P+09G3sWNVxBazdPZrrVSkYGSIqrBYA66Z99t+KttxyI7n+pZdeoq8ffgw9//ybNH3qMkaEdKSkmAfMTLbWXXdFOuhDO6lX7UA//eD7J9H3vneyROqApPEOJb7fnE5r3313p/3234tmz54V1uKjjz5B3zj8B9TZOV6juwTUj/ulRnb7J0VgX8+fTQpaV4XZv8GoaioO6FzW123tI+ijH92V1l6bCUSVHd5rbr/9Trr66uvohhtuMz0RbfeVVlqOttzyA7T99lvR6quvmujfN998i84882K6997HhYRps8iKXBZ834QMWbiAjjiCiQqNSrvzzrvpsE9/g2bx+p0wmTo6lOhW4NMBnuKJG+n5RYN9dBgTFesoUfH444/TlltxNMxYIYylypThIdIGq5fAY7L55pvQLjtvRxtvvD5Nm5bKO5MwJ5z4Y/rjH19XeR/VJWc7PqMwlsQ6UVNnsX3q6x9pz3UN9tFuu76f9t5rm2BHfv7zX6LLLr9Wo1B4DXG4E9Jtmqc/zhHyX3fOVfBZU+eNGTuJxo7poTHjJtEoidJJIyrEGxnREtxGiwxBDQzJYGBFc8X5jO08nOOyycM6E33DtUrMKQm1BqLEKR3LH6lFwCmjmBiTtQqvcS0eLLnqXVqvFDCNNQFqjhewjWUFmXMiY3eSXsoijVhOJJ21yZBMP1I8Q6awBN2ygazC9i6RdAqkplu7yqliFvy71DOxefD7DoBlZMtAMecQUWHzLu+PTLAS+vbciD1oakmA2xGz0PM5nF6b67E1VeHnA5gD/5fPAhwFguLq3ETGQzhqQObdSBqtgaRk3iiJQtLi4slzdRINBrGUXZkjC18vBIWlmhKSJ1sXErFgxZ8x1wzw9/dpenCte6DRFz4aJdG2RmxFWVmixd59tIbVV2CSROqPCmGi4L+uDbVhBHTnlJ++7pW9LEQOALS32il4r+r5ODfcb7Y5+R3IMCBkraS20tqNKMBdm1HYMR7TknM1Rz1j/2u96YY+IsohjJPdV4uM4DHkVIKsJ6OtEuda6vOYjkMaSnwHPRJl3p2p36mpnx544nk6+aJfKhuffTz4x/9+5Y359OzzryZpncaP6aLrTvyEDDbXpnjkmZcaz+EvmIA47Uv701orz6SvnnxtIzIDN4GomLPCdDr2vFtph/evTnNWnEb3/O739O/HX0G7bLYmffYjW9OLr8ylD33xXCE+hvr41E/fPucmuv7uxwMOWr13CdGCvgGav7BvWGTIUG347/ndluQwIyoaREUO2AP8d4SEnh3M47xEVPhDUEgDk3mw+8EAWImDpGg2vUD2SlekWMPY1AtBD8yRcdTrAYymOdc9CBBCATOCQ7plBI2ePd1RbOnO0830QG5T1Y7FQtBoW+JZ5l8NQ9siWwRMtE0/DKM7LKvyRZFdKyQmYcEAHd3DgwaPAw4QV72ksdEgYsBSLDVZEp2LQFSoleMBOolqGdlhxXcNEEWURyIDSeebyyaTr+K6ql1TOqAXdF5+CpfNB2B7SOdTWdGOUApsOC4N79e0SADweJybpFUch3SjdZtSRS4TwD4USIwhtyX25y8nKsyyDRs7JtX3Az2xdRousaJ49nPc7LWwlC4ZzEBdk8YDqo88CoNvOsW3ywqPlR45XKICOjITmuANkgBN5ba3IiqiXosp4LxBr+RCWSbSqCEvLHqQ11oYNlb2jCGJim02oh12iQfMr33lG3T7rXcKKM+AdqwBkZuHWEOurVK8caSAO6O7R0taEKQVyotex7MJ7o/9Zt3CXqkHH7oHrb3uGjLI9977a1pl1ZVp4oSJ9OZbb9IJx59Kj/3uWfHslhRKVgBPxrdQN2Aolc/DxcDgHCYqDgB4M0Bn/vAcuuqy62nZWStSz0T26oPXpbem1Ohm/dA9ehTtsf8OtOrqK4reZkD0B987iX5+zU00dcp0mj51pnjia5RJsy6I3z+4PatlRMUpJ59GPzrrAiGBRnPaFfNkrq+i+IscAka2Sa2N7s5uiV6QGiIdHdTGRTjtYyVb9S+YICEljddzuKP1YTBcxSCeEBXr0fY7apoIBo+OPuq79LsHn6LZM5enceLlXyMqsI1HmdFnDzW7w71GiU4+QMxZc3lJzTRm9Gh68623BBjaYIMN5E2/+MUv6dijT6VZM5ejCeN7ZDyb8h3HJAIA+h2IkFHdI+jj/3ggzZ6tINajjz5GX/7C0dQzcbqkDeoc1S0FRr3GQ+TPvLlv0n4f+iBtsukGsubv/80DEukxc8byAoxzhMwKK82g/Q/ekcaPHyde3ccfdyLdfOOdNHvWChKNJFEbUnw01SXc/+VXnE77HbSD3Iv190+f+CwtM3slmjFjWSG6JMWUW2ut0s2kAE1racV46aFQvXInThpD+x+0Pc2WFCraXgZoTzv1TLr4Z1cIyMakkaSdsTonAqItGhCZW3GlZeiQQw+k9ddfL6w7lkP+NzcAACAASURBVL2LfnIl3XbLr2XMNO2Yj1AoExUiTQYALVg4j/7uY7vTmms1U7I8+eTT9P3jzqTe3iUK5kuaOj40N/dSLLaoVTT6iImKfQ/YwcBk1kfn0mWX3kzLzl6Zxo9nfdRR1He6djOEyf729rNeFj00YSdH+2gxDfT109x5b9L2O25Eu++xncgWA0M/u+gKuuRnN9CUnpmi6xW8Vduy9tHURQO08+6b0uZbrC/7Bc/PaaeeRef/+BKR36lTZhlRB1LYr1+zCuQ5XENlfdpmu40CqMxniZtuupVO+P6p9Kc/vSygu+o4TT+owKWm0mGycJ99d6KDDt6Heno4LZCOxW9/+zCddcbPaN68QRozerzofERWtIrkAqjIhZO33nY92mmXqOO+deR36YHfPEUzWcd5oqJwvgrazTsBBVBvMbF3/T77bUVbbhWJisO/drQSFdOXo7GjOWJDz1NBCzmARqL1+gc0osIRFSedeBr98IeaQo7TbiFKJsiIm1TZowf6afqMyfSpwz5G6623jq2JRXTN1TfRmT+8JKQnQ/outEdtHP+w+G+NaAqGo/VB7Rv9uIgKGN3uUeKA0T9Au+2+CX3wg+8PnsEPPfQ7OuKIY+jRR58WXdHVBUeMWLuE92+Wn/7+Xlp11eXp4x//kJBarBN+//s/0Ne+dhzNm7eExo1jnV9IQxQGXGeQgcOFC+cZUaFkzi9/eRcddtjhNHPmyjRh4lRLu2ROAjbH6rCi0TQyzv0DNLiojz5z2AG07rpc14iJiido5533pYmTpkl7mGyWFERGVmi9AsWApJ7PQL/066CDdqcPf3g/mmzyzr8/8cTTdNTRp9Ebb/TT6DHjxbFE8SP1VgeIqmOPYtbKKMl+NNBHu+66Me2z97Yy3vPmz6MvffHrdMONd9K48T2y9rQ4udUasNRMIBFweFKHRSXj+V1sR/I8dXaxLGqdEE5p5OVRSSltI4o5B6/yRpSx2shMKpQ+DMAiPZGMm6WJGiHNUY3owX1+FtsqnNJGam5yhIMMij6f+yH9CewbiAl9OyIxFaDk1EJGhkp+QR177hM+ILQUrOfoEAWmAeRyvxVgNW98VxdA8AhHWsj5FMMgm46eR/zZWGUHfbECxRaVAtwFgLhGU3BBdK3p4AFnPNcTQQnw7HAlgM3SVhtsiS6QtRnrFUiEtnPCLaV+amVz+LYIGWNWBf8XZAE/X8BkiRjpENAcfUEUfADCbZIUvDfnT+8YgLYSib0tUS9SJNydp+V6XWWyfj3VnGU88bVG+xf2Uoc4LGgBaI6QkLXkimSHubW0StzGkMnECm2zHevn3Hv/A89ASjrRCRZNobJkqadsDSESKRS0x/VIB+iOT0LQcORMf3+S1p1lS+Qf2ArsLpfCMtkrTWbk3UKm6I0hEiOCNPK9lwGssVYy08R0ko3HnIP6hZjXMWE50BZi/PFvr0e4WdAFondF1RhW904lKm677yn63HHDq1GRGww8wAfssB59/pBt6e6Hfk9fOfmaYqFsrK1dN1+LPv2hLen3L75OB/zHOdTbzyFz6RYAomKNlWbQK6/Pk/oWN9z9OB111k302lvzaUx3Jx3+iR1py/VXpoeeeIE+/d3L6PW3FrQkE0BU8Ju+ctLVdOUvHi5uPPmXQ5Bpw3rGf+9Fb4+o4DbmR4WwyCzMSjY7B9hig5LvHamQAPyBXVeQvHogcS/HAhUFwJsv8ia6vIvqadE83EQdLq76gNkTQ8XPB0A60UdWsMZ/F5RRZRL9ppFckhX2LFs50TtCGd0UwAv34ATYiqjwF4fH5OOD1DTJYNud/F16veci4P2IMY+5R9N7tDCxSpPej+cGCbFf9SrdWl3of7gHsmLkSlZ0vARz+blIYZQ4+qXjsGezPW+DPYrnBgafGCiGnYf14TZQPKvxHmdc8G/szQJveM23GIEMz6BGfqseUVHy1JaR1yWgRaksOgGeB2WiolQgNUa81PRYiufbS5NZxlx7EdMRKnMBZdBiONwTG0JskOshJxrfMi+Svs30hs/hGmQ27WENOpE9IZlPMyyCtgGoFFbCMIHRuCYaqk0EM6Z1a85FRXekyi7+xeOUNjPzkrb5ceQxjy2TAZtnRMU3jziKfn33AzRjGntmc2FOzaWNUTHF796Nf6pu4Lnh+eJ1wGCJeCmzLgxFMut1cFBIk2V8+ZVn0b4H70ITJowXkPXoo46h/fbfh9Zaay0x+tiD+tQTz6WZ0zWFDXszYb3CwwdeXx58q3l9K/AyQHPWXqlBVFx52fW0nBEVmh4i5oSF3pN1OZJovw/vSqvNWUn2M825fhZd/JPLacqU6TRtygyaOL5Hio7yuHqSPTeQAUgzUbEnp34Sr9cBOuP0M+mSi64Sz1yOJmFQNjns+MNNIBkcaG5kEs8LH/wl5ZNEzfhom5J28CuotJqGJiu4j62JihVoHKfXYsAzqx1U34Jbvbe86mt2oO4R6hG99/7b0fobri3jcs+9v6abb7qF/u3f/lnS1Lz66qt07DEn0fN/5FQr0xXwd0RZTbfie8zt/PlvSbHubbb7gIALLOennnK2RmtMmWXRGgxipbpc034spNXmzKYDP7Q7jR07RiIefvD90+nR3/2epkyeISDPbntuQZtu/j559pNPPU0f//t/oQnjptJMI1gQibQkKXTPHrL9tNOum9Cmm71X3r1woZIc1//8dlp29ko0ecoMRw66tlXI4Gi7tR6ZsHdr3g4lXxczcEB04N98kFafs0Jw2rjv17+hI444ml5+6TUhi5gI0DROXdRudQ34CQzmsMwtXDif5s57g/bdb2fae9/drDYICZF49pk/kfoBEyxNndasyPWUggfYChVQW0KtiAr+/d577qNjjj6dpk6ZaeB7l6T/UosIShtyCkBWjcQaUcERFcvMWlnaW4uoaHXgjpCv28ud56wv9slXaOTIQurtm0v//G8H05prqlc3p2b5/vFn0B9+/6qkuGJSWvNh1z7qvbnanGVovwO2p3HjuY4E0d13/Yo+99mv0Lixk2nGdE6Jo3UWvCe+f6ISUIO04UZzaOfdNpdi2fxhfXvyyafTj390EY0XmeiRMWcCigsHjxyhRbLl/kFeQwto/sK5tOyyU+kf/vHDtMYaqwcHk1/fez8d/a3TFGwfM15SZOg6rFoS0gboj623KRMVM2YoUcGeqrzuvDcq5FUBagMqANEHksmIin23bBAVLzz/Fk2bvqyQK0JUmFd9cza0EO6662nqJ+wtp576Q0mJNm3aMjSOiUjeWwC0uHyUiNRkkI7JnokTu+iz//5xWmUVrdPy6quv0XeOOYWee9aiiUwueOyUBE+9tGXfz8533sBIADvdcKuzoNE6Y+iT/7QXzZypBayfffY5+uQnP00vvfSGyCn3rbOTo0a0Pg3GGuAvE00sGwsWvEV77709HXDAHnTBBZfSJZfcSJMnz5T7JU3SyCzizdoGJcHpeVjvaOonJaMjUbESTZw03dIZNW31uIYUUOP2fPbTB9J73qNExRNPPEF77XUITZu+PE2YOE0iVxjs40/Qo1LPUVPlMGE70N9HvX0LaMUVptNnP/NxWm21VYK8/+qe39CRR55KozrZeUFrwwA8w1xIUWSJquCaijqTvBp4vHbZZaOEqPjaV79Fv7j9AeqRVGTjxSpHZLqkrszqYUp/LbMAg3UMcPL88L+ZpGB7Ses7xtR8opsSAq6ieQKMYiRn7ciMCAUQCzijW3vkvGg19dTBksmJNukbCkxL+hq2gdt0jAC4Kyit611TaOm5hteQHkHUyUf6JATJCLGdpUCvq8WJGgWaYkrvUbxDxyLq/VRPSSq0jnaLjFGP+EWDmmJM79H9DH8LEG0OlPjOp+tu6BRx9BkUwJzlVexhS53lr03O5xVDLMGfQNC6hyD6XM6/TPJI7Q+sIZ1sv/95kF77yREomqqH50hMX0fUSKopJhQsmsiDzCCFwppgIgPkhgO/WS6YvNGIGy0IjpoN0j7UoHFkEBMYXOCa2yXFyaU2ijpehf3A21iFVGxqOeiZViOjmJDgOdFsEFgvclrzJIllNInzo/Lq+w4SBqmYgEUgNZK8NtGBTS3Ozw+F7U329OxktUgcOcV3y5i1tcmYgIj01ydEauh8Kp1YXyAnhKAxYpN1UulTs5/8+kB/Zd3YWCXkjgsW9O/I57J59lO7VZ7/TiUqbr3vKfrsdy8fdr0HP4BdnR30g8/vTRuutRwNDupiLhXbxj2cA7KDF+LixfTp71xGt/3mqcb1ICrWXGmmCP1vHvujECmvuLoXY7tH0RlfPZBWWXYqnXn53RoRIuxlUYYkmoNrVPDzvnryNXTFbcMjKspP+9/8bdhhjZW3ELJKMe09ps63zjjYn9k65IizOgJ8mGBjgeeWjRt4bmBTFabRlF0CEmcFjIYiKuJBTIkDgNhSINp7wNYOuOiNKQH9s3JQwBlSQDG3UWWpZpSdLQtWlagoFVzOFL0Ol3mSy+6SkS852o52WWhcBc513c2viNZ6dCzyRagBHiuA6D3BPOmAA3c+tmoPOoBLBcItFjw3ftuKqPDPBykmx/JWc5ERAi1mP7Qr2XzZcJACXDGtmW+HyqRKqYKp1p6EZMr0Q6FNnEqOw6TVSwS5SSMhEp8Q4V4MbXwc5gtXZ/Nt+ykKVbMB7wsUN4ip8v5bHW/Ib9rW1uBklI+87X7M4jNqR/yaBtY0ARpiLLrJDLN4gAJRwb23ou0Vb6kh8IWmasnQnBRUGn5PjJNIu2hfljz/ZR6SiIrau+L3eV0Ok2h5pxhpmQevACJFomI+HfXNb9OD9z1Cs2YsoznQGfDgPcTrEOgCr0Zd3R/xehuhKad0PaKtBtDVVLi1kwG6nfbcijbdYgPZux5+5FH62w9/lD7xjx+jjxzyITlAPP/CC/TtI4+nua/3Sp0FKexrHnvQdohUS/R6Za8ZLlGh3rXx4IBICrZ39z5oR5qz5qpidHMtjXPP+TGdfcZ54r0+dfJ0mjihR+tBdOie2+rDz2XDfPU1l9caFUZUhAiPZVYU0oPTP+WfoFPdAT25BunBjFjyJAVkprFDlurVJA+tw5O4rBVR8TBHVMxagcZK3v1mRMVfk6iojTvjx2ybTJsxkQ788C40efIkmccTTziVbr7pNvreD75DKyy/nKydyy69mi4493Ih9BR4TAmj6tya7PN7uNbErGUn04cP3YsmTZwot9x22x103DGnSXolLhav0RourZIV7WNwaO7cN+iT/3owrbHmakreXX8znXrieTRt2mxaZplZ9Hcf35tmzJgm7b3op5fQST84S8Z42lQmQdgDvl09Ph1RoQetQSmivexy6gX88MOP0D/+w2E0acJ0aRdHUwhh52S4lRd9A2isTkDUEwoKKWmy+15b0oYbr6NAzpIlkj7lM5/+AnWOGiPFxydOmCIe/ZJizgA2rHkFTRYJ+cSg4VtvvS6e7nvvu2sgK57iyIfjz6TehSNo/PiJFvmQFwKOtp3sOo2ICk2R9dxzzwkIPWuW1tVhkuSin14hBbAn90zXcRfPYNugE30EokJXoRIVKzQiKoSomL2yFE6uEhUtlIsHwYMnrV0fDvXeNrMUSwsWzBVy7JBD96Fx48bJ/Nxxx1107DFnKLg9ltPZjao6MPFc8HhoBIqm5HnttdfoG4cfRQ/c/5iQFFKbIoxRqRMqTcssO4UOOHgH6unRdcOE07Hf+T5deeX11DNpqhAM3J6u7tEWYWPkk3k485pgL/Pevl6aP/9NKTr/z/9yCM1ZYzWZW5m3n1xBV175C5rEaagkwqCcZiu2UmWWZW3rbd7biKh48P4nCUSFRpCbHFnUNIsCgCSdo+j0I38bQS4RFX8BUcGrjNMIokYF9pbTTz+bLr7oOolqEaKiszPOZUG983wy+D1v3pu02Zbr0kcO2UdqgPBeesnFV9E5Z1+mhCungGobpR7QGbisZyZ3DsgUvdiAOfVlRx8Amn78OUXcZpuvS3vtpbV1GOg6/fSz6OSTf0RTpsymnh6tfSLRYEJcof6JtkHIikWLxImjT8iKuUIS8Pfd3eNkXFgWtDaMSz1tTlzwohdSRurlgKjIIypWkjpHoyo1jrwmQK2LzxzmiYonad/9PkqzZq9MkybNoFFcD8SiaMSGROYCA1KFsJB+9QkBM7lnNH3xC5+kVVfV2jpsa/z4xxfTT35yA42bMIW6uzitX1r/hu2pkSOs1o47t3HBcCYq9gqpn+bT4YcfTXfe/Qj1TJ5tKaV4vEdaYVn1eE70UPA61nlgW591idTJWMKAvNqRtizClCfSUbJ3Ct95B81gK5nRGGpFOuEKhIN5wMOb//+w9x5gWhVZt/AmdtM0NJ0jDWJWRB3FLKIoKogCKsmccx7HNKMoiqKYxhyQoDPmnEfMOWcUFcWEiAlo6NzwP2uHqjrnPae78c7Mvd/3+947n80bzqlTYdeutfZem+WGGHgVyR7rcxRwx7/tnAIpnhXNEjUuZIAnx6zvOXBEZXtk/AT4B+ANoNZqBeCaXMxYt8rwDB09SkedbIw/A/O6lnhfRJsgQccZZvIMUjfBsmVAwKgEVocOLCkk904g1kB8AFw131Ij6/EMluVjRZYN2Oa+Tzz/m8ye7IMRMkolrsJgQ868jF3H4wo+C0bWuhAV8jnqIojEk/U9g/q8N8gYivSeSlvpXs0+kv4dxy/CYCkrCM19xgXHhbyxotYMksOP0NoR8hyiZMHnLs2+ABHD9SUsQVI2itDsZWyUVo80PGdIMfeMhDXBLZT0MZIJF3Rr1ApFK3lmNUbQIMuo4TFi3zHEoKLNktjC4OykAQOu1olmSlgfSmaJl06DP4T+s3kkGIiSexjTCMrl782WQwkSk+nif2tx+1ZcpeSPeN56WE3WtAZT67wSc6I7V3j81fd5jVu2lU+g4PvZPsTn5z+IiugYYAL3qyykOy86gAcVWRJNzVL8p7VXUa9cyu/RjR5+8WM694YnM+o/hBkVr74/n8665jHOpAjtCu4xcL1quub0PXn8cZ0nXv00Ub4KbfmDqECRmWZa2dJMK1qwCTZQS1M9jQyKabtgLY2Gx8bPix6Fbjp1dmlscG5guI3tdfUGbNB9GLhscbpAEw+mwVzJ/FwXbVBwJ50YiM9NYZblCsnZFz7fIky1VNY4NoedMxKb2KHuYfSjZNQ33n5PVIgRi/RBzFgZi+/A8UDHXu6t4G8KwsrPq9cMwW63rnQf80ChOgX6Zf6PRqX7c0AIfrJbGFWF+J1EhWVwhOcNa7Ol4cbni+vbGDHQHojYRwWoHA6n4skGzZ+FByMD64xkwpfUC3T3SjCCYTs43VZrWFiWg6W2hgRCsJTiM8/9O3qrALjRb5h2Io6wvI7VyckkKtoGDmOrLPin3TcclWjPi1Ng99C5mjg4/s32jF2kTTxUmlLqHByfueSirvnCWKNpjq/HyuPzLHJQ0ZtHyDtbY5HFtmpPEqsL7KQ/0uzfqhIVIAWimUw+gyGJqMBjsvxMRkbFcrr4wqn00XtzpV6AgcZMugbziR8/GtkmtsRGTzIOPOgVGr+0jAo5iMKR7JGXQ/sdOopBVuxLM2feRjdfP4MGDtyUzjz7VCorK+X377zjHnrk/tk++wMAtzVCo98iJGUrzkzbREVflofJ1owKlz/G6b0radc9tqeNN+3vSIrb/3EX3XTDdCouKHW1IFiiqnMXT6iIB+3XfjD5jahARkVIVHDNjIefpj5Vq6sUlScqwkNT2t+R9RVdvrrrWNRrzEQlEBV+/mYW2UzyGf/fISpS1q8eUAfvtCltN2Rztq+Ixj3pxNNp8S81dPKpx9LwEUP5oD7/629o8nmXE7V0ZWCUCzK3QT4F2zofRnDwQpT/AYeOoj9tMoA/BgE3ZfLfadmSZilUDJ1+AEa85CzyWKI5UZAbdS72GDWUQZ35X39NF5x7OTU1dqRdhm1Po/Yc6jJAzp14Ec37/DuqLO/L9SUkYl1lPIJoRKyrjTdZk4bv7oG+GTNupdtm3sPgOJMcAG0VaBVL0Lo9XHWiAnu1yGmwBNeeO1B3rT8wd+5ndPppZ9Pi35ZznQ3I1ICkQHaIScxE7arMTdZZh9xP3XJavOQX2nvsLjRstx3dvv3E40/TbbOQ+VROuTk9JAI/IiEnz2jEOUBjAAx19cvooEMBvAtRAYmwW6bNoDPPOo169szj9wCiz5pxF7395qeUn1/Ckl5MVgTRfGJhvTxna0TFw6hRwUQFauYkE2St7v4mdRGALe6gHdDKYfQlkwxNDbR06a80ZtxQ2n6Hrbjv6urq6JZp/6RXX/mQiZi4ZJDZAR6D5ibaapsNaNfhUqAe55E7br+HrrryZi4OXlLsC7zL3Mx8CjmrNNG+Bw6jDQZAbktIhVtuuZWm3QQwupyKCss5mwLkNQAfA7XMmTVCgAE6ZCc11DF4W1LSk44/6SAqL5fCxz/+uIiuvPxm+mHBEqkzkoVC3GlZFdLWVSEqjIbg+kuWXSEX8QElwZpH+/H8adJPSRkVSXYYyxUyGxts2DeSUTFt2iy6/96nqLxiNZG0YzBf13bChGJApaWFo/SXLPmFJk46ltZYU7IqPpnzKR1/3NlUXtaX8vIKKBtFo62+nltHtqbCgKVMWxKnKpw3kVFbBSRRE43ec1saMmQz7tMlSxbTOedcSG+++QmVlqItRSwnhMCiaBCFm6kKlAPUlywE2Gn0O0BMzAHOQowVCbe5ZQAo+1gs/bQ8RfppVYgKjPlyOgUZFSr9hBoxY8ceTuWVa1BhQTnXlgilJN1ZlGWEJHMc9oXJpaZ6ql22lNZep5JOPulgKi4u4of/7vsFdMH5V9HCH2uFqOJi8oEkJAcwekDe9qPGxjqWfhqt0k+Q1Js0aSq98cZnlF9YQdndcnktsn/HEkd+Lwv/FjJONO9RNBl1GGAjAXb7eejtMC8VHTa3x4TERJIRDKZXxsdqF0PfyQGrVpRa224EG/6J4suiny8t4oyTFS0MSEvtr46cSca1NPi/ngCCHeToeSa+sedJ0Jtl7XIwKVIK7Tl1L+vUyWpvWDCX+M/+FTuvOTkq/32WjVLCqKmxmfdI7CecBbBCpKxgH0HUWPAN7GkcnLdx6Ni5I9fawphx5oGTjfL3xGdoGZ8fWbc/00KZyTH5o9C/wDhb/YPwt9ameNuM8NVJ54gKIxmxxjm7uVNHJifQ/yyjpLJDaKusKy1KzgoKkiljz2iEBPrIF8H25IbjvDQDxvwRHjHLJFClBPR/fUMDZWdnU329l8EXUic4LoT9ltCHlrVkGR2cndPUKPJkmjkUziled4HUGMYZ3zcCziSwTLbK1iOTLIrNoWh2mF2RMbIYWJVFYvvIxKmQcazkooSJ+aUYD7ykLiQygFp4PRkGaWvKzuviPSX4DDpeYduEDFDJ+8RNMv1NI9hsXoZERXh7vke4LEPbFF4+VpfJiArO7P2DqIgORFaXznTBMcNo6Jbr0DuffkvHX3w/La+X4iZJL5uoQwauSZOPHU7L6hpo5Mm30JJldRHjEy+m/cBzHyUSEDDOIwf3pzMO2pFqahvo6AvvoU/n/5hoyP4gKtogKmLgWsSIdyA1VhZtjk0QAJEWCtbBzgDRkupT6I7DIFkEcPGbpHc+9FD8O4yDpaC5zUZYAP+KZXrwxqlRSo4QCCLE0g7O6cRJ60SFZmW7PnARAAboRWKKZT0x3RJG8f8uosL6Pe6UiCfgwX7nzVkXSveZFQ3aGVnrESzSbbc2QwIyRd5Ky6gwosIMvLtHcP1oxHqCu6XzKyVRILLphOPIuv0OcNDU1hXibITjYAQGj104vVojKYKDvjH2looYl+sIL+NNagBSJkQ6uMHCYGpEBheX0pRQHJiEqMg83HXImE/BsCVb9MgXrD8SRkLH+r9BVHC8ukYeCnDBUQYWlReplJ4STmEPEBCHkfmhWWY2F+zrcQLj92ZU8LqIT1pt97+bqIhChtJf/ydERZ7WC5C+EWrKL47WiAohBYWokNT0tl+4Aw6ozbTFthvSzsO3YzALwO1Zp59DP3z3ExfmPvbEw2jb7bZi2wZN/7PPnEwFecWq6a9a4oHPwn1sad38IMmNaZuoWI0zIqSAtRYqXyFg84i9IRM0gN/HPopi5BdOmsp1JFCTIj9fIhSlWK8ccBwRbc0xAlnbaO1JIioef/gZ6lMFoAMR1UJUJB4etR/SfLhwTKKHQVQGiPl9MaIiPnfTyP/wHu0jKrRGRUYWY9qu3RokmzzWaesOIAJ1aKGDj9qLqqsrNBPhAbr6ihupsLCUNtt8EzrymP0pP78XZ1rMnH47vfD0mwLed4fcimQo6MbS6pRny6ZFtQf8aQ3ac2+RYMH8v/32e+jRB5/jotoMwoMUULtnF/V1LsjVubA2PfnYC/TXc06mjf/Un7/+wgsv0Zmno4BrHyor6a3yWh7gtowKjCFA3wn7+yLaCxYsoDNOn0i//LSMKstXk3WmJEdGIEbKULSqnBmPWNIH5LY0NNABh+5Ga68j4CekfS6/7Cr61xMvUFlZFZUUVXJNE5Z9U7mm9E6XKF1kaIDgqa1fSiecfCCtv75IqSCy/8rLb6Lvvv2V8nuhkDNqyISgtI/GlPEVoqK2fhkdHBAVkGQZvusoOvUvp9ABB05w63PRop/o+mtn0Xff/CZZGyC2rEizzhnZ66yOUxsZFRX9GADG+k+az20RFfIMMoLsK1tEoAsGitsULQJft5y6de9Ixx63LxdyxwsZKVMvuZ6amzpzlgcyWwRscJAyAxF5vbrRAQfvTqWlAox+8cUXdNpfzqFlNU1Ugdoqrt/lTJJ59JQ2bLTJGjRij+2c5NNryLA55a+Uk92L5wUybECYsGZ/UMjZTJrGqighAF+wmcH/ZcuX0JZbrU/77DdKMwNW0uzZz9H1196uRerzHBmWOc9+H1GB60jUaEcXlSnPrvut8zFZYMYTFSkZFaWB9JPgM9YqhwAAIABJREFUppkzAZcEONp/QB+asM8wLyvIRMVsKq/o2y6igvsAe2BLI9Uur+EaMjvutA2/vejHRTT5gito4Q81VAACKytXiprqDA9BImtiCPJH9o0Y/JRGVOD3yDQbM3YHGrz9QL7EwoU/0plnTqKvv/6VybDcXADwYZ2pNIshGuwAaTE+0l7UgdB6Eirf5n+dWQic7XsiUXEelZf3o/z8UiYt4xJL0kdyDpFAZRAVtXTKyWMjRMUYEBUVqzNR0TUL9soD2mGwlkwDXzePMzSQLVK3lMaN2YlGj96F9y7sPbfeehfdcddT3DZkkETqlLBKTvQcL1lS9TRiRCZR8dobc6moqIqyuqF2ULb4hCYJpOcvNkMaWSw69yiOLTI5ADDR5xxNbq94xk2s3klIWIQeQ9y/iZCgkQBphya6W3J0enD8lUx8u4LUVnMyQdx+OUCCbDFpNzy7yP8AfLU+BCmBiH0BaWHb4POGNkHGTggmPINbQ5D1Cfw+jLeRJ0mQnUhOqZxMkFELoJjnzUoQvo1MVGA+AiQHKGwZFA7wVvmojFWDIH8NgLJsEoybgfnJBELSyVWujO+zmosqgui77hmtz/B+mJ1jv43YD7OlGpRoGRUsveWKnWOdrRRJqC4gt+UswvMzDGLUtoUZHSY/5QBrHxWpGVuaNaHXMWkn/M4KK3OBcf03CC6Mg8l+8TOpuo07vqQQFZhZPA6c3SLnL/SVBFBKTZOQvJFzmtgGk6riehxaJNwRMoGsldXWsDG1/uGTeVCvwsYAplKgpg7UpHJUmBfWh0z06DiaXBj6XurveT/EBVPr/GXiQm0ez5c2iAqbw5bh0hqpknZGYBsVwxslc193JcMdtd1tERWRtWpAoqvn8QdRkWFn1ulbQrMm7cPZCn++7EF6+s3PW5V9sguUFOTSP87fl0oLe9I1d71I0x54PZJVEScq7n/2w8TrYpy7du5MZxw8hPYYvAF9PO8HOurCe6hmeUNGW/8gKpKJCkg/JR2UmalUxl+MqcFOUrAIn9ki5g1RwR3vHISx0ykkgQNaZME6xlUdEqclx0WYoxECaa6iM3Sh9NNKS9WNhkZYRHFYvCZshzN4MPBpaHdqQ9oiKpR8sEOFmNfgyOfPbM64Bxr1PCaJAFoEMQ9apxFXHSQSy2vIx88lUaAmI/IxImyfBHbLBpPMVQZgm7YsjajwDTdjLv3D/9cA5FjNktCxCVuW3E9+MzOHzQVWa3qiyQYhSgfPAyeS54dqtkeckSTwMD43gvGyNSMOgUQsROdenJCIjYvf43zEprbO/iPRl6obqnUx4MjLK3PsVp2M89fxm65c3ai1eBf85zMqhKiQMfVaqjZWvnHtQMITiAoml8x5D/oQ71s0kMcdDYD0874tu+WGJm1tp1xgVTMqfC0ZPxV80cNM6Sfctq2MisryapdRITPDH80iYH+KJJBkwBpJ4bMoLOos89FlLwJQesjRY2mNtVbjr7zw/It01unnUllJFYMnm24+gPY5cC/qkZvLmv433TCD3n7tQ9aA756DjIUALLZ9KIye+R1ExWMPzqaqir5cYBwHbgYQANA0N9HwUdvTJpsNkIMqSIpHnqALJl1MRfnFDGAX5BdxBLoUu7NswHC++hOwFJO0NSfXX2vdzIyKJx5+hqrbQVRYH1vhvbT1GwecjWSKfp8hTc1K8/uhtVdSzVt//b9CVKTZyxVNTbTRwLVp2O6DKTsri+s+TLnocnrnzY+ptLiC5Z2OPH5f2kSzH959932a+NepVKkFrLtmZXlZhHaYJJZfa2yk+sZldMyJ+1G/fn24A4WAu5ilQfLyILMkIFR01ojOPupc7LHn9rTd4C15fqFNd9/5EJ16+nEsJ4U18vcrr6NnZr/Csk+oXxGvqSFEhQAlXER73E5cRBvj9dhjT9CFF1xBVRX9eA2yNFdYFyU+lROmwKoTFRK9uM66vfnZcnJyuC3PPvs8nXbqOVReVk3lpdXUq5fWMuB9sB0drsVVOZOlZgkN2Hh1GjdhBOXm5vKeDTmv2//xCEf298iFPEyYrRAjKlSWYHndMjrksD1cRgXA97323I/Kyypp0gVncfFu20/ffvs9uvLSW6h793whWBAFzb6w2EdZQ34d+RoVofTbrfTQg89QJYgKJgWSiYrWVqIB2CGY6fwf7Un+d+wiAgQ38pzbapv+XIga9wcAwlJotz8udphJu4AI09+NGj2INt9yQwYokImBuiePPfqMFtCG/Y73ebQBQt42ajaFZLAsWbKEzp80hd5840MqLenN2RQolszycQEhjIfhoJWI5KqehTTbXDIDfqUTTt6XNtp4A77+Dwt+oCkXXs2FhvN7lWhh7STZvvYQFfOc9BPXqFBgh4kKB6IJaeTPCRp9zFkXUlwZknGjQVRsFy2m/cMPNRQhKtKCDAn7bCP136CaJuw73BEVt0ybRffdN5sqyiWjonM75OwAQgnhupx2HLopjdhjB844QBbRJRdfRR99MJ+KiytVzktB2IzJ6eVAYinc1Jb0k/gmumeibxobaNy4HWi7wUJUoJ7QxIlT6LPPFlJJCYgKSAt2lVoH7hXP2QgbaNIxsk979yEI3Ahsj7suEwwtXMPmfK5REUo/tZ+oQEsQ5Z1KVJSvToWctZATkaIKgTbMpRBUhG1FZgMyK8rLetApJx/I2at4zZnzKR1xxJlUzH2FWhwi2SQvPi3xX0Z8WIYGMipC6SdkVLz62qdUVNybuufmqU6+SObg3GLkg/lEXI+OwdoVLsJagERdVzYkdv7X9lhARQQID2og2s8iREVAkvCzCPIogLT+HWYoWxFl4CT4DjIoMHt8TYgOUv+hGfUK5P8hQl89Ji2cHNY8QLCoFIM2vX3LjBfSADV4hBwzvMYAZpPmCaWfeGQUvPVS7dH9UIgQyBmF4K+A8bgn6jrxWUilqNHvXKR8hS+6zOdczhbJ9PUwStxPSjRZLQcel0jtDBkROzMnZ2PKc0tNFDv7CZDPNZBA3IROqnS03CdmW8KznN/vhPixQD9Z01pMXGVdbX4L0A+ZdA0QDOa+3cqINastwnJIQdFqfA57yxiYFo52Ul5mULR4usgzaR+r/bZ2229kzcgZxM9vH6jHgD18Cb622C15HrOT0RpBogjRketjIGMC7eRsIMt0UHJRbJHIWBkB5+Zds/SRzUXXLuP9TNZQMzeEeJGzPc9NzB0lVIx8aG6CtJo8gsc6/NzBbziYROesSQvGpkBE68ruyySJypNlfL+VN5h0iY2LzHGxJLaPm400wlmMpva/YV8Rskn/oYNkpNIfGRXBYMAYHLLH5nT0mG1o/oJfadzps6gRRX4ygzEyhrBzp4501N5b02GjtuS6E+PPvJV+/KXGfa+9RIVMcKLiXrl05V9G0ZrVxfTIC3Noyoynqa5BUoDs9QdRkU5UiMkNNimtycBFUdXQmDmH0W9obuTvw3ljR14LQwkj6xFUvzglDcu9AkY2vG+UqBBpHL4/6lOE0W8Jm0t8khlIycYWjpIDt/WbrsiVMMjOusUu5J4hVb+/NZMVApRRp1XWiZIGBulpZH58PEIj5zbOIJ0x2oIYKWRW21hmJirwHXGKxDiGVwgAcj0Usd13XwoHMn7Q1wLREaNqF4/+LpgmrRfTdtHE0kZx9CRSxPQLGTJhVt47qCYCwCMQaab/h81d3jgDyQaeM0F6JUesgKjQKB3WO2SAULVyw7C7NPgjaAR+B+faojpMQ1TsWWv9K32QeaDQ8QuGnvfBDojIsaK30FeUKDxzsqLzRg9XCdhNtE0pcyUG5qbtA+lERfJztwdKirSIo3S8RqWvURGuRWW7Wlu6sggjToT1fZyoiNqtEPjX1ofgR1v35JtqJFvGd9N7Q5JhxEMTe5a0EQdOaPxzvnQAJifVqCCAPg207Q6b09DhABc6E1L2TfopQlTwYwQH84j9Tx5r2UkE3JMuk+/Jus44TrDdwIEcxaxH7r0zS70AZL3yimvoudkvccRtz9xeLD9y6l+Pon6r9+XrvfTSK3TZlGuporQ35fXMZ01/pCA7+F+jm7i2S5B2HB+O1jIqQFT0rgRRUcjXx3NB33zQjpvRoB22YFAMdgba+cj+6JbVnYFtJikAmkFGxtZuxjwIDhsaICAju+pERYTAC+7TbqLCb/eOZs+c4uGe4udpqCOctizaQ1QAwE2sUZGY1M0zqpVVmLbGMt9nXeKGBhp/4DDqv4EUC3777Xfp+GNO5blXUlTBh7itB21Me+y5M2V17cpExjV/v5nmzpEC1jk5iOL2WvgZcyzWVp7zIBtql9H2O23Kck1Yh2FRba5r0F2B1xgYD9sVL6oNYO61196kXYeJRNUnn3xKxxx1CuX1LJY11FPAp1BnWoIROjBwNWzE1q6INp7vwslT6d235lBVZT+VoupOnTqKL8mvmC+YOBgp2X16tguu5Scgir8O32Nr2mLLDdluL1m6lC44/2J6682PWL4KdV9Q5FiyWOSIqGhFG5EoQoI01NfR4qW/0vEn7UvrrS/jDZmvyZOupJUrsqigVzFlQXbLyTOp/XKHVAEQAUQecnhIVMyjfSccxoD9aqv1pRNPPpT6rS6kK3zq2U89T9On3ce1GHqoVr5F/ZuutHRIekbFgw88w+Pxu4kKNY42dLaCDFQy8CFzdWlh34Y6WrL4ZzrmuPEM6OP7yEi55urp9OXnC6kXpMU4I0V9/pYWWne9atpz7x3ZruM+zz33Ap126kQG1qWANrLVYpkYMccD/VdVXUTj9tmF8vNFVgvk1amnnE2VFatxnYyeXOhY6ghFJqcRFepzMZyIKGcGpsQnRmbF8uU19KeBa9L4CSNchtMd/7yXHnzgWc6qQJS5RD1n+svcX63WqAiJCmRJyYmpxbS5+e8V1AmEhNo72/0ZsASAtXKlIyoGxYiKhQuEqMC66NKpi9fIji1KwLEA9DfYoE+EqGDpp4CogPRPW/wfAzcc8V9POwz9E+02YrAjKqZcdCV99MFXPC65OXnUScmZCKisN5D3Yn0KqatWalQk7eEIdBg1elvacact2HcC+HbdddPo0UdfYqLCJI2i0WqtERVJFs18GFs54YHS7IRKP9Uu02LaKURFVk5iRoVvkS+mnZRRUVGxOhUXVVF2t+5CcQYgmiMfY0QF/AGp/bCCamuX0JGHj6TBSnSD+Lvwoqvoww+/oV69Slgmy87ucqQVApNXlxIJDY21tNvweEbFpfTKa3OouLia9xxkvAkwCYCwA63kIsZyyJGzlwCXRlTYfGBgFACvPVfCpqMio+7ZbV/RU7rfqoBpIiA6TlQEfWb3Cc/puA6D0KjXAPUJk2rTehEcoIaMFJaq6UCdugjRaLI2TG7geZmIlrMtF7vvQNRQL+Aw/hZwu4kJSQCzcjYRSSjJIJBHQcZGZNuNAJ7hfBXiRWFtDnyBpI+MPXHUPts+jeaHT4CoegxwdrcsBqs5swVBOCA0LMI9ISaFz++dRPrJvuskfXRehitcMkSiLwsoNztq9RgxTQTIFvJEo2Vkx9f6CWk+brgGokSFSGrZ/OLvoV+URMF/LSgyPDOHxAdsMeYFkzMsoyV7TjiHMHYghyxLAt/gGhVKeuH3DLgrOd3Q2Ejdu3d32RRWsF38BzfT9dmjWY/Wn6IKIXVd0IfAaCPZGRH8R+Sx0QYEHeB7aF+37Gz1QlZKAXYmszrzvmE+kdXWYNCfSyhpMCXmevAKMyoMMzBSg7M3NKvFiDkj47pw0Ke0TSS1jNwwiS0JerbvpNV8FNJLsDKrh4F5HZJPiX5rwpv8LAGxaXPV3sc9rIYGy+2DgDXXVK9nfeCGIeYI4zksk+kPoiIYBMg+TT93PK23Wildc9dLNO3B19uVTYFLwIh075ZF/7r2SMru2pnOvPpRevLVT51RXRWiwq7Xt7yAbj57HPXI6Up/u+4Jeuq1uZGCOkZU4PtSTPvj9s4zWXztIGBW6YL/sS9rQ93iMHY6hago0mLawQ6QwViHnwWMa/IjyJc9oK5RSbbFxHaaJKJCNucQkE0DD6wFQeHIeKNSf6rFn9TZNfCWi1CBlRVvSIBKTuePOqZRxzkOMEsjtCecqeENSY/HnhjRjYq/nP6cSWPCxFBIMunPI5tkeM3Y53LIDB0TbWoIOmtkTOgw+KUg77rCnQ6YTJgZrEQE7VCkKMqhzXQbM8HroB9iGjg+EjxckMGc44OKP1JwCxn00I3QMSR2j3if24/DSCh/PE+zA0lZSUZIRMbIDFakuFhb81vIGQawGcj10UqWkppZhNieWw0uHzzsQBTXWbSJge/6Yow2iy3iJkJY6OYqERuSei2koDytOBUgdGQNebYoE3CO29ewN8JIQbMJ8bUXmW2tdqWsNRsC+12aaY+vuXjsTaLtSpr6TKzaEShqHzPXvBAVcTDVxs6k38K+YOccqeNJ97YIGo0KFTMjKU88Qm7o47+XOWbPKCsoJCqGeKLioqn00btzKZpRYfrp/hqBUUxsq0TeaYQaxsk5Y0Je+Jefx9BEHT1+Z85QQFsZZD3iRJbyKC+tYtAfqfM77Lwl7bLbEHacAcxePvUa+uHbX6iosJQlltAf7DDyYUAjANm5TN/4mRhoaqJ1+q9Go8eKDA/+7YpXV0D6CbIRXdmJ3G6nzWnQ9ps7kuL119+kM079Kxf4LSkup6L8EsoFwAwNeSVCk+x7yIsK6ezrEOD+qdJPvSH9VMSyNzZ/kiLdEgdH32x97QHZkyXmu03HTQ9C+JcM60paEZ9yCZk2nqjYkHbaZZCfc1MupzkffMEANCJepSBvNJpAVlHS+KUbibTni5O1uC4OXdWcTbAr9czrwZk9N1w3jR568EkG+IsKSvmg3j03iw47aixVVpazjXzqqWfohmv/wVH+PVmGCBGorfV69EMGzRvqqFdhDh182F5UUlLMPwYBd+mUG6R4NfTiWZIhiORW8AkR5ktrfnNFtXEwQrR6Tk533mfuuvM+uv7aGVQFIDdWRDtsJcCLHj2zaL+DRrjo2rfeepuOOerPVFW5Gke92/OlPV06CZ5ulaP2XvpGDuTNdMSxe1NFRSm/9/HHc+jA/Y9ggB7jgUwTANKOyA1uIXuUrLbkoAzNRqmtoUHbb0y77b4DAzi1dbV04w0z6a3XPmFQGsRTRPokNv/QTkSSH3QoiArUS4Cc0Tw6cP9jeNy6detO66zTlw49YoLTgce8uu+eR+nxR19k4idH5VUkGCfsDSEq1l2/D+01dqfAHklGBTJcoLefJv2UNkYOpNNJ2ra3EpWBY1CgpZnls6r7FNDBh+xNhYUF3M9vvPE2XTT5OioNak0wGN9xBR10yAhafY1qbtbChQvpb389n76at4DXDQpfuwLFCGJS4DKyfllKpZm2234j2nHoFjwuAMevvuoGevghZLz1Y/KnW3Z0zHw/JM/B8B4Yz8bGempsWk6nnn4IVfep4p+///6HdOZpF3KmAWpfsNRYrKCsmbsIUTHM27iLLryMPnh/HtdsyO2OCHOs5dYztTPGkLewFn7uUXsNpkGDoxkVCxcs5aySHGSmQEs+OOt68kmilTG3UKNi3IRdIhkV99/7NFVwjYrCaI2KFEIYLglneTTW0157b0fbBW2aeM4U4roZJdWaLdPZBSfZvhH1mTL9dxs1Vy9F9yPYbIBUdm7iQKEVK7nw9ZZbrktjxg7l57I1OXXqDbRoUS0/F3wE1IqyQB8XGR/WFdQAP5P1CIPKWrPuEZva0kx1dbU06bx4RsW5VI6slV6lnC1nBWnN9tlYOfKfyalaOvHEvWM1Ko5gCSnJqOjOZEDoa3p7Iv4QyyghYlv3UpiA+rpaGjSoP+237wjWxYfPccv0f9Ddd8+mwsJKysrOFelB9fvxWysejfZyDYMVTbTbMGRUeD8SGRWvvf4JSz91ywGhLBlORgryXqYgXkdImslsdTbbAle4ALRF8rcI2Ij7WxAPiCzs3Qxgo55Ax04MttteCekuA+vFvxKJH/FrZA7BnlktCAEhtTXagVx/0P7WoDo+qwUR7XHrwh65vikunexFIoXk60uyxA3q9bh7ekli5/EEG4NbD+gTEBZBnzKIjj7SOhAtVpfUMoFUvkz60GSgJEsEc1BUBmwMokWz+T4caCROIb7v6p6CfAIYDqkkDQYC6WHAM8YFz81R+h1RoFoIAgTeof6Ii6Bvbha1D5XJwu8ExJYxYwBXMxvMUnC/8fyQyHq8b34wy5nx2EoRa/tMnlVknTiwhCPrDVxvo97aSgm2NTCafUeXTWzIij+D+4BCECFKzqWcQyLBPgljHtoWfhb9jkiR+YLOkvWgMntO7kmDWjVYjM/35s6zqyRnNSGHpC6EFSm3DAtkhYP4RZ0+9B+eRzAZPWtZqAiuYedky0AIMhntORxgHxYGDx4SazvplebXS+CB1rO1AuFcKF7qpmS83HFLiAxXrwWkHLJGOkltGa7LwTZFCqKzzVC8Tkg8L02XcQziYxRsBccTu6z6cG04O6GBChb4yufXP2pU+GHbfuCadMmJI3gDOPCc21NrQ6Rt0GDsJh6xC40YtD7Nfv0zOv2qR7gQN16rSlSYURu9wwA6/eAh1NDQTCdMvZ/e+eQ7tzBDogIZF/96ba7TObQ2elDGT3aJBlhJdfVNGVka7XU+/rvf07avClERrJTEtLrw88RTigJHAbAVEhURGxsAY565lx5yh9YMooI/Te/G1iKWU35mb5vhk+cWgBXthZOETREGnDc+MN8OcwnmR2sIQ8pZOynCHxkBq0pUhBrfSUC59JrvANscsaH4NFNxhiLRBTGiojWoju+gEdASPZP8bTiGMNAmG2ZRDebM6Azw88AVC8ow46nR4sKhxUFNdEJQcLI9REXGULR1NA/6ObaWrM8zxwdpvN7ytG4j4kSFrjel3cWBQFRuuE68E+8eOTI0dvOgwR3lC1EbIE5y5NrBBWXaqkOFP63YahjNpPI1/mARd58MHArubKCIK4jtbcR/i6hobUzaS1LgGsmkZkL/a+877zmylsxwqrCrOnHOeYkUcfUtt3vzGhUj6z6M2r7408aJCi6ryGCFZFQERMWFU+mDdz6RYto9IPMih1RX1DyBLPVN8fYDRRdtUchMDEmzcA3K33D8SsoLaPz+u1NhUQE7l7Nm3ka3zbiLKiuqOUIZkjU4VOYX5dJBh49jUBdr8sH7H6HbZ93PZEYPyAx0Eo1Zi1iVA5ZmVKRMBLjcOEit2wpRkdezFx8Att1hU86kwMEeY/LRR3No0sTJtOS3ZVRcVMagdm4uIm+7SvagA04TiJ7gMBsCvdyexkZaa/2+NHIvL/0yY/oseuyhp1n6CTUzBDQzG9KGY+/ASU/cJ3YHXy5e4c1IJzvLWpyeoGGy58Vf0XE2omKr7UBUbJtKVHBGBWIXI/O79dyJ5GFtH0BuwN2uI7ahrbb9EwM68+fPp1NP+Ss1NXSgstIq6tWzgA+1AJ6GjxxEO+y4DR/mUEPlkouupqWLG6mwABGoOXJYSn1F+wnrFoegmmVLaMyEXWirrTfl5wYBd9nUa2nBd795uaZQ1kwPgvBnoIO++Vbrc1FtyfiR188//0znnH0BzZ/3A0eco+h3WETbvoe1zbVhtu5PO+8qhY4ROXfdNTfRww8+xURFJGNklbUzPTATGKyghwJ7yOBEE/VdvYz2HDPUSVDdd98DdOXlN1J11epUUlLBpGVIIoTmVa6ma8LdJdrvQhDVUnXfYtrngN2pV14e+zMP3P8I3TbzASYaEJ0fyj/FZ5MnKlBM2xMVBx1wLLcTWQLo14Gbr0cT9h3FkZJ4QRZn+rTb6f13v2CyUbIPkKUSresgREX1v5WoiLAhgT1IqzFjnkc4na2WSU3NYhq221Y0TDPyAKDPmnU3Pf/0W0oa5LANHrzDxjRkJ8k8Q3/cdtsddNMNt7J8V3GJ2GzOOlM5hiSiAu0AyTNm/BDadKDUXvnxxx+Z8Pjum194flt9jDiJIG1vD+gh8meQthq/n6xFu8/k86+gX3+pp8IClU4LSUOXyyMgF7L+tt9hY9o1QlRcTh+8/4UnKrogE2jVNGglkEWyF0YzUbG5a9+5Ey8mIyogoYUzjz2x8MrmS7dFVMxOISqSDRowJltLx580htZSyUYUvd9vn6OoqnINKi6uUtIPmYeIMNXAMmthinykLWOAvCbbJevawERd6eorC2HSQLSigU7587605pqSyYTXTz/9TPfe8xjNnv0mdc/Jo65cFBs1TJC9ovthWD9KbuMj0kPz0Q4VAD4ToZg2Z1QcEZV+OlmIivxeZZSFjAUlEdBOBkHN7zZ/c+VKLlh+UruICj/XXQS+yvUwQK1FnfEZfCQUku9d2YtOOB5kaiH31f33P0yXXzlLCKbuWJuBvJwWfRYpZ9hqFFtuouExouK8SZfQa6/OocKiSuqWA5/M+toXsQ39WVmiEt1toCugAxB6RiQBTDY5Ggv+QH/BBwShYSC21IaQCGysMSl8Lj4gR2WvXMnkC0fEK5DJtscF1qhPo3OH5X/sDOR8Lc1wEMYtYmHMU3LBXkom4PlEXqmDA+eZXODn9uAynwPUX3YguIHS1qaOXnpK4HEjLfQkEAS1G/liMjkmmYP+NVBf5oP4XIKbcKpFgJMEQWqGxwe1PWDnm3RdGNDtzjOqaoCgUdzDsBg8igHqQthIDTcUk5Zzh6/fg7XN9Qu0loeTk1IpMbQZmRwYK54zyBoCTtGlsyNlwrNtXPmg1XNoZPMz6SEJ4LGM/+j+IqAD17ZhgDrmyyZIZ8n0j84j26vTvFgeO85kUAUKtVEmQYV/YqytgLYFdfisdvORLPROM1dAqHUyeSfZO3A2ksLvDbK3WFs1KMzjfbq+g8wDF2Bk88bZNXnmpBo9PPaBDGZkCNICznQOu4wMzVriQuBJnajnHMYFuZ86aZCmkJC2FhCgJHNLWHKR8PJ2iiWqlAyMbBPBmNryCBOSAAAgAElEQVT+ZZnMsj+sdB6A9ZHZP+vPP4gKHfkunTvRbefvQ2v3KaEPPl/AREV70vjDiYMNb9DG/eiyU0YyQTHmtFn09Q+/8ld+D1GB36Fdx43blvYbvil99vUiOvz8u2jp8nqecEZUcDoQDJSCbxroZ3ue+Dk6c+wz/BdZIzMeemOVnzN85v/O36tIVBRrRkUIUKrD5dobrKRkXD484MWoDttww2u4A2E0ejtOVMhYZAJUGf34O4mKMNrSRdHKTiJsukYyiMaiFKKKv6Lti02e/zBR4SxprG8jzxWAhBHwz/3GJnvwZL+DqJBfW0R9Zj9ZBANvx1ZoKlxssvJ0/YVF5uJgloHmYef67yQe5Phj88IyU67jreUrR3GQsHMSl3FaRkU8ws//+PcTFW5IOdtEXc6MNWDOffAwkZaLY2Qv3k81GiFOVPhniGYumT4kroHDh0WjOwAjBDn1RpHaCG7MY3MwmH82V3w7w4jXpAXZmpX1zxxO8VQizj6ITcFVISl4VYQej6urkmbX9FCt1sa3038/BBHaIipcv2WsteBA7aZImMXQXqJiGV14wcX07hsfUllJpWQEMBCO64eRXtqSwO4YYWoHUhxAWgdi7MdyrANYO3jnLWjwjluyY81FtE87h376cTFnd1jhaDjhNcuX0ph9d6Ottt6M7Q8kWy4491Lq0NKZwVjUkWDtd9NylYFz/06aVWgDIvHSiIqq8r7UI7cHbbbVxrTLiMGsm48XAJnT//JXWvJrDZWVVipJ0dMVlEW0oF+Y8ld0TdqajxFPXNi4idZevw+N3DuMep1BD933BNfMYKkr1WJHb6b5bTJnJeoJ/+MxglOuh/PM/hAnnF8O7fKHGg2jUsjoP0dUyDT3/kjq2k41E+0jKiSboBvtd9DuVFYm5Nfdd91H1141jQFQkE+53XuKjm9jPVX2LqL9Dx7NNSBwwL7jjnvpkQefpdLiSiHKGISM73WR1RtpsUg41dKa61TRuH1GcP0VIeAepdtve4iJkh65vahLWDhZ7RC+B+CyazbRkcdMoPKKMnftp59+hk4/dSL1qV5TZJ9YViusuyBfBUiCwtWHHDmK1lhTJNW++mo+nXLymdTc2JEzXXrlFZKrwRGLJnc3TDtAWqhj+NSRofEbNNuC5ibabIt1aedh23J2DZ7vmqtvpCefeJ56V6J4rBBCkQOuyzZTv6MNooKllRobaEnNYjrtrEMZSESTkBl13tmXUe9KyViCLeFsB75sdEzTiIqDDziW+lSvxe2EHQQJNWG/4VxHxICZL774kq66Yho11HdgaRTIHnXqFEoKWUZFNe05JppR8fCDz3KNCmSaccZWsiOfuiqS5mboZ0aGKRGUFRAIcxYlew4/coyrr/Lll1/RpRffwM+FOdunXyXtu/8wKioq4Mt+9NHHdNQRJ1Nu9wIqL0cB7SLK5meHvfaAjgBlfpKY5NFxJ42lPn0q+VrIsgEp1LtqdSpz9QeSZJlCQxbtlnA/lzMC6i3U0uAdNqLhIyDF1oUlES+beg3LGKHAPWpgREgy9QuY1FGiAr9PJSqYmBEyNumVPharRlT4UCPb+9Qf4YyKJtpgwz4JGRWrRlTIem2m/hv0obHjRbIRffDoo0/QRZOv5nlaVFRO2dm5EpEqcbuOBJBV5eseZAR4aTR6lKgwP8xnE0umsMm6LaMNN+xL++w7gvLz8wPztJKWLq2hOR9/Tm+8+TG98cYclWVElLcA6eL3IsqaoV+OglUYWLfDGMmSMIA2p9KIipOZqEAx7TLOqAhNoQF3LoJdM+dAqp584t40YMA6fMfPP/+Cxo5NyqiwBvmrMkGh2QhyfYm8xz7FGXlLfqGpl5xI1dWyrl555XU69S+TqbS0L/VABlFXBGRo+J9iLjaWK1ibvomG7bpZkFGxjM49dwq99PIHVFAAubTubNvCjEDn6wZWVUZQ5E4lA6OjSv0AQJXIeaubwDZPde8h2SM1wiQquqVZtOtxvRUtmb4M3rdC0RblziRqE3AB83s8aNwqUcGmJe5n6FUigJQCviimrUSFjTUkmTDfZD+Tunn2WeS8YeCwxlk2s46VAL1ythIQnbNIGGzuJJJCKl3FARTosxaA/kLMGKCP7/ssLMn8aObaOeICikQzSJ9ODNpyuxAkabWMIM+k0fOOFDXJMdRf4HEBGSOZPQImi3wxrg1yKTs7i+dfXV09kxayBYhcGP9XpbbQHs5C4VorkBKX7A0JEBFQXTI2OlGXrK4u+l+yLnztC3yP54Lrv7Y9TCHRBbfAf5tXKICdEYimg6TbmADTWhsjKHof32szdqpWSFF7ZvQ3pKxFTktk1KR2qcwHA9atzSFRodg7y4JxfT87M6nkEsB7fk6VAIO0lye9E40fvxlKJMkzaR2YoLgK2wAt5J20D6bVvUsjlXAG5T28BZiwl5hn+aWEoZVaJz7TRJayPKsVtednMSKIyc4VTIKGgYGcNaOZRKGH6I5OAfHo8DKVqzd9F7s3n9Qs0Anz7H9TRgUW/0G7b06HjtqCXn7vSzrt749oelyiH+TexCRdd7Uyuvq00Qz+H33hPfT+Zwta/1HCp7hOTnZXuvOiA6gwL4cef/kTmnTzv3hygHCYdvZYWrNPCV14y1Ncd6I9RAiuWZjXnaaetDut07eUnn3rczr3xn9RfUMTQarquZuPZX3R3/O67u6XaebDb7arHb/n+v++33iwwFhxYZLbUUxb/Ct5hYs0BMITuy+Mow9BY71UCDxGgPO2iQrrFzlYpYzd7yAqolFiAfOvTrCLElCNQ2jRskFo7YAXQT9j0aXBAEcvoaBKa8+QAVRpV5gltTN7QAC5fgvBaCv6pMwuDzfXqogjseGAi9OS/JJPHDAEdjpliLCxW+okbmc6gSI/4wHI+PUyxzydqLCsmLCt4rynTObIQwVAcCDz5VjqAGBN6os2iYpgjCQRIqzb0pZNEnfcIu1dFI/KYkn3xddHElERLm75fmTKtkpUeJLCnlWcGzUVHDUg+pDsTOrGGZ9bmQfq4NllgUVH5f9mRgW3R5rjn0Pc8FUBejxgn0aSZY6/c2rc0pDxssyn0PHjSI2UQMvIldNsV3xus11pH1EBgPCbb751BfSi9sTWXWhP/PA2NTbRk48+Q19+/jVldUW0Ig79cHLDPSSst+HtBEcGdVhBhxwzjqoVhHr2mefob2eeT1Xlfai0tIL13HF4hWMJXf41162mcfuNYlAXUZQzb/kHPTf7NSorrqCcbiL/Ee4zYpJT4GO1K8hgyJR+mkmPPPAU18AYMnQQDR+5oyMpsD5efvkVOuMvf6P8vGKqLOutBX5zJCIpLWI2Mg9lYsaHEz4SSz+t34dGKVGBfvruu++ZwMDzCRnTHm9DvrSsZjk98ciz9PPC36hrVraAZYnzyNtYt8ZV28kOHBESKBBB9K2JN0wOeIjIajujAtJPsWw6s00Jj5uKj7ejawxok2yCbfmAAp3uyRdcQh+89xnXJmEwNasb769ciHnZEjrwsNGuqPann35GZ581hfLzShy4nRYlljRgBm4urVnMEk7rrSeFgpmAm3Q5UUsWFRSgZgKyNVT+KYhoQwR3VXUhTdhvd+rVS7T78Xr9jTfoxOPOoL591pZC2N17ZhSbx/ODmF5nvT40cq8h1D0nh9fYXXfeS9dedQtnU5SWVGqBZCFgAOQlvdKi8n1WWfCriCNiC0L2dxAI2wzekHYcurXLurnowkvp/XfncnuYNGHZp9h+o5eXd+X/BnBdrMlCji6vq6FDjhhN/fuvzd8FAHj0EX+h6t5rMOkoGu1qkGNrhYmKuuV04KEjIhkVTFT0WZsJLhAQILdq65bSEUePo402kpoOGHMU177qihnUI7dAsgq6oCaG7f3/GaIijUBbNaLCDvQorF1Df9pkDRo7fjfOGIG/8Phjs2nGLfcxkYJnlgyIDlzT5dJL/k7PP/86ZxYUFZWxJBCDkjxkfs1nEhXS16ecth9VVgoZ9+qrr9Gpp0yk6qo1qVhlzTqG9VMiI57s+Rro4f1eicpfb/3eNH7f3Vg+CLrd02+5jZ547GWWqmLSMFanQkCXtoiKeZypI1Hqq05U2NmvLekn61PbVDxeKv4O2vrvISpQ9BcAYgsdcugIWne9NbjHly6F/byU3nrzE84cQPBA166wnwKicd0JRiFtgMK9IrpvSJ8q0KXnC/6ZM/pW30AAeCaT62tp+fIltNZa5bT/AaOpqqoicZ+DLf/hh5/oyy+/o4/nzKN33v6UmpqlyC7q8AC4w39h953+vAJuaevFnsh8Z8zZSecdHsmoYKKiYnVPVOizhIE8QgTIfBJJsrpEoqKiArWDRPpJJFvDSe//IdJGWqQdYJ4qXsCfxRo+47T9HAnC2TD7n0ClZatxnQqQKc5bU/kTqU+hdSVWNNOwXQc6ogJ+5Ndff8vkAs4RAn62x1GR7yxc+DNNvew26tolmzprMW/OkFDQNQQwYZJxFjW5WmRWNDZB3soKY0ezR422wOcAMx2wa5IxySGMiRkVkWkY/kNB7DA4BuPCUjJcq0KyFwTwFhkmDqBUAFwiwO0MJgFCbiQ5e1UAfHxiEkT4Dvqba1C0NDtiCp/jnp07W31DtVGNqE0KQkiltbTOpdVuZCJHC5xbW/EMeL+5SUBxlk3SGo2MsQRSi96eCsFkEjl21jGCCG2VvVrqPDBQ3NLMzyG1ObRWJrI8ginEtQaUqDC5VFfsXGWtkG2Ma1mhZsxZ6w+f1YHsFiNzhAhO9m0UHzHaUscPRIU7z7sfyh5uhadDny++r0VWa7B4o8s42dpYNgyugQAu9K3VEZHpKAEFJlkkW6ydO+3cK31vc4znpK4d7BEIauL1xsok8jd+4aXKgpYG7Y+sdoMxeSPyGJHdJ414WFWigteVSf1G+lJrdmYMrLTHZbC5DCtk4kjWhNuhlKxw0pmKb1hR8aSdzH7tSBoLulICj22C/tBG2LL7eDxAPP1vIirw/GC+sOAklU3S29p64XcYJJAJYiDAUCYv1Lauhc9BIFgBlwZOh5H0wi6sA9eBWVM2Gm03TX6LhdcJEYCil4b2mXRJVld1btsCnBMajqwPGOT2tqM9z/6f+Y6tcGMkW69RMTLMqAgOVaEhCA93yViXahFy54jBlUOEPGEU2IhKKIWQlH1fUqgyeyc5Pdvuk+LUpBIL4XHUJD+kyDE24zBNVR4iAbQ05yIEMt390oiK+EQO2s3gV/JzZEA4GQBu2mwKr+8sXPDlxI72n6f2nzj74fhizqSBLXAIsImZA+MNvYLTgdYrzx6bQJEUb3yXXfGEhzXxwMw5l05UOFc6cj0X9e+xEP083XFOJSoisIf/fSj11R53XJ47API16sJIipAsck6EOrFxkk9sWAzo5LmXEAEfEfOKHx403RdXszRoc9pSQfGEp00CoKzH/28SFeZgar+7KdnOvchPKpuzakTYzwv7IbNPcKSwOSWAuU9F19FzBeAZ8GjXJIova/mRt9USPcQRK84dsguL9BNqQoTST6u6h4XNhL77jBv/QR++9wlHbmehYG8oj8EsWDjnxC4wUNrcQhtvth4NGzmEsrOypIj25VfTc0+/TJXlqA9QQt26aQT1SuJ2Q5f/pNOPcEW13333PZp41hTOvshDQdUuMU1/9UUSNyM275DCQo2KfpEaFbdMm0kP3vs47bX3KNpr3B4sRRO+cNh9/NEn6ebrb6Oq8moGUTkKmwsvesYpwxk3e6SjZktM1rNYObQnzKhY1fGJf/+XX36lm2+4jRZ+9wv15FoQGKMkViy6KMTRtsw4y/eXGe2OOHEb0UqNii1bkX5yxbSNXDPnPqVCBT/jKq9h3zPwEZBNcPCRo102wdtvv0PHHXMqVVb0pfLS3h6Y5GjEFqqtW06bbbk+7TF6Fy6qjfl6040z6a3X51BxEWSJoIHeWlZFdGSELBAgdsM/rUF7jRnGACkTcNP/Sc89/SaTBbm5Vjxaoif50ZX82XXE1rT1oE0iRbJBuFx26TU095NvhahAtkesXQJaNtBuowbRFlttxHbq519+oYlnX0DzPv+Oa1swSZLVzZMkaftB2jgkaQ0n7RO6PzQ21tPwPbahrbfZhJ8REj8Tz5lMPy5YwmPCkkxcxyTqb1mv+ndF/kM320inM1CFWgt1y+mgw3en9dcXcuiLefPosINPoj69BfzmaGC1Y/HHa4uoKIFcHYrcrlhBy2trKLsb0RFH70P9+knWihXXnjn9fpbWgiSNZEgJoWvST4kZFZX9qFdPZFSkkY3J1kK0w72N0UmUStYH8cixC0pkakNjHS1d8isdcNDutNXWA/k6KKz99ytuptLSMtr/wD2ZwIB/+cgjT9AFky6lstLeVIoC2lr42opw8v6l0RJxe4ngoqrehTR+n10pv6AXt+Xee+6nq6+azkQF+g9ZNqnninYaT1sP6/XvQ2MnhLWKbqNHHnpOatFonYrWSEfIXe0yzMvbTbkQ0k/zOIukR/deah9WLaOC7a1mUI3cazsKi2mfx9JPUkzbExUJwd56DYDJ/QdEa1RMu3km3XfvU1RRZmssy62xpLMyfAhcZ/w+Q7novZ0HUOD89NMmMRlVUlRJuT2xH2eJLC1B+iaa/SeAlb5izo+AsrIfsusUgj0O4hTigkFQ4AxNTUyIL1u2mOobltCIEYNp6NDtqKysrNWgFIB6ixb9THPnzqfnn3+Lvvj8OyZEWcKxUxcn4SJtad1JQ4uxV8CmnxerUWFERUEB5izWhjy71S+wKGP2NLmALAj+TKJi3NgjKCQqpEZFfG+R/kNrOduAI4L1bAxbwNl8y+mUk8fRhhuuyz/+/PN5NG7ckVRa1pfJFNTqscLZVmfOB/+hfVGiop1LLfVr8+d/S0ccdQ4TuNkcdCLZGKYj7wBangvArRSMXYki1ShqrRHObFAA0CuxqgQA2o6+EBAcuJRgVfGzlZuSQbZqSGiGD5BBEAVzVqyt1pJTgi4ERxk8RkZCC7TxBYsTnXpfg0XstNzRiIpwCkr2gcSGCYYnxZQ9MC37jZHBVmuCr6e1K6wPuG3cL03ct5I9pnUiTEEBwHUgxcQYi14Lf4T+LNaVqzWieICoMnQSkkkzPUye1bL78Rws+aT9INiwrDuun+DWjGTSICOGwXpul8j38G9A/juQXOpRWJS8RcJjrXJGQopvwzZI15HMH0+qZOIYcjb0bQ/qaCgAnTb5ZWuO+d8pWRVy1pNn4zE3CWGVueV+wtpgkk+IjHA+2L/5llrInrNtIM8FIkh9Jwbsg/swtqBZLrpw5OMQ2E94wAySJsx4T/j+qhIVJtfkyAq3YNKyzfUsbzVQNOtczsziH4Jc5OwzrnfSIpkiMcIl2Lwiu4Ksh+DBdMvgean7lSzoKL4olT90Xf5vIirSJv0f7/9P7wHbmVaNqAhtrTDefrVEPks0ylrwyrmGgVMWsKHWs6HjGPa2vW9ORXwD+H1ERfJ4Rg+ssKkm9bSCNy9s/khzFYYZm5T1RzRqUwyzd0DTNi1rhRymEiyRbSCp0y/q5Moe4NuU/vPwYC6bthW/lpRPuUak3dHJkNgiiSrR+wfGFFEqSS98hZ0P1RyWDVKLWen9fBusjxXYjVyQ3fmEW7SHqEgDh+MHCAC/IVnWNgrcFlERn28hIdXWAUYGyGHVbp8SdFqPQO4wxtuV37S0fohEM8tzCHGbCdisElGhETqc1ghJGCu6x0Q2HNBgjrt5klA/RB9O5lJ8jsu/46RpWjSF9VO6BffzKZV/C34shFkwOtqXVlw8brvS2xWseZvrXAwwCTDVMQpII/zEbB/uzVEVesC2/mkPURG2L4yqUgMg/d8GUQEgbJugRkV7dsu01QOw9vprbqaP35vLMk3dshEdbPJL9isZs3CNWG2ICQftTv0HyEHZFdHuWchAca88K1IsUXKwPSjmOnioL6qNaN2r/34DffbxfCotFoCQJf8CH9A59rEH5YPhCiEq1hsAokKAYvx72s0z6Jv539HJpx5PRUWFPH8hX7Js+TLaYvPNee3VLKuhmdP+Qe++MYcKC0tEP18jCW0ZuH3QMf7SiAiB5RxbgQdxiAtrVLRnfFr7zk8//0zXXnkz/bRwCY+Rk8iK/4g7ynfcf5OogAyOq1ERtCsWVxjdReIIsn6aiqc7t0rmErIJ9thzR5YtATlw/XU308MP/otBekTFi3SFjx5EQcGs7I6uqDZu99JLr9KlU67X4tcCpNuBqT3jBh8NhEl94zI67qT9HJj97rvv08S/TWXpJpY/y8qS1HN9Bpat6pFN+x0sRbAxZ1DforS0lOfqk0/Ophuu+4cUoGZgONAbV0308Pdo63PPvUBnnn4eP7+TnUqQjGrPc6Xa8ciYqX1QEATg9267b0Nbb+trBJw78SL6aWEN96/IayFQKcVXcwMvetu20uI2Hn0HIPGgQ4MaE/Pm0SEHnkB9q9eSgto89p2DmEN/FSMqDkjJqEDxcvxeMnEaOBNntdVL6eBDx1F+voDty5Yto5nT76Q335jDRaWRDSZRyCAqpUZFElGBouJ5eSh4vGrST9Znbk83ty8NoGmNIFQbhT7ML8ymI44cR2VlUvz8rTffYVJ3rbWldsfXX39DJ590BtUsbXQFtKVvpZaRtac1oqKyqoAm7DssICoeoOuumUW9q9agwkIUJu7WJoDc9pyVbIP1+lfTmPFecm/6LbfSQw88QxXlkNwriBWa9ldl4rCpgetyxImK99/7gqXkUExbIl/b9kUjc7YtouKHZSxNFRIVbMkj/piAJElExU03Tqe773yUSkqMnPVzK+4n4ay04cZr0867bKVF0uVZWArxtIlUs7SJ24JMQwGbrdaA9/c5gjzDQET7BNMzJBu9ryt7tst20EhhAxQBnoOsqK2toZqa32jp0l9p7bX70LDhQ+hPf9qQSkuLtS5M2oxYSYsW/UKzn3qZZj/9JtHKTtSlCyTKRCIKxYNTX2abQVTUL6Pzzo0W0w4zKrC3iHERYJkLFKsciQBdbREVq3NGBa7TQWVa4u0yXxF9ZzUqjFSCjWlubqCTTxrriYov5tHYMYez9FN+QTkT5Hhmify3TAA5e4gOf0sko6LtNdb6N778cj4dfMjp1Cu/lNcKsnEwUUxihc88GlDFJ0hTSlAZoJYWISAkkl6WGcvCqAoBA9VK1lhWKvw17P3x85t5+0k1KsKnCAHJDsgYMpCch1YxFQXCwzMb9mvIGza1NPHz4W8eJ80K4PUbOX8JUSGZ7hI8wutAZT2tboEEr+mZSwtv47tcWLhDB8rKyuJ7WDFrGUsBqfE5yz51JILUj7WJi21rvRu0C2sB17AMCJuv0eMiApGaJRtao/6N5DK7L8W1hTzAeBh5YX0A24HPmXzQAthSmFukqJAJLddERonIuJnMkhAtWlha7Y0V4Ma6EJJE6jIyiK9yU+lrWxa3r63RpDLLcRxI+p7VJ0C46Nka73ENiTZe4fnOiNqMdW2At0pfCPkmtTosswL34mwjLYLOs0kJhThRYTbBfCY5F8lzoQ9DjIhrhahv5WyyFtcWaxZ98b+x/nQcDV5sDS8xwD7NnsXfl5OlBsBp2/m8HcNA/e8EF+LPOatfsyt0KDGvrfA7MnyY0FSYxhNcklVmxGMm+hRgHgG2ZkRF0vfD5/pflVHR1qT/4/P/qT2wakTFHkU1bOi5yDHS2dQ4hRtdJsga6xsuXCZGG2mv3snJDFyMg46ZwL6yymC4lbF2CzpyMFJ3lTUnk8cqAjKpceGNxQAV1V5kI8lpqWFGgAc1ZeP3G7I4tuLwykYVbUA0FdDa6UFXM/a2+XpjHr1nGGGgvos+qAHOYG11Qw0YcdNUxHjiHnAsOFJCHcb4dmDOKOYAdB75eZGyCWeAC3kpUK5biTn2cmC06CWV8XJArL+LjTEXqtK0UZfiyN/3M8zAWyZUOLXWAxJyxRWcXmovuZ31h+hk8qEgGJcWHR8maMIoGMfziAam9TH0twW0D0GNYKty0R+yA3m+xqcMO4cv4o2GPZ+pQy+dGXwnsiPFJjkzVfYFfObbb9dJrgfh+yuTrIgSTxqPFiHEok6CdwvCpoYt5ToE6hSxExMhQO1Xvph2W1Y3dKRtwHg96Q+tRVaclolG1SKW32JN6IzTiA9/oJCLtEUcYf6xexPITrTWbj4cqBYyvucio7hd0TVv1+E22dQPDhDyDHFXRQ4mbjrrRGbHJrpQ3L/jJlNXhlvPdmgJ53FSRgVAszPPOIsef/QJys3xxaDlRimGmeRwgcLSqJlQXFhKvaC5npVNHTvpGIXPaIUjV6pkQ8sKql69gvaaMJzy8nqyMzhzxm1028w7WfYJQHF3gHedtSg1k3OQ56in/OIerqg2+uepfz1NN117K1VA078HyI1WQLxg/9GVrxkMq0UyKu644y4auvNOVFpSwv352Wefc00KrIXJU86jtdYSIG7Rop/oxmtn0Pdf/0T5vQokAj1osxu6GFHhGS6/B+K7SdJPyCS55upr6ZqrrmfwQHTt08jkYF5xxm1nBjMKehVyn2KsAFo7KaHIpI/FUfMJVPc8I1PNwGqkGZShQtIlJONsJTKIlyr9NI+j5UUCJ0UWJXOpRFudAbomz1nbo7Esm5obaNTeO9KfBvbn9n+FItonn0VNjR0Y3I/UZlDQAHMUchnD90BR7a15Lvji14upqLCUC78zURZb32kEqEUC19bV0PY7DqRdhkEfvzPL5Vx91c00d843UlA+IE2MzBLZKimC/f2CBTRz5q10wgnHUk5Od27XFZdeTwu+/ZXB3LBdSb8H4XjF5VfTs8+8xkRFa8/iNlkbhaSwa79FxcyqrDoD6fwlEKVfT9tsN4CGQopLawRccvGV9PEHX6YSFckjLb3v/JCgJovsJc1MVBx8+EiWrcH35oGoOOB4rjHBRAWyY7jQtQdMzVdkwrSuhg4+dA9aV4tpz/tiHtdNwKhFkTwAACAASURBVO9LS6uUeBCQD3N/ydJfacehA2nEHkN5/YntWETXXzuLvvn6FwbBpSA7QKCmVokKrlGhNs5su4Ewcl73Gc+OoFilMZJRkf7zNX7CvQn+scmhbT9kExo5aqgW2xSfC+0CsXfzzTPojn8+yGsKmSoAIF32SMq6DtcKohux5k4940Cqqirndr322hv01zMu4hoVBQWlLDkIm5v4UkBPzFb0hiGQi6cFYLnhRv1or7E7874GUOyWW26lhx94Rot2F1Dnzsl7C64FUmp91GyYIIQ3alxMuehyLp6OAuK5XKS9SyqR2ZoagmVU7Dlme9pGibyFCxfSOX+7kH75qZ5KS3prDQ0U005zQCVbJ8yoQLshKWXgvyzbdIOLSNOuXaP1QObN+5ImXzCVvvj8WyoqrODC491ze3I2hZ2PDGyMjlFwn4ysa/WHgkeJn6Xi443PDURvbm6kxoY6QsYnSAMEONTVLaNOHVfStoM2p622GshSe5WVFYnEBfplwYKFNGvmA/Txx19Tt265TFJ1dNKS0buHUcVcoyIpo+KU8zgToheKaUMSy2mSe1Ca+wtAqp5xMfdPYTLB16gYP/4oKi9fnYoKy7kod2K2aPJqkHWt0q6of/HnUybQgAFr8/ufzv2MJkw4WutomPxdssyk7On1tFtQTBt+5GmnnUkPPvSE9BfWSkK2RyQwS+0LbC2yTHJz8ykvr5i65fRkG+dfMYnbIPjJTxE9g/AbKXOYyQuRRcJX4CvCv2JbEIDxTJJxYIAAswbkM2mjZwYDhnEnUeqwugCSpW4a+fC1ACBDJhXvsayO1t2wrA5fb0KIg3BftPWM7+Ac1tTSzDgHyzQ1i0II4zadOqk8qMjXYB5JPRIB9y1zgIH9LlLgvglZKBZxjzYjqpzJHonINxAf7WFJIC1Ez3gDEx5NTH7wPYD3KPDPQH1TM98f/YrP7Yzncv7lEOc2G7HHMpqyXTnHTrEd1CCQvuUTBp7Jsh2U8MPvpEiyAPWMQSiOIASI+ttci8aKiktGFv8O+AZUalRiyrJvrClCIEobOnWW87rPzBFpbCPhgyfQ7AfJAMJLsj98xgUwOye/pWPFxFbHDi6zBVKE+B1nkaCeAsudyZhIcJrUIeHZH6kJIW3GF8J5xrhSYyPvVUw8NUM6TOu+KOlhpIXDqDjjU+pa4MUklNYAiQQEKgGGVnExd+2MSKCEuYJW00T3aM4y0iLXaKORbIxvBvMYbeM5wISQFAIXckJwTPs72RRqJp4G61q7Qjse/x1jZpp14R1M+VYcO+G5HDdBBuuGZ3qb/nFc5X9aRgUmsHWO29iSez72rkRQWKpVCAaGRtCiLzkKLDG6xutKpt3fQF9cV3TR/ICmtlkNuU0oYzfT9W7FqMlClw0JjH5LUz01NdTxI3XO6s7ahknPwguupZkaa5eyge7arQd1MqezPaG57erzf9eXbEa3N6MCDphsRMauYgSSI/uCzSHSXANMBDy1VFEXjRAAxa44kaXdRlaqAhuaVhhKC4UMZLi82cFMOHHywcJSKRnbMyhOiAojJSLrw1K0AvDQObiQYgkLQqKNunGsGlHho/UyDj+xKRAyvdJN0f53zLcy+jZmiNwBC81yPBpVYqmZmaCHgIaW9ijkhGd8tRu1+4Lx0dTIIFhe+ziEPHWktBNNF9SQfXFOZPD8r5w512j2ENAXeSKLlvJLTzYWTrnjTc7XZ+AURoOD+SbmtEokhLuvZR4YuMDSE363CJe5+sf6eVTL0Nkke6hU4iHciUKnK/YD97VVJCpimQjxLTGTpFBvwOag9lUQJK0zMGy30AJJe6rpMmaA+SHY6/5uH1ERtjmcxyFRYSRW/PnYr+HJGicq2GXSpw7GO4jYjFtmIxGMrGjTckvuJ9sdcfa8jJO1KW5OI+vKVkikXkIMOInI0FlEVri2Qhsoe0MmqOCvaQcYsynsSaxoocbmaEbF8uXLaOLZ59GLz71CBXlF7LgCMGsFr+CnQT8AUMT3ATQDDJWDDBvroDu0lbC1K2SeADDZdeRg2nLQQN6nFixYwETATwt/47oQvQD6d82OShThd81NtLx2OY3bf3faetst2CH95ttvadLfphCt6EKF+cWUnR3I1cQHNmgWWoU+FKklT1SIZMtyLqKNF0iKv545kRYt/Jm65+TSlltvTsccf5gr2IlaBReedznl5Raw/BVLK6nT7Jdi5MYeRY3ZpzSi4obrb6LbZt7BhXpB4PDhJMFvicwoLWYIgAXtRpF0SGlxdGhiYWQ9JLpTmScqzLKILZB0b/apXPCAzE2bjz4St60aFb+TqHCJHx4+FXOnp5/4uAd65zjElpbm09j9hlNhYb6rzXDVlTcyaYKIeBB2iAYM+xgAFOqk9O5TTAcesjdHxyP66q4776cH732KpW1AJDFAkzE2KZC6HvgbGuoov6g7HXToXlRSUsx9+8jDj9Os6fdSeWmVyB4pOB2XrcJ3H330cTp34mSadds0WnedtaUo9wOPSVHuEhB40MeXdtnvwyLab731Dh1z1MlcQBsyNxw93lp2SOT5UiQy45uK8xKSiQoA+gO3XIeGjdiepbXqG+rpxuun03PPvMHt6tlTi4K3apgC+6f3s/3cgluaW5q4EOwxJ46jiopSnu2vvvo6nXna+dSnN4iKCuoGosKkn9SQO4CKiYplnJHROlFh2bzNVN9QR7/9toiLaw/efmsXmTkPxbWvnE51dSQkYpcs9uMR2b/nmKEuwwuR/Q8/+Awho0KICoDAHnxn0COUFQj8MQFw06R9084DdvawJeCDeWRuC6CGwtr1DcvomOPG07rrCeBpr1deeZVOO/UcyutZTGWl1VrHBxl3coZLA1jjRAVA5hNP2Yf6rtabLz1nzid0zFGncUYF6olIFp0AJxmvVoiK8LtGNAwe8icauktYI+Uyev+dz6mCpcdAVKTX9wHguf4GfWlsJCPjNh43ZGT0UGnCtKzy1ogKJukbaunwo0ZH6qLsO+EI6l21JpUUI6Oih2YBJdkajJlkD4ZERZt+TytfwHqd/dSzdOUV11N9/QoqLCilXr2KWWoOEpBC9EnUKu8ZfC3vbZqPnxzo4ekW8XPYuPP/zzz/+F1W/pK56cG3JiZjYGMhpQRCFCQG/ocm7jR0OxoyZBBtsMF6rg6VXRFFuGfNuo9efukDysnJYzLRAFDXNTFJq/YQFcgWMNDSb7fSNwK0SVdhzE86cYwjE1BLB/JMqAFSVFglsmdJQQvBfpe8JppZ+umCC450dTRefvlVOv6Es6m8DAW/S7k2kmTHJiwr+GKNDTR8WLSY9ll/PY+zUXJ7atAG29DQJvu5KRKZMs64D0hA1NxAAXbx/YI1rZdw/oXWXLGWhV6yzI9Yo9UOWFFnXw8iCNRT+2l4FgsVaHY5rx7dB2z+CVGhQYb8ZZAbVnRZ769zQwL2fD8a6M9BhArQhgFFFuXuvBkFMqESwDNcpZEkWFCyESxDAQA2Z5xo8WzYJexllrnAQY9KiIV1WHjNMEEj14/aKSGfGaRXSSDfXiEQjIBhzAdBkiwVjUwOFMEG6SR7FPgCXtNhMUyH25iN0JWsYxBmj+CTMADWpH+kXzSrJsiiwPthTQGTkbd6K0ZGCaEkfSlEAGTfkI0ktU/8C42Ss6AjZnQN+iLumcGvXkZJxszGUWTLQGIBiJdsdB5fDfS1fT0kMlwBec0mCmXQmHCLERVGP1u9Gpn/Wg9BfVAmldheC3nl+hVkARcgX8m2xsgMmw/hHAVmJVu7kFyCE8Xzok1G1o9xiBPC2nPWhuGLJjsGjDfIHjPCiHEjK6gNIkllrFrdK0IiwR8hIjJWcav3nyUqYqoT/9OIioblS+ibD56nnLwSqlxvi3b7FQCZFn31IS35cT4Vr7YB9SpbLTGiZMGnb1Dt4kVUvcG2lJWLgnwx8GTFCvrh87eouaGOevff1kcBBC1pbmqkr999hrJz86hi3S1o8cL59PPXH1NR1drUq3KNzEPbypW0fMlP9MPcNymvtC8V912Pr7boq49p8Q/z1CWJbTQdOlBOrxKqXGczXsi1+vuWZqR/eSC0S3Z36lnSh3qV9eWFzkZtxQr67fsvaPEPX1FLSyPLQmAhZ/copOLV+lNWTs929+t/54urRlSMLq7hcWGWXnX9OCojiCTTThXjmHjQk40IC140An1mgjGUrJ8Ysu9aqCs+Z8QpFbCKHS41WGbUfR+q+6n2LALv2j4fvOkxUfudB+iFMZbNASCRRILGojBiBZNCAJa3Ho2ytvbG4psT149dQyIP/MbV9jyRtlk6qDhHBoL6dGDniNkhVNNYo9dXDUJ10CyywTsbmYdY3AuORegouXsFlIO9h+fDdS0yQhhj74zJRhFs5Rla5cFYdNCo/IzCz+Kky7WQsmvFgBGxkqkn6vZBZzGcNxukZfpGtZuosPURc47DNaQLSR44gkFGC3+HDg7Pp7AR/AD2YwHg+XKh6UsDe0JnXH8gR1FfF8FdLIIjeTBR3YRo1Hxwcx7jIKJSbEc0MtEDcplEReh4y3O546bY5Vhmhj0qZztYJIw6nwYaCcEVPINdM8lOhNJmwYLhFGq1Be2WaVGiwshyIcrDNeBtkk2IzCBB+Q43NQlLMOIw6KsImeMXowxtuAYDYCpOEkh0nrjWDFI2NbD0087DhzDgDTmjyZOm0Duvv8/ySQzSWtHQQGc+4qqrPUL/4bsAcJikYIDeloX/y3c/9JJbqGdeDu1zyJ5UVi6SIbNnP01/Pul0BmWLC8sYVMdBIQ5mwYkG6LD+hmvSwYfvRz169ODI3Rm33ErPP/0alZYgatdr+seWZ+R64mCHRIVEwoavuXPn0uTzL6bvvlnINTN69shjmz1sjx1oxB67cno8nufpp56jWdPuppIiyBZINKAPwoj3R3wC+J619oTFtEWKajrdf8+jClq3kjUSA8gtOw3jgyi6zp3Qp3ZsiTxqZFL6yCdv482emN0Vxz3o0oCokMgkne+aUZFco6IdREW8mfrvDKJTnz0NyLKDBg5dg3caSNsN2Zz3wMVLltDEc86nt954XyTHuIg2gJJolDZ+D+kUSPkce+KBtPnmUkvhk0/n0t/OuIgK8suooFcRZ9U4EMrWQlK9Bo0cBHGPNtUsW0pjJuziNP+5qPZ5lxGt6EoF+SVMwOG6TrZqrx25CDayLyZPnkovPPcKHXPcETR27Chei/O//pomT7qCVuL3vVCUO/r7kaOHeNmra2+mBx940slesRRRvN5G4l6UMjipb+uxlu1fbN43NlL1asU0bh/JspLi3vfRP299gNslxbSjElaZt7FN24JcNGtOSUkGJZqbqU+/Etp7/M6U17MH+1333f8QXXf1TKoG+F0osl9xINHWDXxNEBUopg2iAnf8IjGjwjJbZd4sr13KxbWPPHo8bbSxL6791pvv0tSLb+LMGYDNANPW69+XI/tNii5KVEg/uBAN858VpEnq+lQQPJk/k0sr2OmCa4IDPVswXQ+ow7HW2pV0wEF7sj3G6+eff+Y19dGHWN8AVVGLQ4B05zOkzKdw/RroO3bCUNp8i4352t9//z2de87FtKxmBZNKNlcTp5yeCXi2BfbB/HV7H74yiLGxE3akgZsN4EtxjZSzL6SFPyyl8jJIj0kx7TA5JZzBsNO9+xTSPgeMYBIT17zzjnvp1hn3cx/07FkoWQYhQBc0Oi3pRQAxyAnV0qmn7++A5XfeeZeOPfp0JipQI8fkw8Qqe/vr3HS1wxtsuBqN0zocq7p68X1kX9191z1055330aIff2PiLD+/mCXJcnJ6UNfOWZJVyHUCxKe3l50BGeRqkXOAtC86Gcw8xG28zbukdsenspzHZK+VaGH/P2S/NDWBsBACo76hlnr27Ebjxu9Bu+02lHI1SAG/XrDgB7rk4htp0Y/LOOLf13gKR9+3CPa5vn4ZTYxLPwUZFRGiIvYw1l++RkWMqBh7BJWV96OiIhAVGlSS0CFpax79jb5YY40yOuywPZwc3b33PkgXX3w9lZUh66OEpZcYMOdzS/QGtvZBVIzcQ7IAEfByzsSL6MWX3qPCgnLqZus9+GnE59f35eQjEk2oCYL/Ye/t1AlnCjVEsQZI+K5dIGaY+O3YfFJJGMMvLDLffGMOQjIiQgH1jpB9sVoNvHYaRWpJz7pMDvAeKWcZlp0K5H3ExggYLIG4foZy0CbjFAHK4BeqRMcrwefqIgA8h5S1zmdcE6AsR/Cb7r9mVwghgKwCjfLXLF85w4s6g6wlabOB4cJ+K15ghcYVU2EQns884j864FYxCZZ5Y+wIz6xyYVwbBZkpIEmlLgUIKAS4uFfaHmSBafguP6tmf2gEP4PzirsI7oXgTGQESFaZERBokBE/uKdlxVhWsmUw4XqSUdGZ7RfuZ+MZZg0LriRYj8hfSdAQ+sdk3MLVYnZdCABfN8IyLzBPELiFFzBL+Cc8nsieaWrm5+AaY+p447/IpOBTMMtmSe1QzEXLnBCyQH2goM4G1xRZgYwFL0PFxd5ZGgzB6tJyjDO+wzJbLGPlVTnQJ5ZRgbbhO66f9AwggcRCNrjanK1sNhKQL23GFEM7sb7wnpEThrVBloytgmETBpdqsC+Tb7FzUMx6ydyN4Q+t7S1Metj6Dea/XTc+naVtsQd27UxGYCO1Pv6nERX1yxbTN+8/xyB91fpbtTLU0Y9ampvoq7ef4oyDnPxSqlp3ywSSYSX99t0XtOjrj6is38bUs6xPBhiLLARcZ+WKZqrecHvqCm3F2Ags/mE+LfrqPSpfcyD1KK4g3BvkCoxW3413oE4AHAKrBKP17YcvU+PypdRnkyHUBVqEtJJ+nPchExX5FWtQ9wKRXAiNWacuWZTdPY8X8bJffqDvP32NcgvKqXT1jdgwLfnxG1r8/We8CRf1WZ8KKkWeYemP82nhF+9RVvc8KltzE+qS3Y2W/7aIfv5mDlWsNZCye+S3u1//O19cNaJiFIgK3Sxh0ARECxjxjAMBW/7Yo4hDKYu3Ixsf24RFk042PtvQLKpK/hu9lhEV8l1JVxSnMV60SH7ngA9tUYSQYIMiH0SBZk1tDA7TuBe76E6Xz1+fjRCYXTt8qRRJ3JjzBuEONNEobQe0xgCR8ADkNvw2J4pGpqpjYRFvdji2Dc+u567bClEhfSRAoWVUMOCrv/Ggshh5IyqcDrdmbyUqyGoEBjZv2+ClWLlkP0hkOrfARlEjKPx7/oCq2V6oIeFIAZlHQhYpG6+1GCS6ACC+jUeSTmxsPruv+PdXmahw8zG4dvAnj0mUpcgY9f8oURGsPWsWiAp7+XsHRQtDkJ+/aIdav8BsLIWnsGLremCJWw2/WOVqbq1mGB1Zw1GTHrTVf8Dpx042zByK8Jf6dzCgTD5HbmmOeKYXLGcfA1mT2xkfSNS3CaXiJJojIG1QMNoa4C6ZaWP9dRPuG0YLuoNHrP2RZ44+tFq7SC9bxgiPMqd248AgRMVQJSogUXHR5Evow3c+ofISRG8j+lpJglaIChlPkaMz7U7bF+wztdzusdFncHq32HZjGjp8MAM//44XQJuJZ11EVRWQ7SkQMMGk4MIbhP3XBlHx5Vdf0cUXTqW5n3zJBA6ICmQmYOyX1CymCQeOpkGDt+L7QDbk7jseoGf+9TJndUjWQyz61qatZfpk7Gs+wyNOVEy/ZSY98sBT1LsSgC3AkuyEqP0oiejWm+5pjlTP2PulgxzA5dwPLaZt/ecitfSQisGMgW5mc/4bREV0WL21aysymTq00EFH7kXV1RX/jqnH2Tc3Xj+T3n7jEyopFrA5DvKnnZvswASpQmRrrLlOFY3bZ3fqkZvrimo///QbXFS7e/eeHIjS1NxIo8bsSJuobNXbb7/L2RAFBSU0YMAGdNKfj6DSkmL+/awZd3BGAgDd8Pej9x7ifg/Zqz9D9qqhA0ssWWH4DBK3faayjT5l46tErb+ggS9NzbV07In7OjD2vffep9NPnUS9KyHzU0zZWYjyjWZoZt5QiGzYa96hHQCEuABEAjfSNoMH0E5Dt2IAAAD1ddfcTE89+TLfB6BrVnZ2NOso2NdWlaiwSFJEoC9bvpQKCnPoyGP2cXUd8P49dz9Mjz/yImdMdemaRQM2XKMNoiLb753ajQa4JA3Af4KowH3QF42N9bR4yS/0t3OOot7VVXz7l156mY49+s9U3XsNBvkBYgOkj45d8lSJEhXIJKij7bbfiHYdvh3b1Lq6Wrr2mmn02isfssxWLoqRx+SInMkKEklM2z30qdlGcqQwiqo20bEnjaPKyjL++ZyP59AhB5/AmRtSAwJZVrEaEw7sEDC8uaWBTvrLflRZKTJVKDB94flX87zqxfWBuqUW/m6NqMCZtqIyn/Y/cAQVFMp59Zmnn6OJ50yl3pWo1VEu8m6x2mLxM5OXfrKC4Y101d+voSuvvJafD5k6pt9vezfW0bjxe9LxJxzJGXnovxdeeJGOO+YvVFJSyRJEeT0LmdwTuR/x342ol3Uoc0XOOQKusb+fYAt4XvHArBqYlOnpSRoH+sBlafP9JAIc2AZk1tAnsKkN9bW0fPlSWr9/Pzr1L0dTaalgEGj//fc/RjNnPEQohA1CiLPtIkSrn8u/h6hw+6b6ptwHLMtVSyedsBcNGOCln1BMG0QFsmi6QmoSwQcJr3R1CpmrO+ywIe255xCpldDURDfdNIP+8Y9HuEYFk2rsY6QTFU2N9TQ8kH6CH3nepEvo9dc/ocJC7Dd5Uow8aBv8T1vfFtXPYGcHq4mnAZMszROcOWJJexLPHsT7ZGRRpGxWlv0SBGA522ikAf7LmRRSvwLgMda9kzrW3yK4QAgIKARATgngqsr72PW5cLk8MwJA+aztJI0lqJKzTx1JImcTYDFSHFuAWgbCVW6PfYsOHSRIplnqTQheoJiP1eZQ+TABnOE3oG6nLyYuTRSQGdeTegTwz5tk3bCMeEBaaG09I0YAbvNzkeBCuAdLLiHAgwMCpJ4l/rb6E3x/yIzrnAhtfZrjwL6BYk/4vUgHWmY2AHtfN4NBdPSpBlK5TEIldaRIskhAWf0FfAd9g72pq16bSYuw2Lrt/2yXpKVs1yDl1QUZEcjCaNEaICFu5K0S5ItRSwPPjPUmhIf4Q0xcqdw1CDEO+uIaHS1yO51ntncJWC8KFGg3fBqW5LYAOmsn3x7yS1qUXmt62L4HooUzcloU/NfsE7bhTtJMJZeCPpU9089PlmfC2KCulwaDWCYc26GE5RhiZTYPcN36hkbuRyaCuM6JXNNkq5BVbzgX4wS8xgSfRD8xmadEXabigB87a7/tVa3ORTubK/9vRJ3N2Tiu8buIipA4+f8LUfHrgi/o568+os7Z3am5oZb6bbIjdc7KyQCV62t+pW8+fJG655dSxTpSJDJ81fzyPS345A1+v2ztTalnYWUMMSb66t3ZvOkLKSG6grWLf6LvP3mVuvcqpfJ1NvPgL7IbFswTkmDtgUw0CMIkRMWShV9S6eobU15ZnzS7xe+DqFjw6evUs7QvlfYboNr9K6h+6W/07Ucv8r/7bDSESYnvP36Fapf+QpXrbknd8z0BgjZDQzH+zK3e+L/y4aoRFaNLlnGrsPA44kc3F9fUACARsxVY2+BLbFgYIIMxtSJDAtB5FFB/zQSEsMNpRIVt7FbUJxPEV2jNpQVrY+Kn+gQPPgKIuo1ZskoUggxAZL0PZ5pa+61wszo8StIY8CYbkblC1s7o2rAN3tj6KInT1kTxRIXdKzSYIfkRvs+tzzD6vgMlC8GPEb5qBFScqLB2g7DAy3QprR5EeBvvXKk2pCtC5QsD+43X75LmDEV6AweQMKRcdmL+H5Mq6hDZZgq8UeaZn732ff9fu4PbSbSf/FO0RVSkbWoR+xB0SrixecIlOu7/MaIiWLfhOEk2QtgG6Vf/imVUuEwBneP6XSMPvURXsuPv+yZ6j3CamqvmvhFEDiWtEll1aov0u3bAlUigTKLK8PT4syc6H3F709ZS5YeRaB04daaLaQdyPiDo/I2uTd8n3l2NAmfRdWHZFr5Qujg8wRxupa02gpnjbStH1p1lVIRExZQLp9LH786lirLe1NPVC4BhDWeO/9uZZLe36D0yiA35gvrLbFORin7w0eNpjbX6tafn2/WdJUuX0NVX3ECffzKf9fWtYKtEAwersJ1ExbfffUsTz55Ec+fMo4oyZHmUM4GDGhw4eNbW11JWt0508JETXAFk1py/Zjot+OYnBnsBHBkJzA8R92bDVamfSUYFimn3oVF7+6KuM6bfSo89NJuqq/pRfiuR5f8nvkzk6O8mrI6fAgFGRtveuDK2VzvAJfg9j3ljA2253QDaaedtNfpyOV085XKa84FkVEAyK6lGRdrhgSOm1EjFAarUA0cH4syFjTZdm3bdfTBlZ0mtgH/H68UXX6FLL76BKsv7JMomIQIv7WWEMMCypUsX01HHT6D1VEZHimpfQpUM9hYwgVhaXkDjVLYKQMoN10+jB+9/kkqLKym7Ww4dfNgY2nrrgezL8e/PlqLc4e/H7zvMyV7dfdd9dO1Vt/A4GCHCEXxxRyN5C1jF7hNfXwxC3J9qprr65bTbyEE0aDs5iyxZupT+fsUNXKuDyZacWKZHIgOkRAXfx0sb8bxYSRw9fciRI2nNNfty27/7/ns664zzaOniJpWYyiw+Hh6k4Z+sSkaFWV/4i1gHNcsW08abrEXjJuxOubm5/HFNTQ3NmnEXvfXmJ9Sjex5tstn6NGacgclNFJd+YjvkfFm9Q5jgF5KNSign77Xp87KtjAp7LoAuy5YvodPOPISqqoT8g+zTn08+m6p7Q5ao0mW5RcY8ZT6F69dsR3llLzrgwJEOpH/xxZdpyuTrqKIC6w0EADJtEgJYNKOCiXTLqonpzGIK4Rk2GbgWjRg5mOtT4Mxz+z/vphtvuI2qKldn+881ROISU7axcaRuFCTefAAAIABJREFUM8+Lw47ak/pvIDJYyLQ54dizqDC/wtWKSdbtT19G8MEA2Gy48eq015iduH2416xZt9Nts+6nqorVuSC7ZXIZMcArzDtdDP83NkalnwDSX3ftTTR92j+ZoENtAT4PBOsK+11jUz397ZyTaKutZV3W19fTjTdMpycff5nJCkjTIQK/E/x350MGfW5ArIvuRYADMtZMkz86GcwHZN8hJmmWZt9DH8s9u9VYYhDaPCQAwRqsslKiptFnqGsBKTOQFdsP2ZQOOWScy7CcM+dTOu7Ys6m0tA9LgElml59vIRGIc1R93XI697xYMe2UjIqMs4PLkEJQSR0dfyyICplPJv1UUbE6FRdXUtcu3VJlz9KICgZmmxrp0EOH01ZbbcTXXbx4MZ177hR6990vqKSkmjNHRF7OZ+OGM5TBVkg/Dd+cRo3cwe3pk86fSm+8OZdlqUCMZxA6SlrZaMswrERoWuRMKH6bl0OJQgBRksKNe8SUZc4nOer4gEn242XzjWRb8XNi/nPNB0S6AyQV8B0vgNgSpKfZAgFWgOxeEAg2R5FZC5+DAeEOKMzexUWf87khyKK2uW6yTnbmDetoYsqBZEO7EMkvZ3iRzoINM+lvXJclky1zXJ+FCcKgnyCZFxZ5xrXFtfJST/i+9ZVJTRlQLe+rPD0khJDRAPsRSDmtYBC7A5OY+FzFLyTzIobtZGBEelYzGWIG7BWEBpGAvpaACsEheHxdcJ3MXT4Bc60DKbAdAtQScKZ1mIJr4z3DRTgTQie/b65YKPQV8C1kTOK2sAtWs0Lu7Dvb7o9LcTFzzXIJ65TIHFDZp6BtJjsssUEqL6aZDJzxgLFXEizMqrCDFxMVqpQiNlelt/RamJ+Q6+N+ggyVygrzfCA8V1epe4Lx0/XiMlO0HUwaaAFrm8OY3uibtoiK0M43taxgwsjG2XAqRxRqjQ98zllNiuHi+bgui44xk1aJNXL4bm4eWPBEZiB1YPFMPtOCE82NNR8s+KrZtIxnDtZd3PXBs0TwpP8/EBWYTF+/9xx3HaSNvv/oZcqvXIOK+/bPyKrAd+cj86K5kVbfbJjKJdmpeSV98+ELVLf0V74WJJXK1tw4iFBaSY11y5ioyCvpQ6Vr+M/Q6Yu+/ICWLPyKiQoQEpjIDbU19N3HL1F2Th6Vr7O5k2f6dxAVPP1WrKCvP3iWGpfXMDGRk19EX7//PDXXL6eqDQZJRsb/8y93ytCIk/+PvfeA06uq1odXyiSZZGaSTE0mldBC6J1QRAGpShGkKSLYy1WvKCr6v4qiWBEvikoVEKXYQBBFRFBphtAJvSZAQkiZJNPb93tW2XvtU96ZQSzXz9cfJnnLOfvsvfbaaz3PKlofHQfCQB8N9vfRAOrs9nVzxsxR0zpYH3LaW1WVRK5Ykxt91hQwzU6AbRtrLhtTuSRCR5jj0EAHDZy0VrtsrnTb8UGndROFqQfTq9kMycGkhmMJUZHbzKne0EgoIVKszBeY7dSZcI0FWbnIeEOfDe3rYYrCDugIgsTn8yAQH3CavmmpmWIYOiCyopylRIXYRgLUI5LC30vGBANF5SLn4MWmwJZaKNcTVjwSFfwuj8oMAjxHyMJBVMjYKm7WJbHS8WVEhc2PRUhIKQrfmNjuYYc0mwlq+xlomSTuBkIhsNSuhIgYypD/finnlDFGfUM6Gy2nC4fbxqeoRFRI5FV0PDyRksyEm5TkYEnWxN3TzaKkULsvMtDmTfaC0k/pA8e9ptfxY8NbfRrlkDqomf2ptWF5khJg2c+VrF806izLpbyZdvYuYT2yGmIIIpLL2GnTMsiXpKvG8mW5xMmkOVXUKWXbT0xMeXlCsNJ2NbJM9qikU9vYYj3+uL/CPotCKY4yp7Vqje7MDT1956WC/54A7LaH07rj+uRuj9vPZC1F9SlRse9utP/B0cEsJCpYkTsdUHGCbG/H2Y3jEbWL54PxuMXWm9Bhbz2IJk2axPMIUAulQrhGLBvbMaOqdA31HNlt4S7U0NDA+uzG391E5597ab480giJChAp3z/3h3Tpj35Ks1vn0rTmGZzFIM1uLSKqh9bDxpjdRCe++1hqamrkoT755NN07v9eSD2dAzQZ4M14iSKWesxuIwSAK5XXfyZRYbsi6D4HJts5b0SFyFMujUlLNfhViz0q/l5ERaUMikR+AEh2d9Mx7ziItlQg8aXly+n2227XGtlw/IcOXDFbARG3O+64Pa/vK6tW0VnfPJdeWrZGSgflmmoXA8IhAGCURFyiHv+uu29Jhx1xADuHKOv0PW6q/RxfF8DHfgfsFspWoTzUqZ/4HHV3DnJ0OUqBbL3tpiErg3//3QvpUf59C4NP+P3r99mFHXE03f7C579CTz2xjEF6ZC1wQ/giBy9nd1Q0cEo+VLuggKjAWdPdg6ySGXTMcW+imppJLGM33fRHOvecS6l12myq02bwIdujjKiwqFXWeaYv+9lZ33r7jengN+/FZbNw/euv/y197cz/5ah3RM6jdNuYKkfUZJo9Qt7QLLe49NOm1NIyS4lSi76Paw+AGRkCbevW0H4H7EqHJs21V3Jz7WeeepH2fN0udPzbDy3tUQGiwnS635PGAaV7WDKbi16F02dlGYco/WTXCw2vP/1OmqENr++440769KlncEYFQH5pBp/pI1EiTyl4JWAEMlFOetdhtMOOW/NtV69eTd/59g/p6adWcG+EiSCwuNRv5qJmX1m5Bi5JIesR7yMNpd/1vsO4uTpeOI8+/z9fpqeffEkbaTfw3rJ5DHaDIN78GyvPdMihe9C+b9ydv4v99+1vnUuPPAyiDU3aUf6qYJwVthIDk73d9JajXk977rUDPyMaF3/9q9+muxctoVaU6mHyWrLsJH/B65toTUiPijlJH43zz7uYrrriOmpGLxuUt8r02EG2Fwi2ORu10Ac/fAL30MHrueeepzO+eDZ1d43i8k/jx4PIESBUtl0MimFQC+CplSbmWuY+aCZdN8ivPMfwX74SZ/RfJCo/+Hc59ChG+MOOQ2lokBU9PRvoy2f+N83WDCE866dOPYP6+sYLKYQyeqNiaUCxAaXcB/R4V+cGOv1L7w2ZYbfffid9XIkK9H+oqoqZYQbKi5knNhf0FMBD4DIf/ciRaUbFse8nISpmSgZMyKjwvrjzldhv0vkdhejxfpo1s54+8IG3UFNTA0/www8voXe/+7+ptraFGhshp1I+E4ORJ0vXIhAVSY+KdmKi4q5HqQE9UwqICiMLxRQS304CfdKXyY6BzmLu6b7Vr/oRycdq54qZGx9ZyUp8R7I4XHPsPgFerVSM0Fkc+agNt12Dbo0BlNI3IC5kvQC+cz3/0aN4n6BsJEBp4AHotYEIcPyH8xa2Asr2SOm+QQaF5XZSdoflVKPrw7mlgDXbz1zaaCyTJbEMt8wm7gH/HbJj5eWsxI/0XuhncoMjz112LN7HvpVeF8imkBJG8MOsDDhnS3ApJMELuEQ4B26Npj4EEaqrwKWyuFm4fBYIBk5k0rLc3E8zEguqLfQ8i6sqOlZLUdmaK7EUKl/wvEvpI8wHzhhkFyAbRONYNOtbCB7T/ezHYe20ggPrCPYx1aeyIBgryZ1U2pAdIeMTG1j0i8pXqOgRKwxg+IbtYG7wfdhy7F+7nm9CEin+xo8vGTu8wlryyuxurAM32MY6uWolksHj91M87zj7QHFSkzfYOpK5YVVV5Dkky0JKfvP5prLJJI6WmbJ9A1ng/axZPXwO9WNvQQ7MxzEdJNNmxECwgcO+jllKGK9lC7G7oZlDVs1DSk6N4kwOvIzMsPUsIkj4i0pYWpaGJ0UKTxxbo0wzbbMhvP7i+eXBuitljrKsvvv/IVExSCgXteyh26i2aSY1zd2anrvvjzTApZv21jJLcQIxQWtXPEMrnryXSzfVNc8KG7Cnq5Oeu/f3VF3XxGWaIHTzdj4waWi9bvmztOKZB2jaJjtQXTPSfqNR1N2xgZY+cCuhb8Tsbfbmj1CCacMry2iWkQbBUv7bMyoMWHtm0e/4gMc9Ue7phSV3UMe6V2j6ZjtTTYMQJv/aL5VqdRSUKpZUswKi4i0t7eFxVHWKYqvoCESjBjyoHAhmOOoBIVfRRNziZny2/0JEMf+kzFC26xljHw9nUThQ/tL0SZRJgUXi5EUaS8kTh0hONxMBKOO/wCjoY6Y2Rhr4Mk/WfF4vYFMQdKv9JVw1sPV2Sx4NR/+LiS0stjQtKnNOfI/D4cglStDIy9gdt8h2cJpRxwaQOi76Hp/zCvpKI7D4ezMOxaZ19wl3VGtEPyoGedPrxes7Noqj04WMwRg4dRYGh5bjCvOphqBEkUiPiuwrAvWxvqIYMeow6YHBYw37yeH9PpIn2S/p5kmBf12BMeJQQIcaKx+IOxXN8ExaRsmnzcp+Q0SMPLsB3hZBAOPRyq6xWR/2RbYcmgHKuRjYuBsSZWBaQpvSO5GX7WSECQwXNGWTup8wGGDU2qXEqNI6rBrlEtJPtd8LE2Ga/itZEtqEmp0DXbPMIe7/GVbBInzY+IGRJ4Qs19bkUgNRlrOEVF5o1MjMRjkjJdlqZeYIR3GdeTyBJHIyl7mJEXpIf8b3WT607FESZW97mcUzqzfTi/q5kB1atEd1flU75X4zSJpRsUsJUaGln5ACrWdC0AXy8LKPjPA1D8U5ntbwL/q2cS+BBHjLcQfRjrtsy9d/4cUX6b8/+gl6+slnuCE3ALi09ER+DuBLcBp8Xy+detrH6I1v3Jfl8MWXXqJvnHk2bVjbRQ0oE6NNtb3RHo8PGZNcp5+22ArNtKVHBcZ4/nkX0c+vvJZmz9yIG7YCCGNHU4lTjkrs6aG29WvoDQfsTm86VIBlXO/mm26lH51/BTU1TuN+H3BImKwwsFC3X9b5tzXt7emlzbeam2ZUXHQpXX/tH2j2jI1o6hSpUW86x58bKcgX5244Z0vZb6M+FnkLjoVv2peR/zjnnqjYlvZzGRXfcBkVtSGjYmS2melO02hF5ImdZqibPGvuNDryWOlNgLW64qdX0Zlf/iYD4BMnaumSIexDPBuczW2335JO/fRHqaG+nq/1q19eR1egeXXLLJZl61Nic1Z0fnnZtCbXqIT63g+gBM103me///3NdN65l3O2w5QpU+h9Hz6Oy1YBwL300p/QZZdcRa3T0AR8Ou+fjo719P7/QlbGZvr7P9J537+cWppaafLkyfyZlb269dY/02mf/iJnU6A/B4DKUA+58MSN5G6wEjL6u+RnQ77N4FdvD61bv5be+8GjaetttuDftLW1MVnz+KPLNFsKoLSUvyi7dSrLYsPy+TpqgN5x8ptp400kYxvXxvo/cN9jDEjXT4XeEEIy/xJQAtfp7NxAJ777UFqw5Wb8NUTOn3zih2jO7CxRkV4FNryUhumgNWtX0vEnvDlprr148X30za99n/Z63e500ruOzhEVs1rn0WSUEEL0I2wXFXz+wzZB8ch9ckn4RpinIpnPRLsGPZC5PmcSdGygT37qxEBU3HnHXfSZT3+ZMyoaG5W4K+j5ogpF/siOWxcXviv6M2y97Tx66zFCcGPcf/nLHfStb5xH05pnaaNq6EQz3OVi2T5R7sHlc7Zb+miX3bagQ968N2dm4L1b/ngrnfaZM2hG6zxuRm+ga1aPJnKGUj293TR/C5RvO4SzZfD57357E33vnEu5SX1dHaLxUXVAsgnKAyXiYsI+rqkdTye/93CaPl0qAiCy/l0n/xdnaoBgmFJbz4Fk3GTV1RrPSF9opu0bfl94wSX0y5/fSNOnoeRPvfTRcPKAZ0C2AciiAw9ZSIcfcYDUgR8coBt/B92Cs66VJtXU8RlZRIp5y0YCj2TFo+0stfKtLxAHgnBAR8EuLJRLiXq36F3xaRU85KjzaCvFgDKWACd5AvBBB23Y0EanfPIE2kZ10PLly+lLX/wWvfjiOi5rxGQuypyIFCWDZKKiawOdfvr7EqLiFCMq6ltonCMqzIc1ebQxYZ5Q+umjH3lrhqh4H7W2bkL16AOREIDw0aUfgPX6k1gCsbtZ1hER3d9LJ5xwAO211w78PubsggsupQsvuoqmTZtLU6eAiEGPnqgDxfdQ0FSb/fZ2d9HBGaLijDO+SYsWPU5TG6RUYTajIoOgJvMGYFT6AwhwKnhHkZWkP/P6ztlUvNbqc8vzoSQbri0+gpSAtrND/i6rKPMXmDY8s+p7gxq4JFOvkG7WrwbN2a2vInSJlYnCvfEdKeWDSH55FpAFPd09NEAC5hvZgQ+D/uJgO/hbvTSW+4TIC6QA1+/XCHieJwaeg1OezGmEUKKMChkSI/dxPYwR15gwYTyXQhRSRXohjKsax33g2FsdIxnltp/wfMiuwpMBW7E+FBLIJWSP4B9ChOB3HIQWNL73YYwswDyYnyVnN66BufC6hcFqbmIuL8EvZPck+1L9fgmWteA8+65gRwz0c6krZFaBbBkjzay1vFUkPp39a4B0RkV50JlLOiH4SvtPcBBxKM0upKY0uI7Bo0awWGacNCqXvWhN2PGsku2DRuVS+s18V4SnMkFlmTBaul30i6w7dBeXVhqAvErTcEMPsHbwbRBkZSWjDD/jedayUF71le5SlnkpHR9fut90n4oGzpRcd6QdQLVQaaPA4sMcmlz6bBkeK+ZCg6QNr8D7nPkRCCB5dgvoDWSWlVmvYN/aNUKGtz6kZeqMzJtxM/TvnlGBTbJ62WO0aumjNGOL3Wni5EZa+dxD3EgapZ1q6tG80k8fasn10tOLfsu9GmYs2D2kua1/5UVupN08d2uONHjluSVSPqm+RQ4+NNp+fDG1r1lOc7ZD/wpJY7YXxoJm3iueuo8aZ29BVdU1tOKJe6h+5mb8X2rQaI+K5U9R87ztaHLzLKeApAa2H3co/dQ8m5rnSfMz1Exc++JT/F/15EaaudUefI81LzxBK599mKrGT6Tmjbel6rp6iUL4lyUsdGe8CqLCz3/x4xXV/YRWAOiWJSpMTqBoYvMdvw6mZPSo0D/sqMgDaR64NoXHjv+gXR9rLSomKEI1avnfQXRRR9IfUlmvRL/oRH1Qm1/ZwW6AC2pRilGrx5tL7woRFnzvodSOsuvWjAuR4ZwdIYq2wBXjNMjhgEi2rsMiKvhEEqZe8XmdOsvisMbHyYTGceTKVMjY49PL3149UQHD2UXIWzRCqD3tDjI+wGCqePkLs6FjioCxcDVcYDQCqqGxlIK76ptkYf1IfFVaajcLWpKKIym0Tn+M1pO59QdYiHTRWqgwAiQyRcw2qbAWU26HIipS7kHXpCSEoEzGvAMZQVxxdiyyHeOT9EpJe7YoiixRgWew+qAcYaSRJtYjRYUmUot2w4whkDdpZO/hfzDQQZxYnVJpYoeSbyaTiQbMOZHxUDFC1R9YxftCBpy3VsKclqgFb/Ag+i5GefhIQt2DXA6NpcA/QPL3cBudtzKiIl7HSbj9poSoQC+GhwDWTZtJKWjsxsMDyKW/Bd0ioy82Wc0Za57eQMe943BqaKzn391yy630yY+fRs2N02jqlHqawI2IzUHWjepmgXUBG7/SoHb7HbcKTbVhYF/506vp+mtuopbm6VQLR5lJMrdnw1+lkSEoZRDY87eaR285JpZauejCH9G1v/gtzZ4xj+qnNnJknBED9pwwRtFXYM3aVXT0CYfS3m/Yg/cJyvH88ue/phuv/xP3q0AZKkSpht87pzq72JxR8TcQFf56HkQb7hlTRFbYPjZSgJ9fnYyhG8P+/YiKoucrJSrY0e2hA960By3ccwfWuygrdOaXv0533nEvZyvUTpIm8gLqVD7uIWtY+4+d8i7aRZtqc/PrL32bqH9cLjOhVP+67SUy3celRw457HW0z3578DiZgPvqObRmVQcdePC+dPhbpPzLSy8tp8999ov08vK13AcAjbyrxo+jrs4Ozso49PD9GRTF977Ov2+nAw/ahw4/cn/+PZrinn329+iWm+/gZtWWCSJ2WV6pyfqLDgiqu4ITV6rISj5gl7a/nzo622mTzWfQ2044nGprxad44smn6H+/fQH1do+mKXX1TMhIFm2Z8nXAjNpj3ER9vx3pDfvuFrJIf/vbG+mLX/g6zZyxEQPeUoJsXLlNprWZJaMiJSpOOvFDNHf2ptTcMtNlVOQfVsrM9FJHRztNmDiK3vO+42ijeVKGCgTYjb+7mR568HH64IdPookTJzI4cfFFl9J11/yRZrZa9HxxU/Gy5eBzPk2Q0+AIF0GqQzWwpwxUzN5DSh610ydPfUdCVJz2ma9wfwchKlxzcr2P7FU9U9xKRtmzqFspVbNu3Ro6+b1H0I47bctjR/Ty1VddQ7/59Z+52TyyFcwuMLkoJSr0rAXQN2XqJDrhHYdQ6wz4xsRZRmd86Wv08INPUSuyjKY2KzCdl7dUBwmQhNJe//Wx42mLBUJioSTg1848h1a8tI6zPyagUTsifrkXm0wGl9Mo2XO45oEH70pv2HcXAcdBsF7xM/re/15Ms2ZtQg1Tp1FtbZ1+pnNWaEdIbfSttpmbZFRcdOGl9Ktf3EQzpm9EddpLJNVXku0F0LyrewN95ONvpy23lJ4JyBg5/4eX0b2Ln6CpU5TkK9iX0SP0Ci9LVCBaW+aYy6EM5W6FrSW+xLhxY2ls1Whau2a9EpnWK0PMN7Ot7RyTGvNZaZasT+jgz37uXTRvYyE0n3rqaTr5pI/QVJTwamxlebao3uwOFyKynb6QIypO50yIqUxUmD2RkjFCoojdE4kKNNN2PSqO9USF9CWx30SQU3R1PMekZw+CO3ZfuAUdc8wBNGkSSoETLV26lE499fP04ktt1NQ0m2q1tJWv+2ngtI/W7+EeFbvQ4a700xlnfIsW3f0Y1dcXExVl+sk3opbmy7GET9FxUcKhyq628mKqW8K/XT8t7+t7m9vLAwJYuFSSBRqBKOjt454EAYy2XnfsoojdKueYy2rQjAX0FcCCcNNjRLAjEA3VC9hdlcxxNGS2Ek4cUMkNsaXsFMpsImCPqxho/wcDp2Xc6qcbdKJ8YKhEEN6XDyyTRJowS7YErwP6AlRJ+SbIyxg0v+ZSSNLnwgBwXiPLptDgQIwdZAfE2MpQWa8NmzPWyQV723p1sJ2sdn5c+4gXsFzrsRV8LL2g6S2mQljYYsZDpdI+rH3Zj5QgSiFBEFSAJtNZ/MONqkAQ7T5MUug1OfOE+0EIYROuK4CFEkeyZy34z/r+GWmLZ+WyY65Hl80V5AH/yfU1G0gxGhlP1IG4H2fl9PWFMk4m9xIwKZMrsiU7FmdTFQKxECiovVP8viynEy2LJe/Vix4WW1NkSfQx8+zBX9X+p5pJUXSsseTrnPjnyOp2yeKRYEPeW6H6RCQqeO6V9DPfxje5LtL1dq7Y3PEzFCmtEbw36t+eqBjop2cW38R1C5FBgU3R0baSlj50O02eFvs5+DmDsnlhye2EDIjZW+/FhAMmGwTDupefpznbvp5L+Tx7381UM7WFMxMgGCAqnvrrb2hCzVSaseXC4kiKgX5atuRO6lq3ikaNGUNoiD1rq71oLKe+paJuzbTHjJsQel3gGzX106hpzoLEc7Rm2lXjJtD4iZOpt6eT0+j6eztp3IQamrFgoTb+JiZiXlhyF3Wue4XHje+jDBYIiywBMgJZ+jt+VTf130RUxGid7EBlA+tmUiUsRoknKkQ9yX8AibMZFdmtaNH25g0Vs6hBY7Kza9HVFs1gkc7uJDP9xtrI3TNEIPu39Xfh0I4HoijD2HcDT2dRznF+/DNZIy8dwJAkhaV7ifIFO8uKixlzRBnZfGak3ntSmp5uxlaRgAlRoUaJO/GDmWIHH6PeDvrU6FcBmWMUvLcYIvCaNScL5tURFcUbwZfAcvOq3jLOldh3Qq4QiUv5fnLo5ORP59OtS3T0JPuAZ8ocQBuCM14Shzi3PL40l82HXCTc0uoWsixZkzQBtcMvXBkb23c+lVO3ogD8usXM0GCAX6PCzIAplI3COUhXZaREhckvjFRL6zSQ2G6XJSq8I8j6xX0xrqVMtDmOstDZk6BgR6qzgLmL6Z0CWouxJmXOVJKKt3R41/Z09sYqd+Eqrr65K/EQ7hKer3gHiI0s+yASnhK5IbKX0WcmDNnL6X3Ct/8eRMVXjahAjwrrF6DRZ25v5MYdSgr4ucvMq9VBBVB4wEJ6/X67c8QWgNJvn/W/9Meb/sJ9IJApIESFOe+m1dxyWqQNR3kCFFpP//2p99P8LQQUevTRx+h/Tvsy1U9ponqOPBZAIL2Sn3vpCbH5lsio8DXhL6HrQ/Pqer5O0R7CGNo726lq/Ch69wffHvpVAAQ///s/oieWPMfPxf0qNGVeRL7YZf9nExUlkuyc/yiznrjI/m6kGRU1vi+Ku1glgiVLVIR/F5zVIFvr6ibQ8e98M02bJlHJd9+9mD78gVNo+vQ5nK1QA6IC0WVFeiR5QHGquro7aaddF9Bbj3kzA/8gqC65+Cd0682LqKVZmlfHXg/Dc12ga7u7Oql1VgOdcNIRNHXKFHYor/jpz+nnV/+G/ucLn6Dtd9ia1+O3v/09ffXL35bxN82g2trJfL+e7m6qmhCzMvj3V/ycfnH1DfSJUz9EC/fYifXPI488Sh98/8dpyuRmLquEJvRwRnNNtPXZLeMvC2KWr1HZM8eMwKzccIZTD7Iq1tBRxx5Ae+29ayi3hmyDc86+iGon1RPkhbMKykp1WdCJlnTAPt15twW0/0F70sSJ1XzbZ597jk752Geoo72PWqfPZkA6X7IrM8LXgKhga3dAskfQ22HmrCY66d1Hh/JxAOB/97s/0L77vl6Jih7uUfF3ISoyQEtqJpXBiumcGFHxiZESFX6fJ39XO0vfA52MMx9kyMzZDfSOdx5OjY1Sag+9PS65+Epa9Ncl0heIGx1Lto2AvcUvA9mqJ1bR0ce+kebPR78kAcgvu+wnDL6DpEC5JmRHjc1j4yZ0AAAgAElEQVSUQ8qoAz3KBeRGn5WFe2xFRxwpWXa416JF99BZ3ziP6mobqQbnK/aZZtkJ55snKvA7zO28jafT0ccdQPX1U/i2K1asoM999kv0/LMvc8YHsqAmgAjiyNxyvw93eXVEhdjRaLKLbK35C2bRSScfRbV1tTyeR5Y8Sp//f2dRbU0DjwUlqHKZLc7M8wEWFtACFg1733wlAHLDfVmW0jveeRDNnNlMP77s17Tk4ae5KT0IAQm4ERvdgEMBA4uJCsjAtOmT6T3vfQs1N4uc3XPPvfSB959KM2ZuQg3102j8eCEq5JUG/w2LqBiH0lFFJUBj2ZahiApkdiBr1IiKCO5F30nkCi8AkH00Y2Y9vfPEQ2j27Bn8LiLlL7jgErr44quouWU2NwufMAHnlmUfGNZr5W1iABICQw950250+GFvCD0qkFGBHhUNZT0qhlhU63mJ+0tWRTFfZX5R/nLZgEP18wHyl8hULN2qkqk6EWcLgFkOzjIiQTOWjFSHYHGGQ6+AvgYA4z0ErXCTYfiJSp4AZJbATGSaowSSyCD2Jf7EbwTIlvr6DJpz+W05MzmgU/1OI4+8rRVnS56FdYviAOGcDpUKQHjIuK1km/QdIK50AOCbA4xQ7qkK5IpUijBgGXNvpbTMKYa+sjJRXh7DOmlz9iL710g1K08kQLJocAH9U78Rc87+lQZPeTvEiAqvV82nLRJBlNUWaEDk27IpAjFgwauZH2fBcHyMObSyTMjQM+IJmIQ10cbnmHP0DMqSi7KGMh4Dv0VfRbLGSg8HYkazNCBfgehQX8mauIdyXJq5g4AolH1KSALrf8GkmGRy4HrIMg9ZDwWHaiWiQhoCZV9W0juNAeTnHRS5M3yG51hLL5WqD83yEcI/zhvGJdlOUh1CNKHOcCY4wJ7B404iEtmS43EURnbYO0IUaa9cXy7FDbxIZnKz829NVAwO0obVL9ELS+6klk13oMktszU6rJ+eufsmQur7nO33obHjUN80vjBxq5c9Squef4xat9iNsy5gQDy9+EYaWzWBZm/zOj7klj18O4P+s7bak4mG9jUraNmS22nWlnvSpCnNxSFog4PU0fYKLX3oNt6Q0zbbkeqaYraEGwU301770lM0AcZO9aTw0YS6Rpo6baM8UfHInfwdjH/02CqaNLmRJkxu4H4ZY6uQXhsdJTTOXr3scWp7+Xnq7epgYaprmUMNs+ZT1XhxXP51XiMlKqSZdk7YS8F1rzhsjmT7pkCUbWmA3iVEBV/K9YEISrbk+6qV0UfAQDxcgQ8RLWtkY2DFkYREaYqAPWgS+e+fI85EmgcgkbgGknJ6/6A0kTbHxhQ/p4KZAZoFCkvinqXpuADu8ndhp60pU5HJxf0U9OUP2jJlVkpUaASozKlFoyhRkaQVBjXtVLYMYCiiIijwDF8cxcwDEyVEhezYYNybDEhvDSF3OG3bNVITh9PLU3ofGbvJoZEJBvIrI+8YehFXF15o200vm24bH2WfqjjjPCQiRtI7bWcZ5hyAao0+CQRAaHwl6a5GVMj3Ef0rxjHIJjPgguEnSi+z74IUjUgXyErY+utfBn1GRYw8sFqTnnQwo0gc5Gh02HoIXiAfmOFlw/eGsx90kXaya5ixIVElNuOxgaPtsUgmFYFlVl+/gKiIbEA6j5VCuErwODO22BDkurjqvGjtz6AP9PdlzQ/NCYhDk795hz+uvqWJm0uRLi4eo6e3m/bcJy399PWvfpMeRkbF9NlatqZK0mNDknbJ3g5p83IfXWUVqLgvuQQeDdC7PnQczZ6DEpFES5Y8Qh9830do6uQmbuI9uS4bzVxOVLDeZvCqg95wwEKONIfxD/Lj/B9eRIvveoizNKT5LvZmej6Ef3MjVRAVc+mIoz1RcSn95pqbaNaMuUnz6kQvq46SKNp1+X4VTz1N3zv7AurtGqTJdVMlClz7VbyWREWiu53UZoH8QsXg3iwDnM1BMhDMnKZK1/tHExVSksuCBdINibmGPt1tj63ojQfuyVHXIBXQRPa6X/2eo+kbG1sY5OTMMeXJyre81JGG8zahejS9+/1Spgmv0Px6+hypG48eJYWAVPHsCWjRw1HZJ77rCNphR8kWBgF32aVX0SdO/S8mLxDJ/PWvn02L//oQtU6fQw31zVwGBPdCFCRKl7zp8L1DVsajjz3Ojd5P+9zHucY8HN1LLrmcfnzpz2hmKwBZ36i6uOSKRebx6ZnT9UXPM3KiAmtlpZE6OtfRhz56Qmgsjrm5//6H6MeX/II62/u5lwTASAY3XekC00PmgPf19tDCPVF2bCFNrBZbf9369fSdb3+Xbvr9X3j+mhuny/UqZVPIRmM7pTij4sM0d86m3FwYWVS5ngzJFAnZhd4I69e30XY7bkbHve3w0FwbOsXKZUAeEPV+/bW30MwZyKho5HIcZfs1uxJQ0QJYpRaod9750cJRoU59pTPP3SQQFZ96R9gHKP00ZEaF3S8cXqN8y6zEysTZiHNr3YY22nnXLejY4w5lchAvkBU/u+rXdMsfF7OeRekuKVUp0dD+qU2XwR+cWl9DR751X9pkU0TNi52HcX/q1M9TzaR6LuE2ZUqjI8/L5DlOBo+zp5u6e9rp3e87irbZdgF/CJDo9zfeQheedxVNRfbHJCkJGMvRqE2qp6j0S+ij+oYaOuHEN9HMWaJfQLhddulP6PzzfsLl2kCkTBg/ifeB6eVyuXj1RIU8AzJbuplEPPZtB9A+++6h5Zb66OdXX0s/v/r33DAcmS1M+DpD2tuZZnB660tK0Wg5UOuRMvR0s8WBce22cAEdetheXCptw4Z2uuZXv6dfX3sLk8UgTrAX8Z+Un/G9BOMoTF/09nbR8W8/gPbYYwctczNAl19+Jf3g+5dTa+s8Xj/04zB7mPWN2ytGVHz+C2mPilNOcRkVICqCDet3rPWjFFuqp7uTPpIr/fR+moEG6g2tVF0tDd5Tf1Gb5cIPZLdJiL6NN55Ob387yJxpImWDg3TbbXfQKaf8P6qunso9L2pq66mKsz0sS8NHYss4sa64Xk9PJ73pkN2SjAr0qLjrrkeoqXk2TZoEgg9ladxClugU6W0gpYHwMqC81E7SLPycrmPgX8gJ2+vcb0F7KhSdUmmPOS8PMcjIrgdwF2dNyKbRDAkA/rgvglE8iMw9BLSRMaYBWAA+5+dESWMA+wCLNZrc+p4YQcEZFdzTQUsMczlgIfHYHrMeIjps88f481BMVgFaBX9tjg1Q5YbE8Ec5Ej/2FMD7ANq7u1G6ClkXIFLENoA9hTGijBVnJSPzYszYUP5JMi0keAwYh5GCPL4K+5pLa3HPy7Qnw+gx8iPr34nn5jJI2pvAkyf87FqxwWzWMF8lmJj1/ww6FIC/lvjMkmWpn58H4VmPjR7NJbFwRtn88rppxL6RF0wI6nverzYyy4K2OPBSS3ZzRo2SbizjShjx2EOWgJCzliESyC8OiBQshcc1Nqs7fEZSxD5wT7YXlDzM7bvykAAMomDbyR7CegohqQQRy1fKTto+Ltq7qpFkDjUrwzAXK38V8R6pcMHrx2VAUxyIMT8uzWU4VMSQyh7P+rvaM5h+1A2aG/LQz6JP9O9MVEBIX3z0LiYGpm+2I40dL6l9eLW9vJTWvvgkZxLUz9w0nUDU1uxYR8/eezNNmb4xNc/bihtoL33wT9S6BcpFtfJp9fKzD3Fz7Nlb70nja6Zy7wc0x95oxzeWHLqiLrH4T9x+LW+KeTsfxNke+VfsUdG88XY0ucWTGZYiGzWclX5CzwlkjAz09dKMLXeniXVNJVkSAgiiPuPqZU/Q6hee4CHUNs+i6ZvskGsyXr4p/hGf/OOJCqnpydvMuyz6XozOj09fABYHg4TjDQqVkyhcRUehNDQdc1AjBVKw3jMCHkW2vweIVUduAJ49iRujOmm4HQ5cS3s0u0nuG1OxRXIdiDuMZVcaJACzkkoIEFpSN4ciKrySKyIq+Gl8RgUPUtbLnkOMMgFGLYPElLisbuq4+TFFkgZppv6B7R7GSMcP5TfpOoTZj2hxMnvRaJG3Y98GZdJh4GjjKD2FpRl79qVkV3jbGSF8aDPRZXh+Cu56oDI4Tl5cCmzrLCHDa+SabPnnlnRBmTcBdYwkQ+mk0SH6TconimFjjxgyKhAhx8+g99EHzZpGqd1XbAWWgpAlRIXNqYF/TB9ZnVodKJ4rJSo0Ki5EdUQyhQ0oa2qsfS1eDVGRGGVab1MIEFeWwQMyhYZpiX5KkJxMiSNPilZegCCOHM2jjfx461qUVRlRUWrsRc0sii6V5WQPo0Yxf+lVEhXTUO87n1ER94vMS1y7NGo1cSyVdMNI4Mhtt/MCOviw/WjC+PFsJP/o4kvp8kuvpFmtG3E/hzypUEZUyHxwTf+eLpraUEsnvufY0OTzL3+5jc762vdoBpMfUzVKXKIfgzi4JquvlqgwHSOAIwCctbTwddvTkUcfGmqd37P4Pjr3OxdRbc1Uqq2pk/rfGVDVqzXMX1Hpp4su0gyP1o24sbfvUZFoag8OOVCA10v3X2hW7jL4hjreikiPojMq6I2wR8pLP339q2fRQ/c/QTOmzZFsAICvQw1EP7dTx/SBEcUDqMcdbBknJ909dNL7j6BNNpESO8888yx94uOnUX/PaGptncukwvgJRipEcrVoOBJgZWWa1tPBh+4VCAEQCN8953x6fMlSLnljTX59wER6zfSJWTNpVPY2229CR75VyDMQcHfffS/tuddCPj8WL76XPvLhT3EmxLQWKdfGGQaoyc0NmztoxqzGkJWB3//5z7dzlD6cqxdffIk+e9rp9MrL62jG9DlctgV112M2U8FxGwA+3kkjtI7S61WWnUHq7euh9vb1NL56FL3vg28LmUq4yosvLadrf/k7umfRIwz4ItspZCuFgARxgFtnNNL+B+5Om24+N/SdQA3uH118GV16yVXcfwDZNOhRYtlX5Ws1PKIC2S3VE4ciKkRHC6jZSW1rV9MbD9qdDjviwFBz2mYMRMWFF1xKv/n1a0xUaDCOSaC3ETggoIyoyJypMaPihBERFYlEWDCQZZFH6ylYPZDrrp4uamtbTfsfuBsddjgyFiQzH8DP7bf9lX5+9e+ot2cUkxUgJBn4Cz6GlH7Adfbee3vaZ9/dqLZOSotBHh977HH67GdOp7a1XdyYnpt0c4aG1AAveqX+ingMONtAZM2a00DvPPlIamySqHzM0+K776eLLrya+npHM7HIIHoGsGawDuflDpvRwYfsRU3N0vAYY0RT5k+f+nnOXgCwjMxB6E000Y3Ek9+bftR/G1Fh8oqMkUmTRtMHPnw8zZk7m2+wcuVK+s63L6Dnn1tJkxEwaI21VaMXERUa1SXPpjXzQ1a1lmUsnfjwATI9+uj4499IO++yZdBfmKsXX1hO119/C/3p1ntYt3HjaTSIHpSeYV6Mua8DotfHjqLDDn8dve51OzKRhNfSpcvo05/6PK1YsZ57ONTW4vwFURgrAvi04OEQFePHVSvmUHDiKdheRlQcc8x7pYTUVGQ/TAxlemxKBLATMBt/VlWNoYMOWkj77bdryCbDZyC/Tznlc7RmTSc30J7CpbuQmePJhbxvx2Vs+vqEqHjTwiSj4ktf+gbdccfDTFRMREZhtsR2iU5hoJLLoam7g/2i2QtJKWjTBqVERQTlJdNGwAZeKysBnBEqPouSoGl7Zu3r0S8kBLIKhKSRJsMs0wiuQ7aF+vrmc1pVBfiB3LMCvUXVheVsCoC03DdJMzZGSc8LXBfkBpeL1qbKnnQZO06IDhkHsi3U3vf2lgZjhghxVQemq9h26ZWej1Xj0GvGCA8tWaUAN4BeNAbv7ukJPmt/n/aW5GwiIcQkM6CH9w9sKO5jqMSvnPMR8Baf2RvicTHkOQVABzEhmSToAylZHtzbgktpZ/CIBKzQ0ndM0kn5J7O3y6P+WUKCSRNKEPmADG9LmwxmCEq///As8Amsf0TwFTTzgTNm4A8qOWf3lGvIgolfa5VAYo8ZKcOsJJqC8yGTQMF2rAmfB9r/U84PaYRuDagjJhFJgvDsWsGAy0OBkKoSObE5zevlstnlhoKZr4vOk+wdyUDwczdmjAVKyFQYuF9mM7K9phV+2B9wJCXfR3WhZQrLfhfMRfax0xmMDUaigudNs3KLziIjWCy7Ds/EZF8OFwpPWGpWJT7WvzNR0dvdQc8/cCv1dXdpg9FYQoEXe2CAyzTN2nrPHFmAz1DaCZEm6Dex8umHqH3tCtpox/1oDAy1QWLy4vkH/0QNs+dTbdMsWvrAn2jilCaavumOFYF+XPvxO67h68zb6cAhiYqWjbenydOkNmTZK/SoaJlDU6dvTC88chc3mp65YCGNr5lcCArLtYSwaF+7nF567G7ezBvtuD+XpPrXeenGHnbpp/WFQ49GdJH7H0Eg/l5Q9v679nfpKZCGOIlCjWZMSgrEWps2NPncGirZBg/GHhMbEuniXz4yk+/IOlx7EnhgOij4gE2n11ILyJo3c/MkKGPtEWDOqTHq8myOdQ2PMTSUYpHRUovSP1P+t5FFH/q68oh+HeTA5sZgOlGRqNB6fHaoc88AK0UjekGi0+N94xwUHSyZ8SXOqvu+vR/AzOxzRYgJa8CHp0Y68QHKhgUOWW3ozEIjALg8q5cOq5Wt86AfxSA6i5zX7A4ryZQB/kUr+Klwc5JblviGyLBF7alf76J5shuG+3sHkF+iE5BebD0fYukniXrgHhXiwbHg2/csiiIZcjBqirXYqyEqpJmX7BGLoGXw3c2zJypEpixdVLIygohFRtDUcDwzMuLm/xlm24AMNSgtckT2BAQ7GjslQTMZvZKVcZnNIL7a88IELjpLrmxJIKpKTo6MY8RTELgzry/17yUqIOiIjA56dRkVg5pRsWvSTBsZFehRMRM9KlCGB454Fjbm8aVERcgI0/W1KC5zJjBv0DO9Pd103DsPp620OSWaaJ/2qf9Hq1a20UwGSmOZpjiblYkK6EKUe9zQvoGOOv4QWrjHLqzTUWP8rG+eQy8tfYWaGlqkPjo7wXF9oTPNeQBRsdmCuZnST0NnVCSOXz9K9nTR2rZVdPTb30yvc/0qfvGza+l3191KjQ3NNImjTdGUu6RRaAlRccEFF9Ovrr6eprvMk8Tw1qXJn2MymxYRhfMXoBaPQbO6KgKzuhivNVGBNfvqV75J9y56WIB2a7w5zGNQtr3MIZx+gEoSWe97bYmTgXNl8wVz6bC37Mt1uaGjrrry53TuORdxc/LmFqmnXQUgQtAM1VFFOiLit1z+qasjKdOEebrxxpvp/O9frs1zp+Sa06baIv/AUv6om7p6NnBGwbx5YgtL+QNxgH/w/Qvoumtvopkz5nIpEoCeiM4zgABA/4b29XTM2w6k3XbbUdL30SBRS9Fcf/1v6Wtnfod7U/D8oxGuAiVl+LScd1FPln2vRBu6t8tLP8lZLDY6ItPXt7dRfcNEOvHktzJZEfbc4CAtW/Yi3bP4IVq86CFa/cq6EMWNce6w05a07Q7zafPN53HNbHuhJNsF519MP7vqWs4iwX9cMohLqFjJoPInMOcfQHS+mfaHac6cTbkM19AZFSZiArR2drRTZ/d6es8HjqVtt9sqPCemG5k7aHgMomLWjI1pcmEfAXcoFww/lD1IxM1ssXCwhF8aiFE0E1l9YUTFKZ96lURFONvFYmLb3NulSqhKtK001l679hU6+E170ZsPO4BJYXt1dnbSQw8+SosXPUz3LF7CJZsMkGiZ3shg9jbbbk7TW1H+TSYDz3r3osX01TPPojWr26mpqZVJCsmwyTfoTubE8C0+20VfMIHe20PtG9po+52QKXNYyJTB5+3t7XT/fUvo7kUP0YP3Px7GiPFMmVJL2263Oe2829Y0Z05r6NfERMqjj9FnPn06rWsDkTKLyUWcJ9B5Flks2eHFZwt2VuXST3NLelTEJ8Y4hERcR7suXEDHvQ2ZLdU8h3+9624688vnUlOjlMsCiRT9O26J6y4kekSCqABAClhm+peBSQWYKuuTSAy9+fA9ad99FlK1lnaztUXGzZKHn6T773uUHn74aVrX1q4R5NKnCq85c1tZNnbeZWtqaECJLZENREX/8AcX0k9/eg21oAJDA8hnOcN9NvxwiIpPaEZFPXpUjENGRlHpJw1o0j5cyKj4r0xGxZFHvpNamucIsTB+ouiK4NupTA8M0o47zaftd9iCttlmM5o8GYRclPcHHniQTjvti/TKK+u5OTiyRKqrJcsHQT9et1v9d4vilga7UqLwkDftSocfto+WfkID8a/Tn/9yLzU0gKytlTPZ25EVyE8OrNMgJ4w17N1RAsymr7IzRNZTbhOz0XlfWu15Fj25Hvs1+r4/7c1ukIbpgp35zHD822wqnhfrodfXx6Au9C3IRgOq0dvB7DXcE9gACPPRXGJLwHgZT5RJBFxYCSj5UEB3NLiGbwi7FRkNcdzRD058r+zMGeCMS7rGyHYdqwyB+YJtJX0JUc5anBcDyblMEsbT08MERXdXtzQ11gbkBjBj4L4kDpfBKgjKCkA4ghcVA2BygudeSCHY8YzNaMnf0C8hY6ohE9zuH/RKgP8LNAqXBlJQ3QKsHMCexKkFX8foBL2ewXbInudsAVlTyRyQCgnce0cFD89oZcUEn1UHUZ1tk3nLyBAZFrlLQHv9vnlLRoLIPnCl5LjE1xg+A3BtqeIg9nHImFAQItwDHIBWu7DnKTLRiy1l24PFRAVn6HJwcNRLMjfaVN2VbTKbsIwOibhdSlSYTOF5rDF4IBK0j6llK3nyR5YoVoIo61NhZZxNB4t/jwDFAhkzMalA1tqv/m17VEAgN6x6kV589K/UOGdLaZqdsQtWPvMgdXe0cammPJg/SGtefIZWPvsANW20La154XHu5dA6f5ekUcmzi29kUKhx9nx66Yl7qGWT7aiuCSWmyj3Mvy9RMZdaNt6aNqxaTssfX0xVE2v4+ZhcqYRYDQ7S8w/8mbo2rObSVhNqpbnnv8ZrZETF4c1r+XAQ3EwYypR99GtjYE086I2oEBAy/a7MBy5crGzM+El+x/6PZWGkDWqNPZWxuoM1Q1SIjvCOVIBH1eDyHkK8VjJK/YfcxwH3hrpaGlj4UebZ1QCUKUjB+ErK2pSpj5K3AwvrI3UKXVTyMIQuPAOvgx1JatgbYcRzKp+ryxTnyv6mc24Ot4Y3ZMaTbbBowI0bqHMu+V5834JZUQJMHBD/oEIi4D85JH2qrtbmRNSGikC/zn/qwDqZcBHSfBctIxYUv4v/9KOwK9ishu/nHHpnoJkBkCuVxhMRsgy8TmSRg/GkRpcdrNY4WAwVuXtI99QokqKZ9XKeSG0ZAGrzFwx0+VVqNMb5DJEGSYm2tBavyLBqCFdnGQaQBC1Y9EsqN7Kk0QhIybIMF6U/zWqCsAMsqi1Z1OKzKB4H+Lw44ytcJpufzJf0jo/plHTzJkeO7gkvBxJQlK+drZxHoSawtU5FMkaCyI/U8cpEk2fPQClZg9JPu9L+h0i5JAAnsfTTrFD6Kb9n9T7Bo8kkirlKfVYXGinYcCZmb9RKRx3/Jpo8uY5Hiyban/30F2hW61ya1jIjNL4uAs3TYzwtxcY1/bs7aZP5s+mYt7+Famtq2OH41S9/TVf++Jc0vVlAk2xJF59RNZKMCgP84oxHDQPAsaNjA7WjZM1/n0wLtOEogJIfX3IVg/JoeGz9KopsJugBgFzzt9yIjjj6QI6mx3twauFUiNPlNl6hxJS/+fijT9El511FkxCJPh4lMeBYphFNRb8uItRTGyP9lQ8w4Gfq7qKFe29H+x24V2hk3NnVqUfZ3/ZMjz3yFF38wysZtBuHZ4Lzz3pLxoT5POyofWiHnbbivQewGiTJ/fc8ymWfuFn6hGqNuB9Oo+gIhqBBN8o0nXDyEbSjlmlC8+uvn3kOta/vpQaUCUF/ktFFWcTF6yQRj73U3rGB3vDGneigg6UGuL2eevpp+sTHP0uD/VVcqg1AO5d+0b0vTh1q5XfQpvNn0bFvezPvC3u1tbXRV77yDbr/nsf4+THGCdUTpQxNeTnegsFW8MacTsr/MH+OxO9oBqJmljBZsaGNBqiHQVGQkbGUZvwVbCqONEUPuvF5khUy+Nzzz9O3v3UOLV70AJeoaWqczn05hMhM94FssWIdz6WfutBM+zBasKX0xnnyyafo5BOt9NNMmlQ9Sfpn6HUEbDEdHfevBZBxr5v29TRh4mh6zwePTzJIJKPiErpeiQouKVbSM6ds5xeR2vLdojUsfm67dhYsqFT6aTZq+qOZ9nhtpu0MrqzJFsYe7PYikZMyI+hXAVJ4h502p2OOOzxk02W0EJctwRxj//g9ZN+DfF17zfX0nbN/wOAxSL/6qU1UM2lyKNVnuozteRddmfhZDrzCnEppnC7Osttq67l0/NuPoKbmptwDQS4A9OGF640blymVo0TKokUgAc6iNWvamVyrn9rCEevj0DuDe11Ee67Y+hGvoIyo+OUvfs/NtCejTw2y/oKsxqvJuktULeZt3brV9L4PHkO77Lo9fx9lzC750ZV0801/1WwUBaqtLJ97ermWZSQAIIwEcbQpi2w0C7CK0ojIckT3YzxzN2qmE044gjbdbF4gebKTjvm2Br/4DBkHRVkzOLfRGwbP1NQ0g7MO6uqkjw/sLYkIBqCOaOM4Vly7vWMdnX76+2mWluxCJownKqq49FMklmPEX/REJFOzgz7y0WNCM23sta6u7ggWm4MUHlL0Jwjpouw4kNw33HAjoen12LHVNHVqCxMeEyfCRtJyaVkbUm1Ls30Ea4BN0pk00+b3ujqdq+wCQ8oUU8n7N998F11y2W9YzwlhoVHkGkBo5WtiVov3i0WvZW1qjI+j/UdhzZFtJWWUBDyO5ZwsgIWBVFdmh7MgNApc+vbJGQFilc8LJd7Yu+AyZjs27jEAACAASURBVGLnSxZA6ixx8A7KJY2F7MnZLiWh9Dp2PXV0zGdA/X4uI6sBlghMhG0B21Ne6e7nDEsl/DB+H7kv/ndcgDhGIRJ8qSf+GpdCkufC/XBt2I/Y9xLYJKcJ7jEWfTZ0XnAPH+WOs1aur+Ws1Pe3EtwyVRZMKT6zQEEyWK7CgeBMEClVYyU7RPEkBqb7B6hqPDJPUG5W/m2ZCyA68H2Mh9dytJAo/HeMC/dyhAhnA+ha+j4jIIu4Ty/7uBpUqRVCQFCF8t/6LAyOj5Wyc0w2hABZeR4JYouLwcuuOBXLYeh1KN/LBg4ZnhNIByWgIllkGQwiH/Z7fN+yJfAefHfZI9HP8kQC6zkdJq+jBsBnS6sZrsNzq6XOUkICfUAw7/F6URJF/iDzrMMsq0LJ26zKyM5FOBk0MtDkz+Yo9oh0sm+ommGDLGgR3PB+X05luSxQ+4x1gcoNruMzVfz8p2PVHYy1/r+bUdFEM7fcvUStYyL6aemDf6berg2SIZCtDUhEa5c/Qy8/dT/Vz9qcGmfNzwD5g9TduYGef+BPNHZ0FfX1dlPD3AU0dfq8SEIMDtKqpY/RqqWP0vhJk6m7fS1ttNMB2uOhzDwSJnTkGRWSUpp/yX1iRoU0CIcwtK14ll5++gGaVD+Npm2yg6R5KlvNgKB4+LpRB+j5+/9M3e1raO6O+9O4CbFMVsmN/4FvqyYYZkbFUa2SUWHR+74Op4q+KHjehDAIzdF2jdeg+AsauoWHLqUI+VhJCY4ApqcQqymvCI57meGOEDrOuN1lU8d1C8+QYceN9Ih3zMqjsfgZMkYQZH3F3whDqrIStUmUgTISLHdbdSAG0GAJhqAw2sZgl4E9RcoXt5Sa8fKUMXpWgGF537y8CKaYDJhhZWA6K88AcKoTzc+VJyosUjPKQ3S6xeFM11o2WTqvKTAXD1s7hM1xCePlXg19HOlp6Yop+G+T7TOC9MZFwUoFO9j5zYnL7pdXDm3ZP9bQKwIPTvbZmEp7c/jrMFHhMipEql1tdfXcRTZiuagixWNT68XNE3/Z31hqqOkBbzRYizT5DM/ggUtRmdaEXRyAcoAKv8f4YdDG/R6Rhyg13uF0+64EOsk+T/hF2KP+yrads0a7v0r2GTIbl/Wkfy8rr2nUVpg70WC8h4KxGUCvuB+CQ+JSW4uAa7+N8s+cl4Js2ZtSomLf3ZKMim987Sx6+P7HqLVlJtWheWiILi+YeTuemI2K8p7LpuBtOUi93b100OFvoIV77cQGOsrQnP3tc+jWm29jogLAEIP3oTlles9KRIUB+wCEPvTxk2j+fAEO0Sj3a2ecRdQ/lqZOaQxlXZwCD+YAHJfN0KPimIOpesIE1s8oDXPDtX/g+v1T6qTUEhu62qwtrKQ7IzAWaZC7nvtVvONdx4QGuUuXLaOzv/4D6VeB0hHoXeBSnuMRI9dAc28jKor2/6t97/77HqSzv/FDakTEcI1EUHKvJufiis9UvseTXZT7XtSoFnEaiIrXb0f7HSBExWv5uu++B+msr/1AngkNsdlpjjq0qWUKvfX4g6ihYSrf9u7F99BHPvhJziZA6aSaWt+bwM7B8so3drDxPIEQ6OygbXfclN5y1EGhJvGVV/6CbrjuT9TSNJ0mTkRzUinrMNwXR6x2d9KUhol00ruPCkAszp0rrriKfnDuJTR75sYMWtbU1Gnkary67AuAiWvpAx85nhYskH2B12233U4f/9hpBBAZGTooG8UlycpsmtygnUOtvbGKn6vsecszKpLzElGpCoqCrFizZiVtv9MWdOjhB9Imm8wLcltpTjEPyLD65S+vpcsuuZLGjh3P5XLq65uorhZNiKWfgZx7GftPL5zdC0JUdNA733MYLVggZXSffOopevdJH6U5szZhAgQlv4wADA692yvh/FUwB3gI6v/jOdEw+uT3QHcIsC09Ki6j31x3C81snUeT6+qJS8cUrFdZxCGuU7yjh7fPo37KRJFqSSNkmHziUydS6wypf3/XnX+lz532VZo1c2NCBDlK77CecQZXUa1yH+9SLD1yDoOswL5rW7eaRo/pp7ccdSDtudduVFcnRPhQL+j4++5DGabL6L57H+JyRWimPqWunqon1vB+ED2V1uk24IttVgbMIsDkZ1IAMylVtW7dGqLRPXT82w6lPfbcLfTWGGqMJruX/OhyuvzHP+NzrLFhGvfNmDRR+rNYVH6whB3AlL8+dEIvbbXNXDr2eNFVmAeA8df88g80fdpcLoFWpgtMtuTZoPfaafrMKfSe9x0T9BPKJJ355e9Sd+coquMSSdKXyXkmblgasMH7Ir/axeWDY2R8lEnJtOnq7KANG9ZS27pVtN32m9MxxxxGm8/fJJQHG2q+7XPMycMPL6Hvffd8uve+JVQ/pZnqG6ZRXQ3ObRDhyN4TcJMbEWvJGtthsH07Otro9C9+gGbOlN4id9xxF33yk1+i6dPncSZMEVEh/nfMmDei4qMfPZa23mbz4Q6/8Ht4pnvuuY/OO+9HdPfdD1BtbT0TFPgTukr6UrCHmFuLIg3B50tPFx18MDIqUiL9bxqo/vi6626i7517BdVNbgyNy0V/CAAoFREk2pvtzpJSUOGsDj0crYF07FPC1rqCish8wAvnL2cYKpmB/c7R6D3o11DFn2NejLSJGRraSFej17GGTKCbfKuY8x5iJ8BhMDzzsWRP1l4Qf0ImCLoHeA+PV6sQ6CeSYB7uN4q/g+8z0aLkAPu0Rb0DbPmda4FhWpkpzrIYiybjIHFi+SGr0c86E33fuEm0PYtE8oc6/tbIXiVNyrEJwSFZ/AbVaQNpHI7skkqkPROzTBTi+Xv5XEHwgpFXGAPeFzJF5slsTstq4B4oSjRirvBd7sMB2eKyTMhsEUxN+oTEEkWYR/Q4g3xwlg5wGe21gFEKKWKljgVX84EKuDA3HB9wmSpKrPEamp1gulwZt3B0KlEBGTJiwnwJszUgp+Z/m19lJcMMsLfP8W+cp6LLREasibYMx2kA/auRSlJaSubXf0+yJSRrg0k0LKGWdpPMJuv/oEiWbxaubSpE0MVw4f1dZsEU2FX+bODLJMFYkmVifSoY21C94gmmkRIVwR5TFc7zq9c22c8Hked9LcZ//q8SFdW1U6ll0510/p3gjBpF48ZPpM71q2npQ3+myS0bUfO8bQqNWJAPz957EyvDjXbaPxdxAMNq6UN/4RJPmKy5O+ynTa2jddm1YS0tffAv3OsBhABKLRUZGf6wGglRsXb5U9SEjJCGGZlnBQM3hpt4435ZooIV98AAvfzUg9S24hlqnLOA6mdsykPDeOuaZtLEKS00BrXWBgapc90rnIGBzBKUwpIa5/8qL0OC1CmQ8GRR4qh12N/H8z/Q1039vV105PS2WD8OyoGBB6yZK4fiDZAMUeHZ01c3A1miAudv1jRVAEDrxbqjFAleBT0t8gZTlLOYTWHkSiAqtClP0XOI4Rs9a4M2RQHG+wXIM4BQXlFH0LXoHnkwQq4mAFdsIMRR53zIDeEommHC0Rpi3MhzyHjlfj5C2+Y9Xhd18oWcsBFboyV57vi+3cz9lj+MPTDiM0dAhw+z0owbx53oteQa6XNHkF32MTf3QrmK3l4aP24c9fb3hmflqZDTJ9Ns3a1IkfhkFixMh06AZXpm50PGJnNlREU8ODNEhWZUhEe0CGg98M35skPNExVi28ReELL7y+EF79pF0KLEvbdoFH04+77IkzOAwz5QI9GkLExKsctpRjLGbNkx+HskTXXyw3Xk+jKzYccNqX6c/ay3lN8mJGuKdiXfCx8VButl9kKGqBAdbDVPVYqdUckiqU+AWvkxoyRdE08oJUTVkE/vFqoAeMqSTHw59wwYBfYW9tJe++5K+x0oDmZ7Rzt951vfpYfue4SBVQZ7x2bK4ISxRWJXDFNpVCgEsvbG4dua3hikuqk19LaTj6CWFgHeUBv5Ix86hSbX1tP05laqrZmifSSKS1ZkiQo/TVh3GIEATfZ+4250wMH7sNMCR+KnP76abrtlETcaRnkKA+RNVkWHSGNAZDAchgwGBW8uv+wKuuHXN1Nryyyqq40ZGSyzToazYwnRpuvX0rY7bUHHHC8NcvE7NAK+6Ac/pUnVtQyQso7LADQCwvXR/K3m0mFvlfG8lq/Fi++jb3zlHM40mWy9LnT9spojC7wVjSNPaERb0c4NI3B233s72mf/PV5zogL9Gr52xjlcwsh6kjBhxynkA/S6fXeivfbeWaL/errpgvN+RNdd83tqnTaHGhtaaDyyCZKG67JvytK97fwS4kqiiydUj6GT3/vWUKP/8cefpDPPOIdlvGYSer6MhAgQfSZlzdbRIYe9LvTAQMk01NFftXI995aQ8h/53hJ+X+y6+5Z06OFv5Chb3utnn0u33nwnN+NFiRuUjSqSxcpy56Wj+Mwpg8aLzv+ye0HFMGnT0817HIQkgMiN5s2k/fZ/PW251XwmA1FL2/YlIqbRLPuxRx+nP9x0C1137Q3cawCEDLIRICPIvrHeFgw6O32a7Eklkv34sMcRTQyiYv4Wm/BHTz/9DH3wvZ/kOQXxit4ZDKKFjFE9TzPnsNgRcoIJMIko/DW0825b0nFvOyKAyZdd+lO64bpbaXrLbKmRXxWfN6uDRqIvKhEbhdcpiB7E+mBtPg6iorWFf7bor4vpC//zTWqdPpeBWQC87IBboFiBZcNS5DDrrFRFEzOSFdyMvH0dExa9fZ30+n0W0t57706z54CAqwkNzTHPIMiXv7ScFi1aTFdf9St64YUVXN4J4DzIH8gH97ZAlgITEXoeKVACoIX7HGqEq533coZHn83mDbYeZ1bYGNtW0dhxg3TAQa+nnXfenmbMbOVSdL7pOp4HzaAffeQxuummP9I1v7qBZRVjRBN1ZDwgAwhR5lKHvKTMUyHRLGfLlttsREcfd6CTrSvoml/9gaY1z6IanHX6/Mn6h8eLz4lMtQ0b2ujAgxeyfrHMgj/e/Be6+MJf0tQpzaFXhULwGZGqTFTEZobpz/JnjskD+iZ0CWHRsY5Ji+qJVbRw9x1pp522pU02nUf19fVcCs4ymXFlzHlHRyctW/YCgci/+upraNnSl7gZNMgWlFpDhs24CdV8LkgkOUgsa1otYJP1dYHstHesp9NPf18gKu66axF9+lNfpZbm2Xw9a1jtA4aywWZiS3TRRz92DG21dSSah7O/7ZnQi+nOO++mG264iZ9pYnUdTaqpo5pa6MA6bgqOYAWej6DS487jt8LGjHfmM72vhw4+aFc69FDpe/Ravn51zQ303e/+hOrrp9GEamnOzsRvsDOtlLGUSpLyLYUWimhXfMYgtxKPJsbQz5wBLnad+Z5sh3Hz4xiJbpH3EoilpaMtCj+U7jEibTAGyhoh4HQ/D0e1Riz7hDK7QuYyEZC1DflJAAzLc1hJHn6U7NoZdqF9Ogxot9JDRYApX0abUIsfqlkN2ucA74EcgK1kc81k3UA/2xYAuJngwd5Qp1LAdAG+sT98dgA/Tci6ML8yPYl5X7FPKXLIGR3a4w3l4mzdcE8D7mU6RCZg84O04M+V0GJgPfNvK1nMsqT3MBKaR6bkAIaBeWGCiPHt0ZwVg3NBmjcrvuT9Qv0tqkIYASLkAHpx+CBTFxzj+oaInxwrUti/PW4n+kfKQtmcBtKit5dLhPHahyoiIjCRsHLEu86fbP3YUNqA9zHaB43nWfu9yv6P3jlkmsk/jIeZBhA4Ik/9/WbxWNCw+vAqH2OrNPMnlGSLvUaLbZJYVDDBdIJtJc8pPqoSA7aerjxzXLosyjBIVtEje3+ZP/1+6NkJRFPW0uTTn1kmS2H+FSs1Eo5Jov9rRAWyFp677xbeFNJHId3IyJyYs93raeWzS6htxXM0Y4tdaeJkNO/KOw9w2l557mFa/cKTXNKptqE1FzW68rkltHrZ4zSxrpFmbgUAP71Of18Pl0zq7VxPMxbsTpOmotZn5Rfu+8Qd19LoKu1RoRF8GfODVjz9EK196UkaM6aK07DkFUHCiZPRD2MHHvOG1S9x4/C6ljnUstG2alSiLmAvl6TqXPsyNc7diqa0zKHlTyzm0lCjcSCzQhug/h6pp9c6f1eqRtmnzHMO9Ux/38+jMcgG8BBExREtq1XpSAMmaUSMQ9eAJMuk8KOOSn54RIXzIHIPX0RUOCRQa/6lMumP4VGZQiwuSjcxPkIOgahSeC6mIwwY47p2RSg1DjxtrGXAqH4v1O/173OwcAnoWwIeY1qKa4/LIQMgWowdpP4hZbSfxowtqyfrqZy4nZms0rAzOQuzz2oHfjz4EX+QviKIWAi6FZIOObdRZU7NglzpJ/f9ZI10V2civzywaWc8UhIxV1gGn0lSSK7wMNw9i0TAaRQ3+DA1UdTidUQEos71qcZJBlASge9/L3+XK6RR+fK+HtJ86MtQJLIp2HqFqiYcfLmGuGWgUUYCzJDNXj0hf2D8KB1mdTtzBGS8gEUjROfLUn6zrECxLA2pg73hYbfN7lEPzLv6s9n1FiLVv3SdPAhdQFTYdQyYz2nFMK+aPVOgi8xgEqdXjCeJripZuxIyJOzw5GcSCRReWaKCJMKrs6ODVq19hVatXkndvd2c0dDU0ExTpwAIcSB6bkx5okLOHCEzfb1PSA7X2wfg2rGOVq9ZSavXrmIAFlF8TY3NNHVyQyloX7zE+XICAhYDnGyjV1a9TGvbVrNuRd19ANHIiGAwV/tUqAZSslOixRCdu3rtK7Ry1XL+OxoTg+DAf2jyHYgbZ1f5qbElsohbAJkAVVetWckRteg1AwKoEVG7U6QmPiLJ8s6oNtjFeNpW0fIVL9Cata9w6Sdu3Iib5s7TrGGdVxnQKQDLeU7qm3lejICJtZOLY/7NUStURCVv+u0F2YbMAbxZtfplWrHyRV6j7p4ujRuIjb6LLleIP+hZC5AFGQX2TCjzJb0WIlGBElNr167itV2/YR03+JTo5Baqq5lCY8YrCJK9eTHykewtJgR6Jbob8r1y1QoGbeG412Oe61to0qQaqho7MqICN5GyZojIXk0rX1nOcgAHGfLY1DCNry+yKZGf2a1qJArARPx+1ZqX+Xog7RqmtjBJYf1oynqmVFpzu1/5NJWtXNlVi75vEYko0dHLpFBHRzvLEjKXOtrXc3YDAD0pnSGAE4gXyDv2PUgK7D30IcF8SWNdzSQqayjvzZfMA0oPEZT8gr5ZziWIAA4A1GxunM5grxGRDCD40g0FRIXNBgMtmknTtm4NrVq9gq+N50LPC2RqQB9Jhk5BDyEHMAx3r46YqDDDxN3AANW169bQK6teovXr17A8ApBFBgAyVyw62UrUVrqvt/L9c6QAtdhSAMoAmKJXDMrugdhDCa3Org1MJiEbJQA3DCqNZZmADIAAQAk8/DmhepISVy67xskGB0IoKCEyppiUs+FkaqLvZv8GeIfsJpTFkfG1cVm3rq521uvwWTlCO8juWG6QjXFWV9foOOv4zMS4x3EfgQoGbun2wnzFHh+rVi/nvYNsQfQoQOYA7mGZJMnzFKx7KLm0fi2tXrOC1q9fy+c99plkp8SzfeREhTVzz+uEPFGhI+UIaDQn7uPsJJaJzg1cPgk6GecNSKPe/h4uR+L9Pvhl0KPQGSiJOLG6lntRQHdANpBlMtpK9GjpFgta4rurXQxZA+iPe2IfrF69gtcb+wEEI0otgfQQnZ32XrBrRH0A20n6gWB+16x5mfVdX78vHezxILVs1EaATsd9kNUCuUGjbDwPShEyQTFuPJcNEn8j9kbwfnpwMXM+L4gKlKFqp3VtK2nVquVMDEEPS9CQ9orSfTJcfQS5hjxWV9fRlCnNNLkOZRlhj1aFfgoBNNYDyEryGMtZdi7hKUEAYHxWCij0DNABcvR9lUbnj9EeKgqmc417LXVjexVYC2QO/+Ymx1pGyHS+ySrf23pk6NmCamfIxuEsB/MRUQXNzosCogJrBeAdr2i3+VLf0XfEdzhLQWv9s02hfROsjF3O5GE/VHpuSD8I0XN2L5RJtbmz64G48Nc1f8b8QAQCsf0cmjvH/h6mm20PpXtAZFuICsFQJOtCAXRt5N3XKxkPlrWBsaDpuPWx4J4MGsjsM1vM95Jmy0KAKKYuQQaWMaXzwCWmUOoN+GVYB50n9X0Y2Nfo/4SUVyKBCU719TAuK5Psnbbg7plecfgJ2+Kuj4SpZbyHMwQ6Cs8BueYsmDHIBMH6ILjZsjxUT2hWDsbLZT85e1P6V5g8xh5DFiwtcu5tGtF5Rt4JeWOZFuwX6nNI5hnOIAnADJhP2BdKFI6NZcAd91Ehy7vAbvT+tP49YF0yiaEKiccr5FwfIVHB+KyWJNNn9UQF5jVLKpn+yNs3Etz5f46o6Ovporblz2rJELOeg1rjBnBTZ25M61a+SAO93VTXMptTE4tfg9TT2U7rVy7jptpMMmS8m56uDfw5SIHqOvRtyIIng7Tu5WXU39NFddPmaompyscQFmX10se4ZuvU1o1LGm8PUvualdS1fpUKir+vPO84RJY0zuAx93RsoPWvLKPxNVOoZmqLe45B6oFBuHIZExOTm6WEFDJOOtauoN7udgY0x1XXUt20OTS2JDJpuAfr3+d7IyMqjpy+hjeKNMeMdQhFUVoNnPw62maxQ2uoCMIi8ktVXgq4jB6kUZoSF0HlNGotA8Nr0qsY3yaSovQ9T2tgotxVmFrJszJyIuqn/PNmiQq5V9pDwxNzsgpZ0LpSSQiLJM5KRUpUJIq9nKfIlNOSa4ojJBkVPD7NlrBP7Tsyh7JvLKMiHZUZuNHhCQo7V7+/yCnyawHSCGPyD+M9fZWSBERWgypx3GN/Bxg3VVyvl9iRG11I6Ng9MmvNpEEhVxtXVMfiNWrZevNMZsYps6u1SYPAKiGYAZ09CWPSbHMtkRIaja4ZFQk5Uopdx8am+XXNa6Us4WzfSI74YOHHWUH5FvF70vUq0ntmiEpDd82YUKMnfJ/nUa8f7pdG/peERqn8m8bRK/rzK5Ev1RGZxpw+nTM7bywy4Rpp6acQM6lgghlzubF6oiIYY7o7vcHpCCCWJGvMXjCxCe/gPs+XzlChH4KogJ6HA9zR2UHtnRvYqAUpWDOxlqqrEVFqtYoz62K7x10/ODHOaQx6h31fBA/0cwmMjg4ASJ38rCACAB4KYF8CFBcscUpSRp0I5wT1lwFS4bngfOAeACYRMZ48kz6HrTccSDh/qHsOUABZXHCs8NtJ1TWS7RGigfPngeiHuDBijPdxFDiAElwX4AnADoDWAB25vIZGhmWXnNenv4cBWUQL40+sV0jVD2pP/5Ihssr2Jhy5agC3E2t57hGFLoCJ6XL3bF7Oii7odGLRx3E+sHMkPbynu4faO9czWYAa/wCe805BbjZK1QH0DOxfAEuQXfyHvwugpCUuuaQO1nYDywYILTiLAOQkqn48jRorkd6JLqxEHGaGCAcR5BueCeA55BAOotyjhsaNKyalSqY1KAuTIwCuItftGr04gccO0Il7r6gcZYkKIc36qRt7vWM9X8NKKUKu8XuAQmw3FgQ2lY0vvY/ZEflvFwOKlZ66mKiws1ZAfyn7g/2AuvRodgvyBf9mZ1z1M4AG7HlE8jMwPa6anxXvSdP1THCNH5YdTy6a0H9s6wLShNelCz7FIN8HIC0ir1nfcM8PAdPxsgjVrJPq5ynqji4GswG+47mYkJtUJ2vOJX/yJKfM08jIoZF+PzmEdVJszAC9AcSjZBl0CoBR7oXD5X8A4sU552cO2dVxdn2MTN70yTdQEdBSSv9AhwMohTxgz4AcwPsGRgJExNqPrxrPc4j1YpnQMk8YIwMuGh2NZ4g2sRIVDpSQqGdnMwS3LR2nBKhodkVPN5+FaJIM4BxyK3ow2pISpVtFE8ZN4PMCIO1YjFlLxxq4VckmKzIb2XPgUjQ9DNyD7MP9cQbgjAQpAhLEyknZqiQyEsRL7Ds553C2C/HSPwBZHS8g/4RJGq2PjPl8X67owzibMIhCOVFRKuJsRkvde3nOPu5PNNDXS929mOvuMN8Yt+07jA0gGuYcJDbOZiYzg74QIpixfAUipZyK7G2JwAYgKEAbR1z39ip5to5lEs8K8hIEiPSXkWyYrF3ugVp5DvQ6ATkL/b+eerq7A6nlLI5UqSqJhfHgeaA7sCa4LzeHHzOG94H0fcBPzW7MAnTqrQRfMtGCWpavi2WpqxPEYIeQbi7rVI5RRP8bYFncd8RAVcwv5FxI5hpuyC1nnGZjhRIxsS9EJCoMBopnUgggkSgajn6HPcpBguhL5MpvijwLqA4Shv07Zxv5/RaAWiUqbN0DUJ2N5g62rGTkWMQ/mimHgCVIFJcQUiC/gKjAcOTeEphg5ce8fepPANEr0R/jhtGVXvy8Ep1vxCy+jr0B+9MaO1v0twD8o9nW5RJMKIfE513s4QJfHnPNBAeuocSOzSeP3dXxj/1e1OdkFFjkCOvG91ZsSMgG0R9GesCX6RsQYB5ki/1ppZ5gG8Aet5JIVgLIdAdkldeISXCQCdLfyAgpy7rBTIZ5sn6b1mtTlVTISBgY4P1i9+QSVCgxBdB/EERX1LZeBYYMAE+aKxGCucQ1RfeIPjIZZvIB5JA28Ga9ws3PrSSqYGZMvql9wr8dGOD9Z31UWTsoSYRnwVkViQoZqZUBY/uDMye0d4XKHsu6ZTNpBgYvqe4tCUbVsXAvr1iencdtmQpK6GXF1591MVBAKjvImOxsNXxKzmfTtX8zUVGQUaEiG84Yy2DyGUTevrBnCj1G/q9lVFTWKv/59N9zBkZGVBw1o02UMSsUidhnhcGGSEpUhDRlTeE2UFE2NFONhVOaOp15M1gODH0fjYy58acC5ZxupmC9u7x3jsXkj6nhXnmECI2Am+G7oB2KiYoymRAw3eBo/wwefHL1+SPUH/m8AK6WOYRFLoKVqoqNm4LTeC1/9gAAIABJREFUWtjUN2N3BmDX6pfKjBj7nwcZ4vfkM1ubvCFahOjj4AwHVBhKUVaG2XFGVDijN/zOg1/x7z71NDruAYEL9+d6kUitDL05/Nyk34+fGNJQIKfyYLnRieQXg5Ah4l0P7YivqyzlgEMlkDLEjN9DWaKCzcMMkC00/Ug1XPEPYomAVG4ltkFeUY7SHhWeqIh6Ij8uMzalJIFldKVceGKPJYiXjFvmYWj4JDylJ4nsOdwUmGGQ7JFg3KayxDtlhERFsqbucsIfuvWTbnAFvIYZU9Gwys5s0a7l0jRp6kRYRf5L+FGBrJsjPyANaKU5nzT1w3++REc+y0P0jhFR4ohCb+v5YdE4HFAnPR04LbpfasbCacELxuy4KgENJR25XNDzwGhe9tipH5TGiAb8wHgHCMNOeQ4UUM1oDQ/VCeNarWz8i5MvfYXygEKWwPZEhe0RadQocwz9xXNcNVbAG444LNhDcMBQ4g9OCMC3nh52ljCHQdYy6m0YPEVwVjnSHIAMIsrVUS+bezakSy0CGXsZGO2JCnOgALoAAAB4xKAyR4ZVBlaz85rMmAKJSEVnAFqfyZotmtwYaGVri4AZrCvLBte9djtJb8hyXQCk2v390nHMYj8c8F4mLOCAQmbgMLPscQBJtG2GpdHNGdV68CZHrCPH4Hnj+vnG4TndAedzEAAD5BByJBG/KH0QwaqRHTJRRervShbptSQqjPy0rERuSgmQsA/zDlkCYOhBGLG1IOPYxyLr2pA1y+ikx0ByFvosSPuavQebG3NqoCfmk+Vw3DiOSjUg0uybqDPTuuQsfVmiM+gOIfPwW6y56GdEpxaXqh365EwlZKTfL5ZdI5BE92I+OPKUAR4QNtps1IIy7HwqISpKl4eNtCJ9IeeqNSplcqK/j0EtnG3B+efzHdl/AM1Gs1xYSRQ59wWgkqjdGMVrPpP/E+cDN4uNWGZuDcVKF9sfVxdAVYA6jI2j+hl4k4hsmxZrjs0ExVjZpwY2ZsGN7B4LslaiZAQ0Mn2As1/qpKPSgM1HFjyXcXkBNUtN9D8TtapfGLhDdgLvhdgEudizrFT6aeREBUfvGmikYGtfH3QCsixQNhnyIHqCycNgx8BXRukT0dOQV8k0SPWFZdizV2uArka/45pYKwGZBaRFKW0mULnxMoA4rKXoIlmnzPVz/rcBj7peKPfMvr3NjayLt+BtZYyAkDJVADJxb4n45++ovEcx8akP8TzgVed/5vedlPLpDySxzO+AZqpIoXmMlQlAbsAsjayLXtzwGL0PAOZqZoIAxMhEFPvSfsz+gYGPjkz2mIFaJ2qjqG5Ak2WU/lb7l/c+msBz8IKUvsJaMdCNPTooTYVjCbjgoPHZY59xA2Zt4mzlbqJ/J/see90ICQHZB7icDOZD7AMrDShTzfJRYCBy9D/3ART9L+PwmEXmTC6YcNNvhQshajA07BZSgdhWZ/JmcJDLCFl0fgiy0ouZ/sH4jNSw5syGeZhN6fWsrKmRwZG0FV5Y/sfVKNRmtCoRocywBjHgGpzhwVmPIBmklBaD72rb4z0O2NDeGNwrgjMCsGchf0pUKBHApa4UYB+DIOkeBE6CYJBxhv63ajOKbpEMeU9U2F7CR9bYnDNyWP9H6yLZk2b3W7CgQGrBv4aOkTNNdB/KleE9nLvoQYRn62jvUIJEekYYIWFbkf0TJfGsXKX1XzLdAvnkPYx5w9o6sokzvVmviK8XM3HkoSDn7FMZcaBBG1z6SgOrcX2sh2TFav+TTHZKma3iVUqWqBAcQvrJ+O/ZHpS5tk9cMELm/bLST3Zo+7Pe9m/oX0MkMol+J85GtbPcznDbD0ww/YeoKLFg/vP2v9AMjIyoOHrGemEs9TAXY82Ye9mI2UMvmsUuZYnJBdOxlgWgdR35mtntnskgMKKCByLUg49I4AiaoJENmJQ/A0gcmGNnLIVGWPEw5+gVFx0gdmM0fNng1FQzMZZGU/8gGmVlYdkY6cOz5Aw4OyDj+2r+mL3CETQyck4Ddvactw8sqsRWgiMicuV95NmErbe6hcmRpfrUSA8zxWweo2lmDdlsrvOOhx6gvBbeoNSalDA2OeIEhkFsFheMAlXiQd4SEiGdw3RTOdB0jIyBnVru/WC1FeX38h9qAosBK9/Lvnzj6vxnlUB+cSDj3AWIQ1M04bTx/Kk8Wpq4Ze5Ido4tuO4uK8kScIcI9Kl4+pnT3+sYeN9lrPih+pcUPKAYuHZpN9/eMXGCir9K2SGJsEgIR92Xfh/zE+seztvAMYvCHDkNdinRrWKyqraS5eA9nI+czC99Xu5F3Xi9URkE9ddMiYwwgWHPGS0QtJZVQMrdQu/vSQp/I6vxLd5uHG9QrdFo8gaUXCIrH0XuY4bAzJBy3pATwM3pmLDvUpOuaN9F2U/HhZR/S/KK5LQ4liH1XX8ijRBjFJw5117G5Bxz6xH2XH5U4r9rY0UFiaIuycydkY5uF9tvRZHj+1EXFQlwEaCTLrU1eZSzU84RJT1MTAr2MKep69nGKd1I2fYgjP1WJ6Zcz6ejtn0cSBttRlmyOQv3UiGIVQAepo6XnvEMYmCNBJjzxHDc87beqhsCC+PkFHOWlK2Ves08tpD9ZY6i2DMGEto2E5AoAk5mD3kd7OWxbI7sfS55ZrqRo8JEdljGObkjLPhQlxIJT+rzmt0j0XNSZVBlU8J8Ncuy+NJhT5i95PZ5ERhSkRxyt6iE98se5v8f1vOO5EsM6rBTLNeP+9bOEm93OrmwvVY0JDWrisYRLcb4qezPuC78ia05R9kaiGF6J7Vn9euy1gXjiYRMBCVNd6R7MK/XsuC13CtLbPunyv49+12vf8t+p064EgbmfxiGxvsK+sb1c5AxyStXObREdFJSNp6VXt+Ec0AzuXAPgE/x/HQ2aqb0F2SazylHVGTXSEwpRvPUFvKEblxMxarsCaP/pHXgDeC0X9i6heaeCmgC1JLApEx5yJKAjrxERLm1PRl1QgSiWV8ZAAr5zvX7M50s1/PjluuZHornnD2L6PtiXVCmb1Jb1u1MMw8zP7QyPAIQKoniynSFfYFzyC9q8ANMp9qc+K6uLKW87hw0IFMhZwh8S0SNazaO+NAiGwI+6ffUpzEfWyU/UTmwk6z0q0XtM7Co+kSG7WSM3/BllmWciR+vfePMt83rh0oSY+tctnaaDayryzKtssHD1Chu/MmgKpNuJj3O1tWDGVHsCLaUMp1Sxtoi9KOPKL/nkkA5+8nbtHqq22IpEuKJw3jteKbg3pKpgIh8IQTCeaw9LSxLznodBNBdxyNHX5yzSERIVLtlFmChOBBG7TspDy0kqOhKLfVjMspqR2fYbCAoWbU/okGt8+BsRDs3bKxGHMQob1y7X/omKOAs5IGcoZLRKzqC7XkNQhKCSchKfA6iSUgp+TvfL+ObyXzEaHfTDwIg67zpHgtERShJFOUGvA3uHXSX9orBfMqekXmIzbytb0UfjRsHH1/JHsVjrOE09BZnSrn5w/OO1SbbsMclAMn5nCrDMr8SECJAuY4jHBtWPknGDRmwkmR4dimRZPscn2FNxvD7ElgmeBa+pLcMJcm4jy83sBbyBTPV1d0dsidMnqxfCDKKrYE85grkILIpfPYnlwJTjIaxNJf9IiSZrFcICnR9G1gzsXg6Rl8ba0NnGslmtvuABrIZ7mJ61HyXnCUSMBpvaYaNIXu3IIuIS9PpuL0+FIJNnt/rG9UkKQSqtwn+l9NF/prmZ4RnUdk32RRbPva24X//h6hIzsX//ONfcgZUUQdQSwznsmbab52+IRgn4Xy0aBFnExi76yMT2KxxythHuuN9jkbSiKiiqYqGQtbYcYZNOFeyAFj6G8/e+oMd94WSFvZZHKJikEiuJ88pwCsOG/yvqgrRLlKLML4MQDEHQFjjYEBypKV8P9wPQGowPIXhxy9CQy7fcNfKSqXelY5RRsLj01qVbATrQcWRA84xiTNVVisqAjupQWp1zcNTBYdNLm8EgUS+SCMNRL/0MeuPA48dJZ6G1FHJptaFyGh2/sprWrHPqh+LfEm0I6JOpL+KGIaYUyaYYPRk7GRbjzKw0OQnlVlzjKWGau63bkxigMY5EwDLlQLgyfPf0O9WsPnLep5k5TH+Wx0iN47gbPNSFNzMgVG2F1SA5SpZf8PVZJQDUzKw5KDlXRSGw85PMqG633QYZlxFAFC/jz0hlkZyLXP67PQPEcxs3VR2nmynJ3Olez44k5y+XCyHSTsTdyvv+6YAuZmEfp1Nf8TxhktVkgM1rsL6hPlzTdPMVs/0cnEsFE9RdjnD+LlklxjBfiiiz5xOC/vaq8XKc5/uqcxKhXRbccgsqiQhnxyQwHKmSxTlzzvjsu/sZSBAdgxeuxV/Vrw/i4Bakf8KNfkKbmDZg36clcaRzJo+njiDQhoKSCMN7ix1vYyQGC5RUTSeMv3JsllChMgp4HaeCl3ijJeg2Eb4ZsfC1+PriF4OYI+7k5MCUWVFsuu/n4ixD5LI3L2QEM7aKl7TvAr4PWMD2NWz+zfcJQHhvPwLuSe2gc9kKtaYsu9K7lLGNJR8/zW6zBDkRSXdkz1vU51ceb+9+k9NrkUuU4Cl+KpF850P0nn1Iyo0Y/ly0BlMoujUmM0ve9lBxQU2aX5Plkpnfuh8rIRDK+prD6w6eSszX2Rjl8+q3AJgSbTfKoLghYomze7mubEMcxuviZYSEmVrVWSCOeUUfzYUqxcV2rDFooiQivpj2JcxuEbkR8fJkfHaVNb7Oww4G0mX26rekPIBBnaey8IOS6qsObUMSmVbnin8XuXNix2XEeGSgEoWDkedFExVMakie7/Q7i55Kl8GyW4TwcuCbaQNcfGJZHZadrKPuo6/G8GMRtFAc4QRvKLFWL56bPsnZ2/+vBXQu/jeVnbHFjr6j6PEL9Tem0ws6CUsWEwCQGIPiGAuqqCUEWQmTOXlkKTnp+wFAem5WbQ1JuZI6bSJsw+OtP1kz83ElWaO4O/o98D+ifr//Lnz/833FcLQjOQYAGC2q81dOB2d3WbBIBwWonouBN1pY3EGjFXO5Hsot9zHZZysXBIHZAYHMDZe5ow1ZCSEoA/r0SBnkbzSNUemCoP43Icr9g3N6rMYVCW0lM1n0NecAaNnnfp+cgyJ8mb8R8lCtqm5/4iUk0YJUJ9dg/dsXQ2kt4wQy8gzckqyb2St7JUC0xKAKZlwKM+FdRa1IcGesq/tekZmIupenlFKU/G8DVAoU8UllpBZyRk/fUqUylqEjGvNIMR7nC2svc4s2Lanp5uvj3kQAF/kG+PBZ/y+EvDhLNCMISFHUgLOP78E2Wqmj+ouZLZgHX3pJ35G7Qfi96r4PFHB+/VnL9B0RzLv+KD4RKl4PmbkMuIdsWSZPYtl3/jv8DDLDGL9rOhztiFlkQPRZMS0VRvgj/9DVIzghPrPV/9JMxBOWI0u/tuJigA6QNNkWXbnNUsUPdJkJZPCQJKyiRg+UeGj+HG1PABqB7ptZouCZJYetfRc2hSnh+VASHkQblCFhj3BgpX3PEjnD1A72AzUS+dKvxmUpBrN/G9fh1+UMUduhWgs+W5WYXmQAiA9Rx9oORQzVvx8p8d8JaJCAS49EOXeVl7DRWO50i2ILPV1LDmTQjMYjFEW40uj8oyI0eeXc8VFtviMmCyipQ+FA9vWwsBMNgKZrZfUxND4SUE7Tf7Vg9wDNyMxuouyZ3RQehkjnMRJkCZhBk5YRLSGa6n95cdSWV28KqKCTy0vre4fhV6y6I4wKrdOIowZadJU0DTqwKINRMbtXLWni2ZB+tlwiYrIBVqqvpVZCB7IiIkKPfdDlDTGKOmmxfJhMWgpGeGspMxzlxEYBpyYPkvuViKarA8yn1kkUaJ7zDjL4HPBQQn7SFYmC9wWkXFh38VF0B/bPtA1HeLk86Zh8ihGNGokXSQqZICs4zXSJwBMJtIBCPSKI8qgyWEF+3CIUYejb4ia/P9gosJtWO/U4m1zaHwDw6yz/48kKrIiHR3DeD5UWoSKRIXqJzPcswCk07SF8h7vqzowsxlLHYt/FFGRAWq9tsnNWU7ITdeqHeNq/KpfXkjt/msSFZUkpAzGjMBXAN3dHAy58V+DLxjxa3qs/JL/PKJCzgEJ9ZPxiuOPcnLhVXyYZR6nIryXf3QDMIpk3JBuO2L0z1KQv2xipaIsv0L2pz5vmV7JbQqX2STHcEylYd2rc8c3Uf0hAErxYV7+DJms0H9hokL0UCSZhDBHxLSU6wj2vRpZloGbLpOc0xFcSomKcA8jF4baj/ABMt+xFUh2l5NlCRqLTYAN6Ge/cVjsiN2wRPY1SK2MEi56JJPLsjO78DdaCsxAbynPLABn9uXP36GmNDxdCVFRaYocJJvcxquSv4Wo4HLDVvLISsKFZVPsIPiztjclWt7OA55rwaidrvNqTwMP9TtGdgoonH8NDEiJpkgWRbvCgiWNdDK7zXxlWyv2ZRW0xR0MzMX7UhJJ9leM3NeMCs2gsWwBwT+UlsoEo7GdZAthGSzaP0EmQ/alDzyRcWlpLiMCjeDjUpF9NH78eC6fZL0UGOxXETQwHxOOckNSXkzwIvjMGE7sfZXqTsmvkCh7fnYlLQLBbueD37TWoNqViTVyLFQQUZ2N960vBp8Tmk0nOk3ubWvC5fcUrzGMyfadEBVofi3ZANZomss2FTghtgbWIN1sd8uIkKWIfVAwBiFqxDcKQZmaLYFnsHKxCJzs6u4iNPQeh9KS6kPauSRzhyxT+VNIJmmoje+jJKk1epc5GU29/VJ6CePCvS2TwsuTBWdgiIyFlJyE+I31d/HzC9mQx0O2RswU4Qokfu+qbHM2EZfr02mxvGtv670GREW8d6ofOAgi4D5S1suTWl7BVCRCSrIdfbkzy3gxMs2fEf8hKoZ7mv3ne//EGRgZUXHUtPV6CKlxyOe1RX8ZcOlKBknWWKgJyIapi7K1OpgGVDNIUmLpiaIsMuJTMM6+Z6RAsiktxVHvkaQLuzQ3VqSc2lZ8UMjPHZxh5YM0G0UOrKw5JgC5vBztYnPiQDTRuPKGGUU+bROHBQ4pG4XMa0pUhNHpZzCWwDrjFdLtXNOgFGtxfUAy0pktdcVj4Og/SUMMz23UvjxMqHVs64Fa8mNQg1IPGJuXeD2zBGN6cXhgP4Mh+iK/jZio0MPfml0lz68ZFXZP9iWDHxUWxN82d5NiINXLRp7wwaGKqAY+tHukoa6lsIpsSKSWvZJ72KUNMS/QHv8IokLKfnlIT/4eyLjM/mDj08rM6D6wrIqwJ6LQqtSkyLkPdBCD3UVj6zyEX3iBtqgCre0ZdifswgKdkl9TA+8cSOoyCHKGhJuXqM/iNWSe9Kkzz8yufKbygi+bpuEyqUwWYxsVSiAIUWfgUpGAh3lRksLPiScq5FGzdfHzBElEY0x16nwUyK9/K5WAGPUokSJ6tiQZFXmiQjSQOo+qr4wUjHOdni+V8J5KBIb/XRnoFJ/v709U5E8cnX/dCya7nqjwqdXJWoR9WyJwFdayLMIx6F7VHUkkkN8oerJgvLFhZjnkUQooOmFPHOoKGRX+bCqeD//uSDIqsvOY/pvP9JI5LVuB4vOofGGy+sme1aIETUPKfqmMwo0Qcq4wqBGhfZUergJuWD6zWULOwKEhVNVr+rGV7ah876Jn+MdkVFhmAGv/UBPadGxBScVShfoqpMY9dglWmGKIJZullBQIkYpCVHgioXQL5O5h55tGx7Oic0aKZqN4YK8iyF2Q1RgEbliEkBPPIfZxVpBLd6MnW4Yp/VIdx8rlaRkcBIMZyMlGuPo+XMYje2E5p0Vq/ArGyY0kRhx5JY0SQP6SZwi/DeCjZGGbTrRAlQBgD3Mu0twAvz4mM8M/Z8t2UZnOBlBnzd+tlj5GYJH7RY9gwO9wH2+wjKioIH9FKxaw8WGyQJV0phEVwQxwiYCCQ7gSP1pOEeHmCVFiYLYnzMTI1KhuF5Vv2fEIWndltRKLgcvAIPpfsBQpCySEEds77AtKloXZLP48tu96cJL1spakZnuOyxuLfo4l3wQU5pcL+AGhAmCZ7+/VloGitn9DIKoUx/KRbhYQJUGgQl5Yo2h+PjyTlqYznCVkUzC5oJZI0L9CxMhRI3OBPy3g0PskNrdcJtPIFWSTjBG8wYJj5bn18V2B0BSc1/OUyZO01A/mDD1peERhLuSCRjBJryeQD9J3I2TCWJkq/NY1+cbn0lMBRKj0uCh6+X0d8Bfs3zFjqKevV7JV+tEHZRw/ZAyElLXAeGLfWOlL1d3dzeNGVRBuvp4EjTr/idAXSvSf9KmNgL/Jpd0PUgGiAr0sYoaNBChK4GxsTs69bbS6Ct+74MGNkPMZFUbiccaHl3vNeuO+GFqtJWTGuAoPUa24wAvdEzYElq9XlVGRVsfwtqVBOKHJuAsi/luJCpN723uB6ASZqdkoLLf/yagY7nH2n+/982YgaOlhZVTkiApGHxU8sjp2Fq1qpSU8AKGHTig7oeympZRx6aecEaPqig3cAtXllIeZrVy/PETfu9/rREcwU37Byk8BECv7xL/SGnn5aGk1pEV7BYUuBoUaNTmlZg5kUb+DWHonADqeqOBMDwED4wEV69t6oiLinulcsRGg88vKXFBerQfpJDCgwSlwZ9/wzLcoQ0lVRUmSeMCHb4tTEVJx47ODqIDCxDoxQ66N3+Ra2bnK1JNMNoxy77Jgma2khpkdUhqBwQRJxsCAHLP8hSZ5DhQtocicnRPuLOvnx5ESeRgRNwJEWuRYGCWSxshzp/XU0wj1zIntHf4Sg/8fQlS4RzSXXM52M21TOfcptXGRjIzx5nC8cCWQP0dUxNuahZvKggdZVb5GsSNV7AwGQlXMUDVG02juYJxq1I7Irt7Wyg4ll3fPpkRLHGR0tPPvsZYS/96Pl29WwQXPfBwdeHmOOP54jfT6MpII8vv5is+SZJyps5bFpQKBnAMY0n2WOwsLQBjhKIZHVIQIMt13otbjc3jdlJLPxSSWzUelM9uTPOF7hcv0jyMqRIrTvcXzoOP6Vyv9FM9BG6CLdHekRdk6FIMqet7zIsa9yufYa0hUlO3JPJiU1T3pv18NXJ9oUk+Ylp0V4bnTM0sylORJfP3kSnL/KiDnkZm+w2UI7aplzzzkxCoIqlMiOqKktF+FMRWRc0ORPd7OMmeznOT75xIVdjTy3FjPnsQej8tbPuWvQmq8SZSR8SL7d+R3iCWaQiZEpuRMXnAzzUf4gWU0ZhKFDEXOnJCGoPwt6yOnPlPhpig2U7REkJvdSgz7EPuibDOWrl2Z7FfYXylRIXOUEAtmN/G8aX+W3LNnWZton9n+StZ8CGA8GW6pnnSz4/sheH+hZAJ5LIVzUh6W9/+x96ZrkiU5dphnRkRmFucBpCE1pCi9kkRpuIjS+//jcLoyMjZ9wMEBDmy5fj0quytHiuivOiPc72IGg8GAg21d9mkvLvn4Ub7s5I2xCSK5rQk2m8saoIeSKuOP28gnHQV5LwvHDw9bZWz4PmnabBHsyA+nQPgIFq/noX02IsDO+zUww55gfpR8c9EWjcUp8IYo5s5reKuOhYD5zjGKEjysz48y0pAbdFSgz5Vm7ujZwDVDhoHo8k02Yq7sO2A7hqAt8IMIALEsASsnFP0hYjIxHuJFpZNhnIO1RGwhnLHsdYHyVrHK0XzYezp4Sagqdwj7H46BslFQFuuz9ZxMR+a4r7qgcN4IAWz3mH2Phs6oYqD2EJcWdlbIZc0ScUA9nC7CWJ+tdHMG4FVQrl3iDofgK/vbM0GsWbZkvtD+MLDa3soeFwTtLco+A0uP5Fh8504RLwf12XtCWIaEj4XZPIZz+Dgqg8ecFn5d2ITGR1wTLHzY9ZER4ZkcliHyYlUx8Hxm8DDIKR0VyQtoIG/ff/n69WI9YjyDxvu0oFepBsGm8rmQHXY96cMeHcDwzMsYFVqCzuQVD6YAPOfXyfGMN5Cl9X1C7z/iqOAjwVc499nbBHsXWUdWaovOxlscFSs5xylpRlbuVZURH46KHfk+Pv91KMCDJ2I7CJbaRn59vry9mDB6urw+P15enr5f/rf/wTIqUNsujmP/hwKYHlj33gFVC/AVB3c174pGORIVbcLHhfqkDMXh489aaOthGKWTwsGXbnQTn2HUDsMEHKwLIJ3Cy4SwHWImOH1MElFV60YDxEowoSeFHzJWq8/H01WuGQztRi/mHIdjIZ1ZX84jB6JvBgFGjwxghHi4ZhN0G4wVG63pPmxe5YdI1O7Lev0KZPn0NgBuAr7VHNsPAx+DNDLK50FBslOCEQV2vTcSusM77ED98vCl9QSBUNf6wHSIjL4sGikKopI9cSD4Qepz/pwNuFg2y6MsIpVRlYqeLXB9x/JAnEFQyYwg7dwfgj1Ax5iPIxwpmHecnygRHttNwOF0Csxje4+joj1F1j+ouyBAV1bBMeVgosPJPw+lFKmfOJhBiqoRD35Tg1PjzepzHLZUCNUgaAkewx9xU9Db90PUgl1mVAgoofMHm5ch4cp17FzUtIU8KRxcwQtZO61zu8Xp9XqJyiSNZEW25m6TA9X8j/swo3tWCnDb/uIySt4gWDACNAE8yP0FiEdq+ORsOdhfHFvMJffFjY4KlwHuRKbxUzK89mxfo92ormdKLH2mi8ctZNZ1UdMefg2XyqXNYzTmHSn6NMp+tdJPPIFMTIDlhpI8Q+3ekWxbrCzPShq8MBIQbaBaDUdAnhjPQzFo21frc9OfvCn9VOBCv3cPUK+ZxGexASp2bLUsfOKRdHCeZwRmgq4HKOTmJXs4bqNj7ACxnaG+2wRAKU7tqLwo+rdAhsdeccDktsdsr95hln5DZdMlWHPQ/2g9t2sZFTfSYzMRBpMoj9Io5pmvt+4A07OOmy09dWF2iOYZ8FleADtBdAZykSvctzCC9KjwW1Vnrr2q8m1Lj81rgX3Imp6Xk4e+AAAgAElEQVQZ3wHgdTOXL9hpD8yHaRZ0VGd0o3fIaPao6GPi+UVZPeqGIm1OzJOOkzYN1TkUrIqB8FoGO6HUyH5f7TMtDhwVG/trDuSLQS0y3ghm704L77NhjYg9UIqR4fu53Orw25FkSyqVjVdkvevwocfbuKB3l26zFfveDzKsjdDlTW5Z5Ltlt9t3HvlvoLSDucz66fb5tN6rPRg6ypHD2fjv6Uf1tDT7iFktDr5GWVkPJBGnGL5DNgRBZvbG7EOhDIK+wp6Mdh9LDGm5a+rqDuVKE2WIQ9CAnN6dMd1eYW38zGogcGw2eAQOomcBSvAgWPVyuWePT1+kwGcc3DUnRS9LZvvPsIOH+4fAmrqQHB1rXlXBx4FI/jhxsT2CKegQ8jMsr8HvthbM+qDdZzQ0uqAkFXQmo4ut4eP37wjGzGBOPAOZDta7AfMiaG06OEsj2f32nB8/Hi93d+h3oWswnq08j9/e4KxiHwxgM8jm8ebtz9a8He99+PKAoNBwCJnDgu8wnrA5/fiBzIuRh23ehpV9+WoZG8ZLdq/1Q3m6fPny1StG2HPNQeL2uhMUfRlQIsqyarBnvaF8yCLlqZWss3HY9VreCfvVMkDKCeC8yvK/8Q7avTYUlOFCH7YWwNcJK3Tf6e9d5x5lLY46nlGlm9FpwQbyjo8aLpbOxrR8jjOZN3KSDlwdD7HDZiN8OCrWx+PHp78SBeLIITAXm3vbTPt//KcYPAQMAZ7QKyPit6KO27EWG5GzdwFJcP4SjWXMUXFkBwxfOmj4hnTIzHqQclQ4bOZIuHxvoV7tEMimQRdzRJTBXiuHA9QO2vv7L36c0dtuB4V1fAJN2GLK7tRx9Em6okXDOFMlI7WYh6gJ1Ii4AsCIzA2CpzxgGrgh5WksRTGB+PCMI9AnFLBJMR4AyDi2oXggAqW/q0r7VGo35pwKTtznB4UpC57RiiZmaK6ETINSsKvhqSppfQdp5L40RxWA32hl0SOW0vj58z1qJIZzheur5U6gbJSzQJZgaT50JwW4ruZdjYadDkZ7iyKJCAePZvKG4veopenLsXFU1ObBbzsDHJbvgaCZQbd2cX7dQbqRa/Meda6lhIjSZPGdRVOA5OQJOK/Krt7v0zHSHdPGQY77qTbKLFYAhmYR+EMiG2egVAN30/7E9emUlUhIWwekV1dOV+7nzVpQeR2XdORtn11EGGGmsgr+EqkbO8xjBjpDIoeDM9OmaXqkBdIlncbSFb01qlFqlOeERvYTQ4bOlqgfuqh1VTcraEDectlae4y9KHSf8pmaDQfDpRRA7tE/z1GBvb7/0R3XF6fYm9esgRLZKrVdG/3LAGeUFeX1yD+7zw8mICKi5kJjrnhf5SU+Hd8NA1qAwjCitwDoalB0Ugz7yM+WZSS4H8op0fojyUszn++wQjbT7HNT5+6w+8+AjoNzYgQRgppbwH52VCAgpOR0YbOr42aHE+tM/jRHBTb4MXuuaDzKnOiXBb48w+37a/Tsmq9aOSr2jWFx/zi/844KghvvmZHeWyBJjXUnO8Z3QT4dyK7N7gshMWzJeM6wSKOMOJaYEXAhT1btYrX8ew4jGBZ+UHVUxLoBjwvZxlKvS9nVxR91Hied8Ks86hoTXt8X1/bOiv0I/GyI0jIqWvZE1OCRzwiU4jXs31E0DfinzWOXSaF2DvVwBq6VihfnywjQDpRiw9Z0VFhzWq3fP14/0jHN7h3nrPVSe+y2TJXwvPL7yPv8u5WWlbFjLyMorByn8fsBxyxUx6uid3qc9+YYTouF/udyOHjiJcoZTY4KPlxInHY2ZUo4d9DMHbXz7dwzENmcOGhO3G0LlWuqDyWdxTnBIShAOMkiN4oQvGUgsh0wHpTIYEJZB0Zbc+0QtY6SRm6DhG1egWBxXkVlCN9HNlcH7CtLhFiGfc9IdZT+KacOxHRDdFJuUQQxQI5r4Z+7TQ8b2Gx+lgm0MtT+d+AIAKxfvV+FlSBiyDuCwYDz2A9KIQGXgeMicJEQg7ombLDMfW7v9oAcn3s55jA3NCqxoRIL8HVgYFMEx404RGqHERCJUkg2PmQ0fPliUfKgG5/LpslwfBguYdcgo8DoYFkUBvTb3z+sNHT0F3VHRtrToOuok9tz4HgjxlANySlHHfOIPWTYw+uLOTbu3Flgn9t4bC9YvwnLmOAauUMhAmTJJ7ZW9rvN08qXsSF42sRm4UQJdfauYKm5dMiZ8yjpH7hgeje6lOD+MzrYOuJ9dRJkWa/gVZbQdAeRNeFO3ArBCChWjrPF/2X2iJxtKQMC01P7hQ6HMk1Gm61wkMJMjY+fMiCa6244mJdEy6Bl3EtZoGe9WrGrU4QYGqt1kPdcdspZ8VH66VgN+vj2l6BAakynSj/9h7//5xCMAHIhIAgsi0kfGwHxePgZDbwOuBUx5k1HxRRbU6DAeHC2q41oZxNeiJDAtWvL8ig6ZBwbI8VVwWXEOOShlJEI7//dg6U0UtGxa44cFXFoRnMj0MtqOMZBNNuiUF8ojEMRoGaoYAVnv81Q3hjeELwAkksw68GYalj8EsBNKEXOGRlh0DNwcIOtwKqNnYJWdIjRFlNCFIBUhrJFw6Depyke1fNEDdhwZjhBMB8exKZAQEkN51dksTA6pIBozqAic3Q709kSDDqctCuwo885GybHFLfmjK6dGiq161pmRg1kXPRNQUiPWpcjUQ84anXc3xmOzEH3d4xrXeDwyEdF29lGCYVkgxbpnm5v13HLFwZ2617n+2DQwPlJZTulj0f+jI7FAwCLDfsGea+2awP7QkHqU+yyI6dwxVFxeMQIHZIGO1mQAD9k3cTQCxmrMqjtg2AnPz8i8y6NmWtn4rTuOol58Ckh4r65dAGvII/XM0bAR1/9hzMqagEvlzc4nWs/sKZvOWkJbipOP8qWOgtmuUzeTfL64XGN2LXUs8PrxL0nL1Hl3Vk/M14GTosFyCi3MDR3vSi41p23eZ4GRainpKAZNynlzXh+x/l1BsiTR5aztjvXd3J554TxXbjrGbGTjbuxburuVsTIKvszNDEnT+2h1SsQXa3n7+BsXfDJrZG7q4jyOWKyMsokJjQzLn0YB+tZa6E8cd0PMk9v7EFUModGL3VL6l67rVR9LHbOpJVAx1pwT19zPh7x4OhwHP8+KQLWokgypsBm1CuuOW7mtzZwt+kwW8qeHXpetxanTUFrzyRIZ+CQRYce99SBtlzbCLoJy6gQwMhmrg7yDD3Emt5zML0EeKL8Cv9e7VOf9OYgYQlIkw+5dKMciIeuStDmMYaAsIx49rK++Imd2EZWe0gzcutcYWQ0wNMOviqfHfG925cPAIcN0HX7IYLVzjAOM07K+dLvKorO+9eb2MZ+0D18zTE4OywQFKZORjwYfEaAC9HL1a9gNT+wAUatZWp24nT3OaoGMMocpY7ZvDfnGu9KhwbPQV9O0EvpqrQGDy2MaQGRveyulGIjQA6Si34Y5W/sE+8lYHwgpXNICwKGvFezzspZgEbD44/JCKvtbzOqXgVV09+Gow2iEe2Pp3iEuoOy5dzyz8NxwCwSOtt45iafNKMksjFmBTSdGR51uCqPODrwRBY8PaM/Ix9rgHnRHqWpvMKFlwdir4Y4v1KuhD3GRvAszxTy0fRAgvAmL+134wOjJ3nbqxpEJLtNwZuPG2AfzaFtDarHA2SG/qf7kNkpPAsRJQ9cwRbZ6K5Nk1l+jRVFqnIGHDAWYGqOCqMFsyQcbDf+Y3+RLgGxB7zMV2SQSzltB/Yjs8TwO+9d6g4IZGHgXvARy1TZZyUPbB2GvrRDAKCD4rLJfduZsyKcOLqXTCeG46T6aLgMiXUc9wQdTKzMAH4OHVX6naqMoePG1jVE5+WzOWa8DBRQSsiOyDiK/qDmOCSOxBuND00G04FjtIJzKDCDcISAPxCMuZSZGyHIDBv7WnEpZrwTrzo6n/g+uwZrarSFjakOC6fFR0bFcn0+PvylKBCH9smMiv/z7/8iigO80xRs+KVH4SPolYYRJ74AlHh4MeW60Wi8voOLn+/RfMojBVxIIFoAyqPdO95/mHs/RXJCQGEak7HqjgVckHZU1EK3skavz68uECF0VdHpY3LI3rzr0STbhGDPLFgorFLjlh5lFVAOqjM6ScHmk/z3oumMSL2og29h7CkwyUOaDp6xVBiGQDdWdz5AcY7vPbKTWRK4q1EiUkOTB03Bvo9SXHaAMVVUbiJPwOkUjoqIYvEDNQ1AKN/tYBhBoHiGc1n7bm2g+twa6LvaE6765oFaO2heuP7KemethVCs6eeLPTEq8IxYZ+ZCOiKSyxo6X0ZCfD+mRg3PP+uo6CQP0/QKGFdf72UNRglnYAgxROcIsFaOuopMgjKjf0ct1Y1D4jCxJZeU81IZo7zR+Sn/SjT9DOrMXSd8NO6LhbGUe7X11Jhlcj01gIThktx35Kd0BL15RM9mSTuPxTMR/WIrUS/hb12ahMyIfTcDoOM+ledVkGvbiyHtl1J0yk7Tx68G5pu79/ABUEAgPd5WLFrwTBeE4rQeZQqj4tpi/1KOCp/lALxTno7yPgkfiv6O8y2arigxyMakLz4v43xY1pBh4M3R4NhnMi2Zw6NhaSidc1Qch6TaoGr2ecTf4qhImbxjzrEWfJTmHBwPV/fECJpeEYrvdlQMzixfW9JIDWfFSwdAZieIEiBcBN2s1vvA5yHrttDrUs6qRFsL5tlRobIk9HEdHPuIhSOegRrYf2uu3c2jO1FqrFsn7obFdvuXezKdHwFEnjHQd/vv/Ofbg3D7iENHRdgIerPJAkROn3VUgJspKxVgvs1RoRk3i+lQp+WZc60Hw2YBCRADTww5q9mfuVdDwzhgtJY97oFxc8YdZ9KAaQj3Oge81Ad7+yFAwABAlhz2ceZZe6BTxdhZCsbtryihcpbHlD7TPQcmqjoWc9cxC2HQN0ZHiMrV7I8i4HKB6cabaGxLW5r26VLWkc5S2YBA7l42LhwGkclHMFKdJWpfqWzIIDLqEMOau56ousLGUVHjhfMmy1Q7gF3BkCUrAUAze4BR8l7Gx8rrRKmicraAEllmKaoaWLkpK7O4pmt3arsspPMmbnAbxXWLKmvqcw6HBEsLU3Yw4tzm+P37dy+5PJ6TpvbQFgY5wZCrc7loa6PYZMUfqBcE5u09BOsBpmIQrAJhTg0D6FMGQhL6vvvx49H51TJLQAvoZvbvy1sA4eJIIy/ZM7nnsY50CAPYZZNvgvkaVGN0tOff3SNQl30WHu4enE7IijAnDCbvJaBiTQycp4PJnAb2bjodLAuDNPeG2l6GvIIp7bk2DnN8rBtts2RXlUMjvgQa0/GIcdmYrGzTt9++eemzu/s7lCB6Rnkqx9YG/Ae435zNofuSzg68wxxQNg9kkBDTse9sbrauvlaRcUOeODrrtZwW6PV6+dR0PJH7YZvbnMBDaGBu7/ai7TC38O9b9YqwjBJkIEEWWrAlgX7t5UPZ0fgjHXS36RJj9gRKh2EuluViPywL5hU4lpID02F5ce4HLfFGHvtwVGwI+PHxr0SBYPMbHBW+KaPxEgHo9OQTnOTeDMF/BBy60KByGIdP33x9o2cpp/y4p411IToLiV0A4RiRoquUxlIqB/Zcghw4MAvvtMbYdrB8ciPEDys7IMxL7xctBFec7zSG0ehJAdCFQSuOCtbK55gpdzkoKjgrzlvN28cbnncTlH7QxgTZj4PPmkYmBojrN56xQEWsa9IjaK/lJnh6FM1Ke+8gVqTw2QHoTcch2P1A8dIyjEDCiJvzKoFeHFw2R1MUbM4VsYa5TxFvAtYkuyej6zzxe0UE0UEzrgbNuVL4+r6YV2/nqIiJ5ntnG3BcNe442XniqOg0Ey5rDivuBz5jwefyUd8L633RFWPSEau4/tlpxHV1pxkUrvxpUZxImaX+kusX5bmwlSm4DmpXb/UUnU/tJiglnYb+7mR/gYL+qKNiIOVeBs5jUp4eewKlj4r0cSIqfwRHReknyKf1DyOsGgAmjX51CgneUE6LvMauWxjH+drOgyIaYh8JD21Gq88/zLpoYnAAF+M1vZTYysnd+WfGjvmSX9tR0fhoYIGRH31GuucaVN9vVkeFrlztdalpPZwRek1hVz/HUaHGDN4znxX1/s2maB8XTwMPXe+kpdHnl66yGuUFzeEcNfbHYaXDfvNu2XeH++LMdBfXHO27tufHg1AcGwpgrobBeuCHZ67euAFeGYSha99ZusDounZNVzgqmIHVAzr8+W3tkDVZ58sYFbkm/hlHRZ6NAaQtn7Q5mg/g4FabWd/xTjYJOV603AMh20N7++r1PKgfjPvcdh3KoJicJ1Bz9FYHD+Ml7JtHgOTIUdHFwaij7SkJelfD71toTp2JdgcDdBIM3nnFFi+xZ2W5WbGf6mzoVKNTw9l/cFI6+TwA6y57/qFfX/RlUKfKbv/GHvLIf7ODNYL2ilNH9/noRGiiQ53nG8LnWUhQllHBdewjUngwIooms97Bawlmglx4hkcNb8ZC+wgqcfHYbm+r07fN+xVljLQkDkBg2s51te5d/13KHDfHxOCocL1u2Gg8kzzDwTHyclSgHO+ASMReRDQ49AIHQQPQ5PjRtyD6IlDHCFDbAGoDwu3RFjW/+mE5KvvOos6RkYlAzbGMpNu88Rx7tpd1jUhqz97yrASM0X7s2eaoQKR/V6TII0qnkQaN/uEP3GrxG9nvjp5whtFuZ5aPbd3El8yhGBkrc4TNp5SfmgHA0s5Pr/YOOHPIIwa+O9j/BX0ivGH1p8+O1Xi5r8/WdBtODA98ZUZXZBLANoBzwspJ0xFQeA97NaAXA3uDsqE1y1/Zfcxi8LJfIeswdwZpoq+EOz4eHrLZtv1tvR7mH/S+NF4B38Cxy3nZs9w54k5F481wqn3+fPkR/Tb4HXvv0K6y+ZJ3MNa+L9RRAXKHLPCyyDjrxkw/OiXoELW/zfGE+2fHl8ooLQ1ofGGYm5du8gOoHBCosFIOH5aw+nz3MGRU4D6UYAJ9KN8h780xYPQF/di8nmcl1kLPWJOdayfkRpQu+rTiyi9Wjuv5KTMjXNaK/Tw+jxiY2lB0nLUyUB8ZFbul+Pj816HAbY6Kf/zXf2lZBRBgPOX66e+ywuXMAXAZhDjrqEjAtL2qUlgpOOCt5kWDVjIpHXvzgAKaG5sZJBCgocgDHWiOCgss8CZRLy9odBXRAnXRoFxf0OiICgjpmvX2lsBYRHRSQVsga2kwaHrcwHwrcBKwJJRwRArRC45DewIWZQxaxgV9OxBFsspsAWewVqSL3hxdAW/8HAePjhdXR3S13yC9SvzJBCeZ2hcHifToIIfCoWIKynN5rGMQu7T8kXPWxpNGz+Jtaz/4z3VUODWgnYGm4b1qToei9jJaJu/zx9RsEdG+apw+Zx01dhOCgVa6R+d9SIh1eP0JR0VwBqcu+lS3kY2/NeKvIvBSyWIGhcsypBnTyGTU1RHYsg8e7mMcFRz+nWv4kxwVKpE5tpSVW1FoM+xprKQPbhnLw5iyqIstoJlEC6JJW496HM/GyVGRhvB8slAEjidOAiV/A0dFbLOcxhKYFdJIVYs5Q1GIwf0CY0D24sDjRXZe8+s7KjjN1VmEvV+gCkRaTXq39yYjiroGNZLI1vP94EDHyszWDfHHHRUmM+c56jumE2V98m/R43OJMsVWML76z6gv9b9XxiNoOO7cv93fBFZ0r5Us2A9Mrx9rVo+jRw3ptiGvT3BFFJF/0/OGXhhnHRU9qEPOYEWafOzMAoIMUeD0Buy4tIYgLQ1130Y7qvwBR4XuGYLN14lfV4x7rsDa3VO2s9i+9lZHhe07ArweNSwlfZabiVmBFmUci3Wt9BPPTgxadevNaFsbIFy/d+YsqugIdeD4izfL2DOy++QC2igYHIfoZyDN8zmHB6YzJJ6vssGdGAH62v2oVQ8gfpQhOn4dKrdURgbH2tmzdk5Y6ou6x+bAApHKLXt/JlRqACHkHJSSbBsQIu5TVk5z38A2RDg7Z8T5ShuINCE97XsrbbSTETgT2DMRzuyjUmbI5ph50HQh6yHoZWvMgSdBZ7S921pggDVV0mP4nPfgjRZI2GnKrAh3MLyEfh8gKXN323sD8/ByPO6cgBOA/evIW3RikM/M2YBSPwAvCR6z39q40rRH7XPtJ+fybMhwGPk+1zT6WtrWoW2r69z2N/nD5UDZd74HB1nwMxwVdLzoWuNcgp0F254NktNCGsRj9Q1kj4W0Ks2eN8A+8AmeA9y7dEhlubGImvcMCuvF4NH0cF6Q/jm+cKB5ZlwA17ZO3tj5DeWdDPvxrAs2D4/SR1Y2jo2muceYWeD9G+x9FtxpThTvp4mIfv7QcbfWl/E+NM0ufdPOF28YHxkb9mz0Q8CPN8GOstfo54k+FfYOODuA5aScjF6io/xQmZH7LkogOc+EUxFbMfQQL6cc2W0sn7ZwEPJ5uo6UVZ8yWxRXaYAKHUheni0baX+6vNkcWGIqcIA8bwwP+vQ5nGBoog5dGYG3dFTY31r9RHUqjG1d+mknS2nfcY7ENMlDfBczcFieepQd9jeDIPz3cNC7M1b00o+MihXlPj77xSiQmkuVPInaam+vz5c3b7TzdHl9fry8PH2//OO/+T0OkAJBVanR0k+2EaEGlUKim1gJccZR4dd4aSkBaS6fLj+e0MyHB7N9bwrBzlFBYZlAmzyvbeAExKrEg92TAGaA5tjzc0YFGiDZgcPyWIpOdU3JjRYpo+UpWhEhsVLQnKrSrNvHRMu8pDlcKRElTi/+aQY0j7KNw5W3OOz5jqBNzsL/tgFVwyJNhS7Hjr49ALSW4hLPcYOadK1GvT2NO9WRNMHEiY5IFhrm8Q51JHi6ZUSz+VhVeFNxj0wSb6g16P7khZUhx8Okg/E192NwyN70M0o/dTAitXMgfQMbXEOZcH0DdnaOitRORmugv6Noow2xlUYFfvVD/RyIsDIKoVTJO+BJzcyJHLpQKCPnUh5ACTJaqKNiN6rRKKq3ixxrY5Ir8vOIZOaekD0eSP9yW2sjaV7QYMl4PtdVlbv+QG023ODA4bIAN0griapRhxmAYXHgHaCcCrbom30eaYyvqZ8SIks/rcjEnU3Zg2sW4jRvPgIkVgDEdD0HFno7gQc9AyAzB3RPhVDsyOTZePEM4PzLcVSA7sf7m5FyPu8DvlE+b8BkLmw1jIbhupKBOpY/7qiY62PTbquzrHHooVhOuEqy9bqB1rl9QddP1VRy3hlrfaUbXh3s3oGaBLJ1yShDlzvynIjPW5UNRrk/ApDQIwPaj/fAfq7a70thKqXEeIj4o7ZOo80kwuBvbK46qNQZp6NiuyfC0IaxDH52QImgd3MgExwcS8tNQY7L6a/4A7q/79pwgvx1HBUqF46A893AS2e/pufkwXqSBnXZH3FUmL3iGTuHss/A3zqbsJek74oDTzjD0saJv3NWwZJjQ1j9njgS7KljR8Whd3LsUTHuuSvyuw5bgFguLzwymsFxR0sUkPRiUWyfu21gtDO5P5QvTqfFptSNvdWi/g0ATcAs6tvvuL85KgYBtRMfR5zq+y6mTwA55akE3iiFRuccap5D5pm9iSjjcg7ovX6tR2hv9Czp9UFZQJtptUq7PQwRO9e/39nluQc4MrHZl++FC2XxVeitbnP3TRbfCLVLXkJvQHQ1ZZRFPRPURiCOlbSBE4vzMNDRgU6PMHfpvT5yaNBGlJnt74yGjlLMLvcD0KeN742wxXFlnz+/AotguaBWtluYjXzijiaHFWpsozOEg8bt5lRYlH7KbIS4WtWKsM/pOAGIimwP1vwHkGw8SuU3ZF6A3OQB0L/6i3hNfgsWZWk36scs0fsGcD7L+njUvz8ty4gjY+Y+cRzyRpYFcydQZS0xsBTZNQDB02EU77c5InMDpf+MdoavmPPC1tHWzsZlzgErY+34zUtUiJC9upd+4CYGlJIv6YxjVgcyVNBn1t9hPSqi747ztfdgKeck18OeBwdIrXX2GsxyR8QeuK8Q5Eb+T6wu9gYzi+i4Unk0zlPPcjwPY4cDQXh1cITa/H1vWhP2KPX9bHuPzmpmy4QN4o4A50WcN7nmogdqNgowH5Qs62t+sLcXiwi5DKcnn2nvp3OKGTi5j3c6Q9g5zBZkNpVmUzhvfGRUHCkSH9/9GhR4h6OCAt/BclMiYzOnGqPCQupE6wE1aGHlqOhqAWhEJcB+D2CRn1uJpTgQSpnBwV1n/yAo0ojDoxNwjgMxH92iVntUPB5BZTiO6RDcLvQv1gTr3pUCglTWswLCel55joHC58uXh8uL1c+LdNLpjjSw493iGee1kNlQbFCrbu3ZXfMhIhmsx4MNGEonazgO6mo6LZCOSoEIZU3LJo0CW8HPWmeNLE8wO3UUGtulGOJOK9ODqDQfK9Ma3cveo1iZUWCHokcx3N1l6qjdz5qAPBgsssB96RYNEdzI9RqVEHWEFF3ng+pWR0VxW1+tHdjhUUax/iQd6TTrxLhiOu9ajwruxEERkJtiRUo9aNGcM9O/z1GxPvQbVeiUWmTnQGmrq6HrMsWWX3SKjZG24ANxVIyI9rCh9o4KXqjybeWcse8xpnTe5a2ukq6C0/yKlaOC9WeTH+JZth5MJ59lQq2fAuFKKb+HPBO8x7t8rf0PKq6Do8Lv3ZjmaQR2HkTdTTGkFgpbrii/M3nQmQXDzncXc2BZa4ZqsJHXRzohFm+f+ZXX8zXqqLAsL8nU43qrcg/+JT/ECsazCD79S3dU1Bw3J9Mug3Dad7FnRHjm2qdTRx2Ai/Jtsv4/o0cFHRVpqAXbr8+NwU/V5pc7yz9V3jyuWjsQaeuoUCE5ytziP+M18uMOxOjjK2D1jzoqKsV/cOflcGGAq6NiZ9Pd5KhIfQe0/MOOit3z4lxpgUDjlrjqqKDMJXAgTVFPOAXXO5CfMsupy/XtCa2CV9nr4CXkKepbh568grcAACAASURBVPQ+eM6f7qjg2HTbsqSO96WzyFuU6uBZv5rOstQGlVITX2wC7O+Zm46DDgR25je0M06i7Hlfaf54KfscLEnfom+rdGUGHoQMxlA3Zz+ERzpeGBm9i0CPHZnD0ce6JMBGd7Aqm7J6o1rrQ9BtnDFiXedoNgLAZ1DE7atsyFtXcmkY2gK/EWL0fSUyO1diLirHfM3RmkEQR4Q7JlVPKoNaniG6T/AKbByUILLfUe4XtfTDuo2IapRjOsoOJmi4dlQUJcCZmx+r++94AgDUBo5K9ofKAbcIw3EDJxP4qZ+Q3FrWs4Df9DF5r7DgkcIPWG8NADr5y/gP4tkirYF/uM3pZWt+YDwGNIujkHS1Z/zwvhRWpjicRRz3sPvd/o9muKbmW79Lt3EdXGUGCxGG2Nv5ORpq0x421fK33/7V5Z/+6b9lL09UPyhcoEWha0aFBPKtzjt89jnUf8UZuOdkvUX2k6fsfgPmDfNAFgNAbZYtYu9OA4apX0vCVgDDWHfrhWBBJ4R5rAQoS+u5Q8ScNtGY2zIe7Hle5unTZy/j5OV1rD/DF3MmWNYbgGM0r0ZEvQfCMsuA+8IcR+HoY6bNjyf0qWBZJ3eKhqwwZ4RhC3aPZU0YL3i/ovs7z8SwZ3gJonAYI7ASzg2UnLI9q7xcNH6NklolE9g0+xmlhaI3kjfTNif526s7Kb5/fwwaQuZa/xI4Skw2oJeSPdObTHNLhf3Ms1r7ufA8gUPP41jjiKM9i7Pozc++z17Kyq77y19+d1FjfDCdOZFtZSxn5ZzQd8Ge84w45hiY8jLPKaMf5+TyOxxiKvvdFR59ZnD8GN2fkcXnMgkBBcYDTQ7JvtMxbx3R7QvKE+BR1YvCsCc7Z1CCyvg0y+xH+Tb4aqKnC0aUUsTnGJkvaAoOfm+q2IejYncafXz+61Agd/WpjIr/+A+/uwD1CHvbDuadDOGLzRmnUAIxHYxWkAWH22zWzICpvynex0hzKAZekxGyvzaoy0B9djguSs2Q6ElxaARoROGkIDQA96hVGGmYGukLhRO6otc0fLWST3eX74/fL9++fYPDIhojhR5FFTNFCz9nTTw2WcXUYRSgbl70S6CgExLaTLN2ZThr6GCAWp1EqF9Failgon4NKgdjdCIWpSshCawxbTNT1UuByQPsbaw9GjyU+KA+PAbqJ1FFciKaRAFe3oNvNH4GvCV8SraRKSByK5S/rHvKaJixjBPSd+1nLm818HYowhW5q4bkCgzCoGw8nvlh6cLB13aAM4qAQ1cjMwtdCYhOJb7WJ+90kpTiwVRwgjB9n85AaJdmZSAoY+aCDqIv9vW4JjHvcg0JGJdp/7XOpBQKVEY0SChWALPJ953OzjeDyGoyrGk+MVbJXk0ARJwCNPBI0FYCaZh9rZ2sRZbn2EWXzzJz/dgAklImF63brlCx4IZ8OHBHWR4vyS2UjYbn8dgjXn3nxTtzAeJaJ9KwFlyH/DgXbUe1fELLWNihkZun2Met3q+veYxu+SxEaeEr9LWpH+co/JmEIu/JnMdbdKs0Z049uWe9jFktur8GukbUkU6fGW7ljOnEWWcX7LMdaAzrUxgld0D2P/QV917+q/zkRlHP59wCyro8IXcIVDRbYuFxBIiMdRVRu4VimoxWa0EocYZ9S98ZSagBGufIm/IqmT6EYgKNtwQ4zO88mk8ZtRsJJpmN1ihxdBaWSbYHv/SeMxTZ8YktszoD/TwNoJEbvhw39kktMIz44hMf08RPVS6Fzynnz0bmB3EVRBt2MkQRxe6G5w6gwy3JjrDl1U1Hjqkz69Jky6ZYPiJUB5vmyCGzoUeCYauBbZbC+WZwOs2ErxJDW5qrLePvV/1r/n10vXcZzL+G+7bz3qzETuXQqIfdrcmj4SQTfcv3QXw/RnrycfnqXFb80vZ16mkFNoNyxQvQf6OMTIDKVcY2ArPEZkrHhpIwfkfdeh0HULja5yMxJPNFv9qIa9efNhtsJ59gtyBoCywEebILUOvtawq+KjvTgFBrpFuampVlSnIM4+sNpwFA7mLjcg6DDMQWKp3xyPmtZNRoY80YYNS6XQuANuzjoDszEXyObp/FT/BTObAP9t1qe9aDmp7rpWeY9Rb0c+BZAvxQicGcEXbt3YjTujgwGj0//Ui9w0sPRalpzBW8AMwCPTz9yFHYN7IIW19I2WO4r3icOpE1GPbyRlEOGs2eAd5y2rRNiffYNdlcOppQW+DmtfM/2JiLAlkYcpYZKiU31B7ETN1JEVUh6EiC8yZ6LQSDup3pz1WpwcyN4jQGNkL/r0wWBpQ+Pj5GHwk4HSi9ZdNUD4LAFji+KlsOnIl4EbMrKmsAjgpzLDz9+JHZUDZ4c8hY5oxNx7MSHIe693m5o+HzZ3fEEJg3R8l3H/P95ffv3y9fo+eFrbuVgXp8/AHMKQJeSeGUTckf0rtM5ILK336SwV5h2SW3msxZ4qWp0DDaswxHGSjnltld5HnngcgMmSSvPcN639wb0I+eMu648Iovo1wObdicZYGzGaSQpdroKFuddTz+I7OCzlOXId4MPXAqZsxmebOL05/9UW2dv3794rQ3erizK0rFNR1KzGOcaxU0Q8cpM7Zs7rb+LtvdCcighk8fGRUbveXj41+KAoNSj5MZ3vpF6af//e//yUdvhys3r21+F9pqfDXtctSKVeudNeCtoyKcAC7QLU3t/t69z4yGAVkXDQURb5+HnSr2I+iKiJvSpJEeCcAP6YiIXkYTm64wqwJpB7cdAtZIybzEdtj4M6JWobIADZz0O2RJFHPEIOLl4eFLNhij8pZpbjlc/OKHnIAOS0fFdILWIU/gBXb1xiLkkg7vtibi3VHBKAfzJpUCmvpgdyPExzv+KEXCh5ZGYfWo0OiQPFTBFgJqBvBCzW3YjzgMOBSNVskP2x0EqxK0nuoSEiXwGLeIlxozGMZ90P/2NRWHIPlIa8yS/9vgFD1TtEI2GVSGI0dFPVH35mzrxvrm5WQOOVEn2cd77N8+Z5hOC+PfIndcsRz5CbPw1P5w5HD/5uxGw2jlqBC+Wopq1FxDJgYYMesc+/VNUasox/FZqoN1OVTNUYXyukInTxCubKetOzMvjN6EYbtZlvyuyczJ+TDfHivRom4gnrkX9u+c+XiDqsTocvxnEN4N5cbGhMfPpKMCdC1HBccZ/5YQwVshUI+np2RRqxInWzwmzh2RaHjuIJRzrkq/Uc4za6QTZueo2JUmgQwc9m+cmSeZ9ebLRkcFqFtjUCNYKbAHerhMdFST3mPgQ1wXZVEUnL4G3jb5uWHrM2x8+J7F1joibhsGBBq7EcZtNz7whpW8BlTomerRkiMQHO/S82t8/c90VIw6n71Ly+gwYlo2PPYsF4xO0ENHBcs4wRGycgLmHIVZOk90WXDdUbFbtJ3s3S/ytT2gdzp4fMsNvPlKmmID7yXTYBr1ZnrvdlToGZe+aumC3d1XayLeSI/bV2ifBXTzs47WQVgwAeEycrqObaDRpqHw6hhjMNGKgAC9AnASZyEBe0ZxM/CMZxfBOw5s4kshjjVI1VJxAE33uWz7zJM1xSnPlt9u+INgdMnMrb8cMqnpGqW7ZPa8R4zDlqx9WuVbRtp3R4Xn7aw0S7+tgM5ZZ9DglrOygXXXqyHzWq54BoRbYVKup2JzQBcddWTk7dZhu1+mNQpdIm5w7FTA8pe35whGsywM9DVocx/3mfdHQC/FdOaw8kHIVAC5qDJgWSSGyeu1MIqBMWSkWlM+4NRxNVQ+Z99NL9MTTMAofe49OMgsY+QeEekvLw4SewaBZSl4Y3AL3gTFZ16qT0qWY6FYISED71oD+85P5hiyBtRal99xmAg6tc8dy4qsAp+TH+JC/+APd/w54I1y2NVQ+dXB9d++/eb0ZQ+IpdUbTiPe6+thb2NpuwjuNJ3C8J2HezRQDsZMnI19Tnx+Np6o9uCZI6+vnjHCPet9MuL5JDVLuXnPlMjSePTm3F/d6eQZJQ8oT+X0eA1HXzSZZ0kr38ehl/F9/AwrK2urGXbae0RKANP5ZXSBnJ51T2QSRfZb8Le/x/tcDLzkf6IaBstJZa8Xd9zV9emnCqcJGo0je0l55MhRbG8znre1szUynkcbd2RKZHZglPuybCk9G22c5lwz2jt2+PWrZNWUM7nbOax4AlzW1ytsR+cFa+bOiiu2fp7FFbiK0fEjo2KvzH5886tQgCdnbNorjor/49/8s3jSkY6EW/icQoRD3C8OIgEYV4ruVCsa19MjDNnDBmgGBGot77OOitjJiZ3JmAzIi6ZHGvHjcxVBaId4Zj+kgwRe4ueXJ/dkG13scGZjpt7cTg/jOIsiWoJOHxNNdviYYkyPez2jhOwouAoP47zsrFkADq05tTp0EBENJ0oAQBmt0zW79u4Al9NRknVp2QCvxmC/IerarbsiRnMgjCFHBUmMjgp9zoj3dXr0tZ6UpDi88hmTQ0PmkAdpGEYtwoBPtusLIETnlrmBaRkDen08I5QnOMoKvO/9S+b1pTKX4PkI9IgiUNEzY0bFqC8QwFup6UOkdwP9a+2K5hqtOxgt7qRQ61BSlPVjcUI6xsbyXVl/GJIIyt74jmh7k0ul/LnYL3wGHRVnECCpm6m8duSomE8HHcs4rp25NN/D1dk5KlagHvlSozmugX9Y6aGUTkNpF7StDZfTVz/bSBPskrjJ/9ms14mjduWIgVhaPZNZa1EyTPkPTDaItHiGf6zjpczP/Kd+Xx1RISH7vqudRnlBPjigA18PqxWjXZzBN1UJDGBoxzsnyP+uSxpo3Ryvg3xK0KrovXph8mwY5owGRPDCsBjpj8TnZ8TAyE47PPLDUVGr03hKCLaSgFspeIagwhA7QxQGbjWfRQALmizyFX0P9BHhuaJ7LDMqSh+i7HNgZXeGcKPmXuZEuiw4y5/rjbij7Obqk5c3J9TNEmAt43bg8k7vXmBkIcFPTmLFNwO/QZcXQCTv2bzjRkfFEel2s7jmrD29HO9xVGSWMs7X5M0RZBJWHiNz40BcDpNznp0V0APpmCBAhFNZgO1QF2n7rJZr56jY0Y026/g9lnpeJWrK57kQdifr5YPnIgBpQ9dZ/Iw2DIBsqFZRRm8TtwY9otdn7+FPfeY5r2EQAJT3mZtHfKkgJ+u42xqymgHK7LxcngzEHWiu7/xrOipwZoTDIMaAnluWNV9ZEFQEHTdw4mIdeIKwNr7NCbQHRc3pQDuOATTmpHizMseZ/RkmpJfXYvDlIE9jU6IsTwHGAIirpwlr6LtjJUZXct3WEn38DLuxZ1nZHQPRLfDy8fG7953QEo65r2NfOEfRUZDOA8zVcB+nSdskg31n5YECf2HPAZZPsnHSiZLZIXfhnNGHht7OqPXM0LByX14m6M4zGwwAtr8dpxFrpA1PHBXZJ4dAf2T90EluY7NIewO7s49CvNMdFN7HFI5Ej5yPd2J+keVyuaSzg2NjkLHtCzgsXr2kmGdffEbjcAfYIxjXMYaoGEKeogylA0j1ntrbIU/S9i7HQILzUSWEza7NyZN86z2AFtm84sSz95IGXprL++jooQz5CucYeJ0OCHdsxNiaLR68TIeG7Sn73hxUutfaewIbo/PRy0LZ2KIhu3Gl90KJiif2r9M/Spyx3BkdSD4va2h+/5C9g/J9aUIWr9sawgFHnkaZPsoMc2bZVI1vnDe9PBoEyoej4uhU+fjuF6FAiBV6O084KuCcqL4FFNw8XAtA6RHwpRxrE9XxgFwpbmHchXphz3eh8fbmtf242XnwuFI1eNl1TEcZFTkHpvUvDmCCw/S0QmijBIg9G3UGcWhRcF2NDIk6clRF6KgwSWPPNQ+op4J6bURGdBfFQ5eEshLeZmWwwtpHA0//FkeFpQpGmhudDul8GDh356hoIHmkSY7x21oeJjRiPD3tbDHsR0VFQPBSBmQ08T3Xu0BNAHtU5ueNGE9rwGqjZi9BEZ555bl+wPbG2DjsJKI931PlpSbQNaJhCJ65buuHGU2aWse0i8UgTP5TI1GZRqKc+Gwq1N3urve0aAk5RblbqwwC7+FYlZZ7R4VrqP41DSh5N5fIH5V1ekIptkZmiHpBzVJ5x2idSckrBaWVp0f+0BRx7PlJW+bG7Kk8w4NucVSo4bkC5OcI+L6vRwcNHRUd6GePhD7QUXZdc1JwxRqpYe3Kg5Xw8fFwzTVwLXZx0Dq5romPeW+vP5llBK9bAWIovefnjWqDKbQac9a8w+Ahy+ZI1JLR16m184cyKpS+BAEKPPvZjgoFIM/wytk1mvbh6HQVeaYg1AgSHkVEucyzpnzSIHMHqgwHVYBgjR0Pp/ZHHBVHD96BW7u1aOn13IPz5n3vMi2BuHrYerRcozpHh3aj420LcfLeAR85KgroxJlynBGympts8G3pJ0YLVpPLs46KOopSgYK4ide+DwPfcdRGlp64vAEb7xiUFaNY/WQZkAl3W8nxPWuudZtjjjrcd/9CHBU7X/9WVjkPr2nrwF72fQhQaDjTWiDA7iVpogqFx+fI0ozr0BwWcZ+f3KLYemQz3x8Azp/tqKAedVaOMaMC+716gu1Kah36mNIhi4CGyjDalwFURwXGTq/GLKxbYKOu3WYTbc/sWDNiEvYom6+W+6kSRRZJ/NyDnwLk/1s5KjLmYQqQDIkTfAgHAM4XkKTvMc+SsEbP1k8kHmpAqM+VYi2i9TOaXvpx4vASF5mUvc79khgIHBXcI8ZbzEig897GmGXUXHfiooJfPEr/BUGbBtB6lQkD9zdiucZWg3QujL4gThE6KtpG6Q/0zA4rgWRVPz5/Qi+WAHXpTeC8POPq88X7AHjAW8ojsTsdWI+yTgFOm4OJJZUMoEYGx8u29FNj8dhbXtrHy3khE0J7WXh2BLGkyA50YN8cMC/P+R7DxNhPwzMBwolBZ4eXMgqHRsuoiPJuzIKp96OstctwM8WjGsjrc/Ro1LKcsdwSi4FP9Nwb+oVxr5pT0Uqkf/3yFWWuoy8r5jALBOdvkUmZmWTrMl4P4xyll1j5IJqEw1H0GjxVQshKjDrob468wFjc+SOlzUaZzKBlL10V1VOYTeQZS4JDTCVpI6ASgdDDXgtnkdGkgqI13g19cWy8LH/nzjcGtMZZQDlh13hGmZWUi58PR8XZE/bjuj+RAqkFnupR8R/+/r97qhma0KDmWUZd+CxEkUn8sB82GVW2OICXHwXAg2ZG1gD51bMVWJ9OyzC5E4HRJHLQTM4TOc8IccFjjpp1trHTIcOU5MB2KMDcE82IBK+pZyVpmCIHYepgfTSHUsdFRWHGQHrQFSRRLA2MVERiULnGISTCVe3fncXkS6MX8m+bc+/5YNch7VNqcIfQm0A9Lpo1sHKawxqAZzzA93RU9EFX+nSKzR7dRIMieAk1BTWqcXR9kJ47DYicUOD2uPnWAZha6mtU1qHIl1E2RCnH3NMwsvJY7PSVw4xavU6/2RhgCi/d4FRIAcLXXBsgkeXYYl1YOmME+OjQEUONVFLjrYH3K2Ao+a6isLqCTcelUrx5CvpSmHbkGRXF0DnE4K2SF4xugbJnyplHA7kSYIcy5dyIYAx7IoC6HfdwX9JOTlAWWpnAycWXphqsf+Z1qxgI3LEGF+fRrcdLnsKzSDtkOhRNc0cMjJ/KYMxq56jcHV4eDcWBMStrdFbEzbMpuwtJGnhnBVZfgUavHraNmCvK6uERv4dCHJSOxSuZluyxyKjYOcVGoCT3ZJquQtwyT7fAkZ6tzbk8IBa6tSZabcAk53xJ4b5K459wge6NvmQ80bUefG2Abe1vmDSIMnJvbcgGHLyLngLzJCAv5zJYq+n+io4KUm5yKrYJ7BSM/aLeegf1GwNsGPn1HpZ5D+A8hGjma12Xi0VTZ9wts2ZjQ8iDUbaAStC5qtwKy0AseYhlEHGjOPVJ8VhRiqmDhVjpPZju7qb1qXMUlLMOetjU7z9c8Ovv5vYdhPHw1M3cbvsYonU6CuIhFSW0Oe36kK4GNS3ostITsHTriexW9PDdW97ZrEUASqDNmtdP7ekpC/a6NBmv0Hmt9BjtVcEjeuJ9eWjbx8w0lwbOp8/Ng/11fZb6FnMLLO6wvgvXHIELfccCqew22sB0QpTt3jPd1dHjgC8B5eW75VxeBA7RZiT9efyuz1DMmbLZQbqMnga4x96BAMsNsK4nYdyVqQBppzZyxlzPr9dKEpNUWWq04VTwEXdbPgISmcGQPVDyMX3/APt4zobOpAGdMijfzRwHCCcPopSy0IZLOK0MgI5ytsqO+CjoSzxAbMRseh31/tmg3ntbZJAYAFFEkMOx4qWj7h+cytYAeXcKxmEIyjKQ1oP7pbz0FHHfn2ajR3Ni9JFEdgdKXRktUBLIeATVL6wE1+x3hbZsU0dwKhwfjFGy6X/9+tV7CTiYzKyKoFXjhLDBMQdkQ1DPr6bdaNRMBxP6G/T+qE5DL6P1UqC0GP8I5DWnC3jEI/u9OfkdrNSI9jdg3a6xz1COC6B6ZmT4WlYWjdEQjbSrogkygrBG6hQd540gjziNB8eXZxdEWSLP5ggZsu/TgxLs9qPOF5R1q2MPwwqdPvjI9g540XrD1B4pXuf9b5e74C/N1FjJZQaHsieOOeLsd+tZYr+jhLsENWoQafS3tOdqg3WcmUFnz4rylQsCFpv6Po3A7NQb6emLyyFXwlljzg+WfrLnf5R+OqWGfFz0p1Igtt3JjIp//J9+b6OFbJwjwSkzu35aDQUlZH6e/fLkqqZrdAA48G8CWK4/5aiAHlU/MUg2z3l+soY7d1n/kamCdMx4cyH3qr9crMYcUwqZ+mcHIGse+uHj3lhp8hdv7gqz9lnAwfjqSiYaIJniYmlb9mPPtiFTQBeNOasuSvNwWIYvMCp/NCYQkwoto4AfyPr+fAXQqilVOSqE0PmrOlzkFQkIqYLU0sND2cI9fVwlwffjbVkVG0vAmg35T1Oy9820DfRlVAujEdgkKhV7jtX5AA6gNm93TviqLx0V2GNVaqzSnCc2rqEPtR9ZMmoH8JEcNgoeqnC+KOKsB+TaQK1smMgkiSFin64VeHw8PM8dFQHyq9Ln0R0VEaDGk70DjgpLiYaSRQUahBnfMRgAay+VCouMRCKdOCs+aTTKn+mUGiRdW4ccRmh8lBHC47XvZrqvV2J2VMx8t3aGqJOCwO3aaTJMSv6EQqykc4p1Wg7XNy5oXrfFewRRL/LB43ubkb8ekkjAceVS1HTHL99KucnbYnTK40KG0VGRstGja2R/xx+zo5h01R080mtUcuvBY0aF2x27rf2LOiom6SGO8cYN0iBy4qgw5hlpl+t/xVGhoHU5KnaRp8WZf9xRsV6kHffv9u8MZIGfkgdWgPqGP1bSwGZ8DSsb75scFcPRMb7+eL/fJg12wJ46KnAkHoOA0FP1fAZd8/lXyp6yrAb13TVtI7NDJV6rbx66EEXQASn+2o6KtZMCC3srf+xOHYI+KlOvrdP+BFtTfDVWddIq/3DtroLFeg6+gxh/dUfFjm8O9CUFr9v4hmetA58GvUHuOXO6j8Ml/RN2VrBTezAw6pw11HUt5KF7R8WGUAeg9paXt4y5fgeB5eI11Tvmh4lGEKBrCSuPCH97Q/li16Oj72GqNCFXIAgTCM1MlUDudms1jTGeyzOXvNMcTFd4TSscMKOCtfwpAxTwxSsD0G/8JUI713+muTs4tnt1befATqySWkbjl+fnAMuRHVHzEOB3dNZ9vlx+PD9d7iL6nlUeHJhmF0SWafK69WiybO+yH8MtbBzu7Eiwv5+q2WsgyrMRqOcyeOaKg9to1E0HgpYj9ulaxoFFmv94gqMg7nv48nB5/vG44fJuBzmZQ83NjIg8gwc9u8lSNCo2cJ14CUB2nJuMsie24h8PykXpd+hHhTkjwt5+Hs3eNGfI85OX6mFZpuRhnSEdFRE5b2C5PdOwJPKm7QFmPDiHRnkktcPI19os3nGoT9bX4t4bl5uzwhqfe8+EKDFka+Bb1prKe+UPc9Agc8Guc2eel0fC3HxMRjvL4IjSRyj3hEbURhtv3Bx6jfOC0l/FeGQIIbAZjjPiJt40+sePwHTKebN0VFB2R89aBn2y9JO/fzwvAkZwFjJHxdMzeo2MtmLsZ1QxAd7G7CHidas9706Azxbc/Mmbk9u1Ti8pL6ZnIMpPwXkEen8Oh2E0+X5BM3U6XSFOZ/vOPvfsCesH40HacZ33wEHJUM2ycUdaBFRzh304KrYH7ccXvw4FgvlvdFTQQQE9pVLU8Td7V/TUzxlQdzEwkALR6Xn0+A5VUCU8oBktDoGJH1UOELFgAtA2u39Lw7Ft+np9Og48u4CKWAlUGh10OiSYLgrUKMTcgNEo2j5EFeOh8FXzHktvB2g01ubHQzzlLQ5wlKoIrz+jJgagEJknQSkK6BCwvm6xFvBAD/Xlh8PWHuOHqR2wJiQj5c1yOfWg4thLSHctINODhYZ+iGXpro6agTsgxPNJBv5nyhyUD3svU2PXqCWiANpoYwzeUCv7clQ0RfHkyLN2cNthYXzPSMjycmv0DLQEh9D72lMLK84/lRVfY8rfktfTEBkUfKdb8ncNY2uLboRVtFmTcY7w0by3c4/mmNQoGDVEOCpGoIF1Jhka5Y8KGeFUDd7N6AIxKJqjapIZOtFeGiC/kRTpkYYjWDBKpRmo2QmD/Uqo3G2jFb0eCmDREnMW4JGyIy4ZgfImeylZD8CTLQAa99ZSh6WRVkdnLGRg6L5eoGujsZq6m853PAnqdHAjpUWljDzbx7ReiSbhumHjc4u7SkANe72/YwWqIVtPzg65ZW0ck1+DxkJ7H02Oi9FP4Ac4JGcajDWc+fp8d5PXBzHXB+CCUiFr30qEFMTU8fqseLXIXme4iFUxQCo4wIEYDwiY35c8sACWd0AFIlG1/xJro193YGzE7emPm1Q5Qb9bHRVdPxvOjz1Od3r8HHd1/gAAIABJREFUdmE2t58CEkpf1QdqFgLZ/Vqj7t2AlnWRfQsdFGhfPGxN+vOOivGRLPNY5xqkWW5vOc/O7BuI9L5gpfbJgbKQD0eLOTpoKCCRfWyAETNGKnJxEcZ6yC+j80adhbcw2i0OBH+ukuWEs+oanVbfn1m7kfdv9czvIlW3493t64xIrQh7glA3JuLsD5EN/9VZNJ8TPeoaeyTtpWGSri9F1jsDyxhoJltKyh+REWZqEThMfiQRjui39VivV2N3efX7y1MxWLbK9mT1AxqLt2wWlvdxWlm9ddDUI7FfrN69BdCFfAtAloBr7lcvUWJnregpDVTcD2i3V2/+XGwvOpwcMHSwGJUUvOxMNDSGjgQecZk+0E7fv3ZepCWWWSqIGofdjABIRFxXBgvAdPSlnPntxTJeLtbz4cE5jGVfNKOClAR5LVtg7ovo3/i8SvexZ9l/GBsAdPTdRINlqJJVPaH4kRnzg43vfY5NPnA+pXHeGWDeyhdHhks2aC6h6+tzXxkBOPcQjGbMaE4Ci2B3JIPYhPWPeIYjwcZvYK45SAywb3pM2gRAGKzcUmaIvL45jmTPJUhvDp9v3755BLy93nGmISDVvrOeHDZG+932DLMGDJQ35wmbodvrvQTS98fLt69f3elh72dmDLIrQEeU9kamCPnSgfIIsPSeFrYvY03tXu8/cXeP/iCWzRJgvT0I2QufYs7RsyQCYtkbI23q4BdUtohzPJo30zGTuhvLobOcGQCXLE+Wjd4jq4U6OII8UbqKMoXlr7RqCR1OLoek1BW4XfTEoZBDkxefLt6zBv1rory6425llY09XxCMC12AVzHjAs4fZNzwXwY2+xnEKjSUnZ5FAgel0dr3XDicsPZwrOReptMq9rx9bnsSY0fJO6exYZ40n6O/CNfLaGjBk7ZH3LH5kVFx4yn4cfmfQIHa0AlQR1ra2+vz5c1r4D1dXp8fLy9P3y//8R+QUTECvEhVi5S/jMhOM6rm5ZtHAZjhUEMcNN4R1wayi+NWakjnRlxqxBCK7v1+pmIEAQZbY9Yca04cE8E9rV/q7oPyBqdA4z09Oqw5KsbVbVOvuoQuSL1kFMbpwjlBkhq3Czevp12gKhWllVNo6LsoZQwY+T5H5+1gIgeLozkQD0l4oIWu0OqCX2ZliwoULqHjAL+XowJeYl4CDzjA63oilGM/+KQZOSNTbnVUvL69RO15cgTBAJb0GKnCDImILpgaz9X1ruP6wAeQmrRyZZJglhp/Z0SDHGihParRW+ryz3FUtB00On0mxwv3XHeAEUSH7Bno6jRCtA6UC+wRlpvL9S+iwmm5cFSkZpFGb+32rSxYMb/LH+W9mZajZOHf854ceKDUkc1iUx7NAxPpI9GpcX3UkVbgTI3aM44KGgWTCDsBhOr+jpCPOWwpHuyrfPDMkZ8re0f22OSyxsNHfp3OsQXV1/iC0r+XQCiHgE5xuF7es5KObgd6lFp30uLcWp1dECqgTclcnqHAI3FnCtMo9bd2VKxcF0E/WqV/0FGxcvIT5FBD4ixop9cltdsYaw3GsokJam1KVyUPLIt6bzhEGi8T3YSh8Os5KuZw9s5DM4hcwSQZ3BEbbCVL8dVOk1iLOl0jDRrh1dMJ7FlrQV94rqVsxeodw75tl6zHeoujAmNe8cb7HRUAAlC+gj8Zvxj7crE9t4pDd1TUCUKn9oFv+lAZ8ZIWCxlOEG1y6L/jRd2hguG8E3s9o1i1a7p86mUmbnnY3klyxJurQ2otg9af4v6f5qjgwRrsU+fZThIcUGjJB6MsqvthJ4UtKuzLzIIsc5O6hRbl74ewW6TBswaKGahHwK0wLwG/NtNIHrfoVo3W3fD47ay/p+uu9BOO/5CHesbd/nL0TJDgNux1Vg0oOwm6OjTLyvzH94wSjl2bcjJU/CVlKfvmL/fZWDtKGfjOH0b/j84AZhMAKIT+FOxWKiz9lil0K5q5HXcw+Kh9uQ3D4Emz7VHOGg6BPq4CxocYzMvrJzQJJ3DNiGp1CPFZtLPXe76cMLSdeZ/tA3uvAa5eJur1xaP1lTYFCO+oXdHxhpxkPwEjahDUwXBRl8FfUVo8zEXoqRd3ttDWr8bOCkwHFuC6s5UpenX6GhBNG9LOT23aXDxl90RQq5TvZNkcYDH33kvh9++/R8kmyCcHfc25wcoZDI4L0NjGz/4FiUvEi+07Oh98r/i4o7RTOD8oV9CHxJprs/QSHWjh5DKH1Is5viTKPvZg9jKI/hn2t5dIfnl1ulpw1MOdOWQQlFF7FxGw6Xx14FtsCZEvBNaztDVlL4Cpwm3CVmEPDHcKOaYE+97Lhwm2pT0XyOPcL8aXTcbowce9ufjMPrp7sEyORy8P/er9OC7u1CLGwIwb6BeQX7QXEDDSs4VRAQXZNVby6fHxh9/jOptc69ohMZroMeGZR1aOyktrmSMq+rvYesYzmNkGrCtsOvYeMcenl3GLzB9r7h7Nxu0zZiKR31gV5sNRcaCTfHz1q1CglK8zjor/9A/f28CpmAJkwIEMfCU2tSsFJSUKTOFjulEIc3M0dEpZVYAjozcmu1K0Ztu0L5Z6GF5LB7Q3tM9h9gcWUBoRvyFweDSzFwOeiodkC4LBYOsOnhoHDFAIFh7aKPNYPSLWo9Z6xnj/bKySHt104cGN52pE7sbG1oPVI0CQrmbRBWk00IGQ81ZaLgCA6ev4gEP1NFmhk3NH71HBC9DsCE4wF8Y2RjcYVpQLzm3rw8MEh7xzHbNQ2jOGeRigzr4Zm4yKrgyFo2J8d5R3UrCRb7oO2HE+wYUc71ALcWSOxYpMxNoB2U01lbl4hIazYj2dAOvb1BshjJuNo4KR3R5dwUwtB3LJjHiP7xt/FJSckkHs7RLXv1Xdt4z8u1kU95JWvnukUdlUN6cRWf9QpqrPr2P/q1VbGWx0bJhrtcvbsZl2KqFivF7nuXOEy+dwYhs5m/w0yUx5j3znjxE+1xmuKbvwhV0BUNdgzyC02pKG8giRKky6+p07PYwremTFyBnPiz345Nb0TY4KH2JEQy02/ea4iRGcdFSc45A4geKZP81RgY0pnB+yhsIj+TGiA/3reW8lzf8/66gYV2mkwfi3UUQFsN4/cyg+Qf+u8z/z1S3zaHiQG6qu2yGb0kWDGMbjeyE7Nrt7I4ATuDyYRJeZq+druaiDjMPhHanrUqJkI8v+DAWOztM6Hyqoe6x5ROPd8iyAl3pH7TsY95WBjevOaCHXePSWER7z67UnqYOn7B7J1Lv2AH5/24bYPnXvHNwPZPvq9wLqCxGxhy7X49o7brTMZ93L56ezNP0QkOcIShP98mBdMjAq6n1nk+LNPbuxIio4bClWKTjih3fwAEG59lgvvbPYSnFmIagt9A3amIm8DwPcjMkpmpHuCI4YnbcpV2OfUy6bQGAzWgNG09ZtNgIB0N0ZMhMyHTArGm/mYcAmv2KQH7EL71XiyfExXs6RUeELHaVJE4KPyzMEcg8gfA0OIDQWx3sfRGkmd+gs7WiAjpZVgUh//DCLwHlT9jHexAyIWY5mFoYHyGGNAabDUeIAdzQ5tjHCvounxjT27rPe27HwG8NjDIBFn9Nxr7K8EssemZw1WvwIrMHPkegH4bOLrIUvX75G1oNFlzP7A7RNJ2JkRqyOHR9P7AvKAMtQ8DX5/PnyJFkQnItLmU/h/GAQQdCFa+LVHSzjSLIP0A8CmRS+9uyFGjxin//l99+zPJU9kvxAx4c5qyxThBkUKO0T5+tL2MHelwPOi2XWsGfHvKJklfewAKZkv7sTzegRjhEH28m7MVfghgW8M7OkjcXuD13CMwYyI8RKNVv2CBxTdKZA16JNX3LL7oMzB6WOyKt1pIozWveA7Le8Fp65y8trOKaDD81a9qoa0WfVLbq2n7C4OHei1HDsGbuOfVh+++23y/fv3yF3C8iJuD2cTKqH4jqUajKagMdZossy2Ky3BrA29N2JcUXwKx0ncHqFo86y14LWkAJYW5b3Mt7+cFQcHdAf3/0iFMiTJlJbccj5IbLIqPjPg6OCRsYPEzaf0Liq1yiE68E3djt0c+c2OhiQOQGgfnt4LyG/UmC7EJUIs4BrWxkkaxxjzZsQURClZHZmc7yrj7dHEGIedfB3ZYIH+Nr42jkqTI5q+QsX8n6gupicACgQrehKz245NkhWGYfX/B+dEGPvhWHcS2XPUhlRVxMNnaDU+CHS0kuvAR6iWAuo5wByesIlq8AF8qppHG72RlFBKgeOvXHa7Y6KpKsoHd1+Cy4LPvAeFQbcBGBea0EwRMAyB9Q5SGV9OlfA4GPG0s5Z0J4g5M7xaimdOKj05DwDEWwdFZub01ExaILIO5FDHptMWHm2drl8SIeMknKDRZbA1Cc7oKuoFkGQ0EfaHjprwM5CGhaFjrScsiyESSkUUxPezl05lZ+rJy5byTSDeyb8bt8zYwXvrfu09JiCa+8BiY8OsgbcXXNUbPipffwHHRWjE2nix2Eya1u3rX7H2Rjl0sg9XC/vIDepA56iXY03Lt9+PBTseGLjMz8q5BzxS4NHfyFHxYqPzjrL9LolG9GBTmewAgkhLHeFfZLmS0fFmvsBYP7LKP00q0LXzm3oUaNMUZ1EqQL63eqoWEleaVI+bISMLgvQYCfTjmTVte+2gPDSuWs0XHFUAHyIkVtIm80OlwwdzA373fqYrX5uyf6AbOE5DOM9nfgRSXyNNm29N44KZLwgcAAlNADaUV+65R2jXNjg67c88uS1DAgo3ZuOizM6WnvJeqlPjqMu+zMdFWBF0St0Ibbzu23ibxZcsvhp52Mcf6QFwSUNwCAAud4v4M27T1a3HIAZa5Tz7O08vp6D62EacHDGPXsbORpoxjGF1TlInNKtCSYmPQAD7nlt8RWeET3fvBQSAEMXH3Gu8jb/1KsClE7s7w5AU7GAzjKvU2K1v2DTd+w9jgo2TscQq1QvouIRrU4cA9H0+Gz82TvWoqTmJJQA/I/lkMmXRl97/ycv44OS1daD4q3124LkR4x1gaJWWohlcUDnGm/xxjgHrJ29//7uwWlhQCgBfYt2Rxlk63tgJaasnwbKIs+0YFYDsQpeoYFinH/ZumgEXGWNfDwByKP3RaxP/M5o9gxCCJ4y/MGi1+moYBkclO+K7IxohJ1ygyoz7WIwss/Z5m4Nsu05RpOH+y+X74/fL7/99q98YvYZ+ccdDOGosGh8Yiw+xnQa4Bobp/GSr9f9Pd7x8oJG3J+Q4fD43SL8P2WpJmR3xX4LjMVlVTgSnGcYWBnlwzwjIfpeeL+WyEQhH7sGF5kI6I+A8m22j73c2OVyuWfUvtFYHBX2u6/YyAjki+iPkLLJQfyXy/0nlIYjz9k76KQgIA/9ANk7GHd3jiY/MHOEDcnDWSJDwPpkSfsemEKcCFkG1n8D5ZMI6TDDxfda9jOqBuKE5EpPwj4i39nvtraPPx6bM0Jp5jip9hOLuVtWC/mLjiEbH/cn+QpTBn+7GhiyFWXbrMxYZGu5YwM4GDNTjPbM5vpwVOyPwY9vfhkKxOF1skfFf/m3aH7kd8Vh6PCgbQb35lZdvTIexcD0u1Xx7Kdec1SIElRCr5SLFHjxCOjMfF7V5TS8gDUE6eSYDbkQoB6Fw4jpGhsjkDV7oveIGE9vRpVj5EtATG5xMJUpYKSlG6fVgLzOBUilAieZglZCvdiLxCFQVQqE0hSH7lCje6vHIlsBDimMxVMSPUVtBjDKgJs1HAftc/362uHR2isAVMyo/FRe8QbUlMSs4DWOMS7nEQp2O2zpFKlDOHW+9ow+JpRxCg8aHWoS1EKlPekdClGuRAIP9Nw7J+cS0hQ4EhmjzvAeR8XNhrbyrwzumqMi3wPCcIO0OfNxzIbOCCQ3fqqESin94c77hIwbOCeoFKlO1ff2PhJodEfUBFexk+4YiyiQLodoVJDf5DnNkJH1XlZ+QIp2cPeCFQI4yc0UPESNLD4nn1Qd0UH+LkG348PqFJisa40dOj90AR6PZk8DRSBYueHbftHtmm+y5/OPPPYGug2jWotAHfsfL/3kym4Ywq0eKUEPEdn78UAOM0ejZIue1fF9yFXISZM581p8aqXpFusva8U3r7hkxxtHRr4+5xRvtXO/L3GbmYKxi8H+/9VRsZb7Gvk/8gfPu9U+XgA6TuvbHBXJXhIg5/mSuYbHMomBLS4ifhKKfc1RobonRrdxVOSYVgDsmgvZWBt7ttbjRcjNdXRcgQDhEZl2iJM2u1wAdNcov8+o4GDrHHPg5h3OEJz7NfmftMTXphZ6dx08dLy4E2Z1ph09catfnxiGXPIeR8XuDbu9sqOvOiravYdzu23iO0fF6sBXR4XO0Xlss0YEx1xKmYMiomnZsFaXlWu8za5ShSVs6qtBMbeR4/2OCilvhdKSB3y2GBPpRxq5o1HKE2hfIcpdBIqN2phqDNU3EbvqNkeF37ORUUe6PR2l6qhAA261oQGsuxwfHCzK6wmaBzn3500FBY5y3MoNv4S+B/luNKtSSaO+7M1+w4lggLSBqQBb4/y40VHBoEgG96HWPfp2IFMRZ9XOUYHTjkbvoB8LXUCriIQXIF/p4dwSYLWB9P7eKIFEvkqOiowXNIKOIL8oyWM0sabJFqTKzAyjG4F9f7BmPfnehZxATwf0w/AG2s4bsCutv4SVkmIfG5hYAPjN+WCz92sDTLfX2PX2+aM1uY4yUfzcS/1IppI/J97nz7U+AtEUmdH6bP7NAFEvbWV9ROxaaeDsXBTZ/vb7t29fLz8ef6BsmPRks/GyRBalgjstPOujykthcizNBHMj8Y3gOc0isbU2OnpPjMenFihrPOX85iWLkL3hdnQEMbjzIp4JPKcadXtWVPRr8EyVLLfN0l0JUmI6qXqIzmC0sYogkeFBuqPRNTJ0sf4ItmYvj5JzgS/Ew41XrUeKOQkYbKvnEZ1J9kxid7yOOh32G8al+oRnm0RDdDpHDG/zZxqdOMFwRrAXimfS0FFhc4msHd7n+/mjR8VtCtfH1X8GBRKxOZVRQUcFDwzKAI/BCqWFQtq70C+jNq44KuScW4G0/q6IBGWKb5bqEUdFKZPwPlsNQXemtGjHFc0D5GOkiDsFqm+GNuDKOqhRK5XAtjdCWh2E+rqOokT0fylKOLBpmCrQCUWG4C0OJhyoLJGTh428w4UmAShxACi472tYaOaGIfF+PzxCyNtB6V7gAZBM4znDxHXSPTtCAezSswbzj73VW4QNIkjUUeGREd48a502joktGiY3HSv+YH1S4a0EC/wSi5YAotIiBvxvLROEVEGoQnVg4h5dqPi9Abd62nYLY4034A3zs+O96QSsJd4Z2luDJh0BeCZnpMaLu/pN+RtbUOQUFvPOIeGJnoLs/qzi86r13ptEGxm1rBH3kM6S2lWZS2JdFoayBR5wyUoyBVeRtvEvZJRAyDFlrRlL5SOj8Q6PgtnCVHJiHYPX1PEgPHYNdPMZHlqyQtFr15GdY1xFjT5JGkNMi0KW0kCINOIiHjDXq2hS68pdHs9gTVE+UoyUHe+vMYQmJP54RsWbpMdLA+2xxrZH12z5YhhTOJD9rItoo3RkCIGurbHsjGGx9vRuR9w13rgCJF8bX51zfTxbaRkH9MRWG1hZn7MO9VwvSNcxQHAa6es79it7KAoWX+qTztDvdkdFZcnODsd5HiHF84zgSilvjb+jTEjpppjmOUfFCBzdSr/d9fsVahSX2/eOCkxnluOa6TbuI0YPF7hm+l7JNpxKeOapjAqJ1OU9cPCnB3NXHeuQpDtHBfZAyOTUHXaZOftXuL/Zwa4S5O91VJwQT20grsf4y0ILyJK373BUHDLa0e7oO+gIkL1VqrzXUZH3KTg/sze95puZr27YVmgTlEwAR5uw2xr95OLeWb24dHZEuzsArxkVor/4r1nmU5TFlRz20jb7gBdINICAf/SHT9ARUU9VJw3nynJDpcUWvUpfmEdl97PGP4ITe5Q0yMPSbi8ewGZEQFAfhIvX8ZcAPO4ljHfofBtD8O8Wm9x34o2OCg8IfEGzXq4nx0MqeLCiBT29GC9gECkb4/eRTvCdSuNyRT/iwQ6Cch6YFPgporHv72Gv/vjxFM2S1xCK0dgbLnsz3s/+r4GS3jDaaV48BSB9X4mAPQGMFgb427+MNHedMxqLQ1Zutete68BfLzoZgWSxkT26O/1Y0dA7pmvvZK8YexJLJyVwHXxmfAwQ986xncfHJ89KsAwQZoc8PHy5/Hi0yHbsayt3kyWzJEDXhuw88RkOS8t6MJDdslvMOWE9B+yZRmeLlrfPUBYL5xHHCwfFy+XOe7dETw0/tDA5ZqzYPrJnIegT606g3iLgLUPkt9++ZZ8D7L3KDjE55/xkFS28j4g5Gyw7wJ5lz46S3KFjZ8kxa9wdDZzdsfH5c0TXm5Mjeh+Ec8qBbS17ZnPwjIooGxu4F+VY9i+hvRtl5hyfsQohnulh2SjgW19bayx/FwGIgRmauDDa2f+8+XdkrLjTLA5t4gwMGPYx5N4SmTqKV9kb1lTafujMYbkvyEwXLi5fjHbumHLcDU4o2OrAnmwMxhO//+V35y17Dp0WbGyNUljYmygxh1Jc6gj0pusX9DPxzJZwQKKPDTL92MeDzeFtnNZjxGUB+SN7WkQ2izn8AiOkbPCMi9ePZtp/9Oz9uP9vQoHYxWczKv4delSMBnCr+CPj1oh5fvz22kEVPsv3vKiY9flCgZV6pFtjXA3B4RHXVUNtXCsCcFqTLBAX6XcwsL3hUaa2W1ri4+Xrl28lSKWpmUczvCEqgkaozykBzo0Cv+EPKoqe/RER6K5wTIpeqKlprSENP38kmrG9isYIDV25BwayZtCUMMchDCOaziYTtnZgQ4hXbemdweR04SBzPojKQX1DPN+jKKJupR2COjEa86jTh5qO0ETjnygx1fhKCPOp9c0I7QPa4CJKSZU1UpHjIYBFoNIMJRwofle+pxxleMK19/B53VgjX2CuPRKcfLdiqa3xKhePHFq0q29Y+okHfJZM05rVdEISwHTrgLPu/SXq9eoQ7eWXipcJjzsKEw47gN0uo6K5sCrXmPc0s+bAaL4kESrnABDX+jLOL7Z8KLTxMMoJ7sXks5hHKGdd1AnNs8eNq4bF5Lyk6XNlLISQl622lkEtIkn5YWpMXPcnWUPYe91UT4nWfkZqEK1+R/1SU3+xI+ongQd+3hxqatLLmA5k6fRVAxhHuvAEAwjBvZb7a2oYjzlMwKLyXvI/ZvoWDf+OI3hJM6VdAJAJJogRLNNQOVHG6UiF/vZ2tAjzsy61WvkJGvGdG9YKSZcv3suYYZcODtS8bzo3+pyWzUizQMZKFmyYJj7WKDkXuZO3tt/fgWhy9U5TWTjZ5b2rke30pL0upN8oP81S8YgSBZSVo23FnY1ThdxYvwMmwSaLIRRd9pGtsS0P3H7HK3v2W8ro8fojfRLXYq20fNj6nRqswuwErfVczyrdOp8k/Secuuuag16KZPVzq3NA10PligL/DDjKFd2Bk3U8ij4UfcmSdtq/bZcvtabrzdkR4oSZn1i8ye/yrG/SrWyxYvfgAaBhF8904xkSvzeHnp7rARKR7gXIswRX0Sfl04a1taa+XqJ6zihftGwtAst2fI9Bwy5AoFTJglH3rbcz813H4xR0vcDWW/s2Uf6+T45DJ8c4AcZBm8XrqoiSX5HnTOG6Oxm7DxgpkedAZDSZLb4Je0Po6lH10QgWZYyinrmViHHdCgCY8QOicX027uz0Xg3R0LYC/HbNHBdM4vopAksyYDEzyqKcXEY9d/twdkjvdlBTVikofb09Mph9JQJ4NEDa7HCC9w5Oh32Ye4LAeESNGw0NJLZ7H758cboYHVenD0ZDfqo97vR1HomtKr87D0k5Glun+y8PAaQXj2K7R4ClBwAClDbwmRktFh3/z//9ny/fvn3zUszfvn69/OX3v1zurIxTOMHK1/+WJYcDZpaoF2SDewPn+we/00p5W/Ahmjrf++8Gaj/9sNr5tT7lc7GI87mKgWUYMEvDoAFGyzNC3HAPdxwZ+B1ALJpOIzNAS+lAj6jm34jCB7jOc87Glg4byRjAOIt/6Ij8/MkcEcBn7Dl39/GswCJsDAYSm6PD5uLOOcsQiLI6xHjw+MgWoU3mADfKdyPbwpwKKJ/1+R5zNtp+sfX//nR5NtCYIFhIF2BDoC1/ciphwltjcLfuomG3ydFdRiUzM+2eL7Gm3As2L8djrBfIjyd3eHjj9yeUuTJnkPfCMJ69f/D+C7a/zIGTmR/puGf/O5QzM9LbPLGXPl2+Pz5eHh64H2HjQz8Ou4m1jEQXii+rIbs7d8A3lLtt3rLmXu0joARgSNy6kJM2FvsczicJblWHH6T/MnjDaW6l2u7vcs+AJyFLKEBsD5szwmhm/4Ku0fQ6sh0UN4wDJrBEe3Zl1zADxdbl99//4uP/u7/7O9+nNg86oHzUbL7OslrmYA6G+sioWJxnHx/9ahQo5RgRAvhv16Piv4SjggfDbjZplBA0UKOwgTU8ZOTwGxwhqgCvjM+to2I3uDBkxq/Hw+zaeymIKMscjIqD1D2VdnjEYYkaktX4Cso4BCYOo4jwCICPjoo9t+wNdztQmelA8CMBo/bAgABijSpKPZRt1zsXKrbYXT0CnIaIKKJC6zqEMQgvHRUlc1yBYeqmRxVvfq44KoyaVG7sCX4wth4mcuB7LeUqd1VpenGNDuKqo0J9IevRq/2Ck0vHAkXqk9dxjLlvHRWjo7C/r4DGbpSpoQquk/uu4UCL5ZjN71UUftGyZRBI5DhmXg2yuV4NwGgygSPfmw/dMSVOOl3HiKJOu58Hd5QpWTkqMltB7FHcpk3jlFhlco8khNGpAFsEQuX6xz4K5ZXKMBxVvZHXzlHRMnd26z3gkckXKRdsXHsG2cnkLpfrfleasqkceAZ/a6T29XP+1cvwAAAgAElEQVTSaveuHBUd6KhdVrQYAVi+azHH6aMxrWG8wDl5GLzI2WUUdUWP8/wgyA3O0n1q16LR27t+ck2DX+vwAhePIL9apd0d1P7aOSp4jqkkKjlbIlDns+PZccbjud++D1AE9JOfGSHML3eOCsin9wFc6gA+46goJ7+OegVz/a0dFV2m3cJ9oxy/nW/PvE3lqJ6rO4hwo9vcPriDO/oZ3y9cj6uDyjg7VBaML6NhTj5zkCwAEufboaH4JJ0yW3Q60PJVP9tRUSIF61T8MQdgrJ0hlUlChwf/1fm6DdMc++cX9wzHjeu5d9zMmlI/+4cnxeWpLwoy1cRx3DZgcO1hLMs7ynbqiJN82pBo56jAc+smlcnqqKgSX2tZBj6Ac6HL9QNHRRKor5ZH1k6lC7Ue+G2r6zzFiUYJqVmmTafTsA5rwoIaM00Yp2BP9V4Fd2jAbHqSA1QBgpEEXrLo1a5DiRoEbYUjyu6x8jJRvoT16lk2xoGxaE5sQKrPzadzo6Miqw7gPouG5tkJdRUBZSjdGnt/JMtGXDc7lJBFlA5yQDvmCvmHkihGVo/aDseB9wZ4fro8uMOin+iUu/Zo+96AWkbg49nnZYc9g/slpxPCwWntQDfkno0JvRgsjro4gWsHQP05y86gtA+yHAxodlzBAGZzrDwA/ARt04iIbPYAg4PX1LZxbCBKxrACAcDbLyjnHA5GlsDpGlVwcGTiIfMhskY8eDB6vnj/CwDoXJv7BzRuJkjtmRs2EEu08DI3vul8vsxw8J0YtiOAdeAsiOiP/h9BSGTiM2OpxsmtjLFA3rDske0vA3kra8qyTADqMjuCmE6WKGIWgrAI1xYBWCHDAvOxuaH8E8oX2f9YiomPUD3ct+OGAZOebj9XT4wdt9o86awkTalDMEsE+x89MpjVbbIZEf6ZROCgPN9POYWKHuA9lAZn6STYLaS59aaw/qbQb3S09bdnSo1HZzga/Y7Q5RVXmOYdD/f9GL8nTheT0V4oLjtH2dScFWtHRfaHuVwu5gQyhzEqjFjmiDm4qiSbyXN1ThiPcE/Yv1m+i5/HEWHrgiwqc6ih1DowNNDCvjc5bz/ekyLmgZLsKM0PhxKcUclrH6Wfzgv3jyv/LArw1Kcn84qj4t8io4Ln4DUnwVrvoJJi3+KA7g8tWpxxFuwoNwEZTQDNmgcdFTPAppFAMtpUlHmgluHlYJJ4+v38dc9vFvWT3yGJeEBAkIaM5smwnORGe2qpeniWOS+yQU97Fp7RlBs9FFcA5ZgKyNGGApW31y8ZbTCuCepFMlos4CoBmdbTHudtyiiVDqRG0gBzZSKMlhGYp4ITq+evWgJSTfFjML5aZ32UjXyyAdTw9NgQ5w+di66F7olyAPF8Hh0deTV5fLCa06DnhUNGhX28izk8o6Pz+QMlgrfCESH0dcNFHTUISPEfOtXUGCTfdIB2NbLByq+gtgXXx5x1KV35mddEJFIFUakgdObRtHV9xkYKZs87MdwaoiuOCmjzkY4a+zUUNVeK43XlZMCIE/hKgU1JCwkzgRwLkkJmqfEz7MoN9rA+GwjKh6w05TqzaCYYbSfaMbcDR0UzRH3sofT6a3XAR2s9otyQFB1XGAlGHqh3tMjPa44Kkwmspy31n+PNcIhdoIzOe21j5euFIR8IVCn+vjpr57Ow5FLj8EbSfqKDx9ikVwBivywZNxi2A8i630dKr/hLryF4IW855KcjR8XuxiOKd9A5nrBx+GE9WF6yAKKVEzBX4Bb05GDmu6je/S1rN1mu8yGVz34579Hk2eUjcH0Ltjic8ygHro/raC3Wdx/IzINsjgLbQ0YPzgZ9l46JfRsaeHF0rzxoy8eOLO5nt/rmWAqNyAPWYfUpxcbqHchDrJ1dutVwll5f1uUVZ3SefuMIuLRVij9ELi4znEMEtj6lZ0ay38FHAQajHDni7913K+eM6rlUls47KnoADWa205+CNoNMve6oWDSx33mZwhbBUUUdrOvjoON0OjX22O2JgE9nHoxofHsqHRW0D1ln3B0NkTFvkc0MjGM9f5YBZjkQBT953jB7okBFlrC1IXU6He7rRRlNFhtiBH++/72OChmA8qMtvztaoo69Y99WE//5OaLfCRYDMEbpqSjLFTqIPy/sWosW90wMA/ScxlsRuD2JUmwOfOWy2cuzAB+wcTv4GEGMk+0fGTwsWe3lklwwRu35ALzdMeX1ccmH2mMKEracd8R84KAgnziYS4eSZwGgybDdi14CEfktoCvGUuKNTZBRTgq0ZuUCRnVnnwhXdfFOlq0BThKBsm9wElifiYcvD97fwcv9ROChOUEc0wjnD0odEcsQfcBIQrKJPKFDn0C9l3YyZ0n0SiCt3TERthRBbZxN/dSqc7u+08/suczKSIdaOEBs3b3HSJTSllT2Ku+44DZzHng5IHNoReS+OgLHW+CAMv6OklQht4wHLTPHMmlsLCirhKbfGVAajlCTM8/PT1m2yIH3ANUNpCcHegkyCZaw4F06ntT5uttdb+Y0bS63zmt0oNHpBvE8SKkwcP3j2JQaCJm9V8IhR+yBc2hPc7ts7aiweXrzcu958YpspOBHiBbrIYPm4O4AYg+TcCxUikcFlyTmEWcQs4CIbTEY2eV7OFMp653O5qh7ec1erWzIbePUcnkfGRXvVBI/bvtbUoCH1g2OCmILYigvjXJVMRuQFiCVvzrMDdHzXDgtjPBRCF1zkigVGwgDF+SCyKMq1qCYhbGh8yjg1Q+n0PFoNHqz6WeFgocmrKLr+ugiZVBLZowD3kXV8nDM5tzRiGeOiiLtS7nhAalG4PheKHUgoSq/cZpj1QmIBZ3rMCHNmBrLqJ8qBJolsI5WKJ8PhTrnHI2QKMxdIbiEg2iwJ9xRkaAgjZ4KEeug7wKgzH2g7NR5Rs9N9WshiZXRYxUdS2VuRfNqcCvrRa5s9AjFVPTWeT1rD7jRovUdh5fv9tl6z/d9NfjyBoi4rqUeQUXdD/4hkmk9h4lS+EAjBrp+075HPAs/4nj2PXRWILWCJPGkHBS+25l4YxaGq8N5L5U0rE96NdRLnMZVD2sUmsx4H8jTnETH0BKul941Z44n+jYmYJabhmXeBJz9WRkVg5PX+bft8wVRToO+ZxwVUq/cl1QPt/ncYTp7OYQK2G8iK52Qg6OiI0PHq9McFcWb4x6/vrf76dPsg5GWjNqOTDmc750sfNooh844KsaxksLaiI9EWZ36/O7Pd1TQuMZ5QENst6C36D9HTPFrOipqxCsH2h+lyRYgDOm4fv5aTnZnQT+bd/jnfj0K/AixhZI4g9Oy7u/NX31H+/UdqGp/b3Tr5eyOHBWbzXSA+fqwj2ly/SyirpB7ehgH9g1kjINrHtV6W+mnAz/SwVa6xh810CWoUlrDEMGNqGLO6yxvIpui7yOVlavfd5M7cmIs1zRVGWgxZx0VqWdkD7qIwN5kKYKhOgMcOir8OYOjwhlqwx8bRwXoNNuLI3hJeu64eiuHSvkDACYZEnxznnNWmz7KnxAEA2gPPYE9IdRWg2NCslUi2ttB4ipGOrHD0e50G4yBeFEKykmLivZlK77XUSEkJ51TWjJyPSKHE7ALIWrgodPCIvU9wjj6n6VOhWa5bFDNGvFGM7Pht83TFxuG8ol6jl7i4vT11aOuvYQOmyZH+TCAxFGS1rNDLAodGR0FXFpE/qfL4w8rn2OAKLIpHr+jkS/2/LgnqlRZH3I0gfbMBzqpcC8zeFIPcSdC9VPAcghHZANsNKFGTbHP7mgANoCmyTZvZC3QqQynRj2qSjmhxNDv6A8RzhJ7tl1v2R9wyoXDxZ1A5ejknsm1k6HSOeHAcpROMtp5yZzILnIqxP43h4hl2tBRQZqw3DRkoDrJe3k9+14dZ06eiKy399vQyHMsIcX4T2RArSWz8zWziaIHhzsvNvqCn4XWZPz52d9vdDUaeGaOl9yyjKMHp2tVucDc6HiAkwO9Iw1jsvU12hkvWyYS+9GwhBKzLMwZYpH+epaQt0eeTPGq7MVgs2Bv4FAMgAqeDTme78j7A7OiXI31ejZnnJUQ8zkJT0VppLqdknq/FnBGWECwVU8Bb5r+gb4cKAvl/0bj8Crnx/0m/UyEII1e3hcIjin+2M62Bun2bsuKMQeJOVlJazgKw5HrDhnMkz8fjor13vr49JeiQGzFrA13vfTT0onAhlZyoKZekYAu64lHCmiL9pKDdWsAYaz6/tEgW5F2Hm8Af8t1KEMxzqk4JErCQbcRkDVuSbDFhMm9eVYLUNIDDQfyMMkENE34Y2D0xK7JsYdcTDC5MIuGSUgF7kZLTT0XZ4AvU4xNVFqBWP7ZkG6NJ8f/a+1CAWHYBIpNmOhg2OXaptCOrBMiXsUHOIjTUaEAfGOxDs674M/oEhHiyQSxJjWj8vaPiRG5tj3KTvEBKLG4UfnJD24q+43yUPmVbzpfD8BhnvTtDnmiEUMJkpblaek080HnyYaH0CDYPD12NkYUxoU6KvLJ/hyC9qs9wM0ooMD4TnWwilOt6KHPHd6Rmos8P34djdR6zc68A80rCiglZq5e7gcNbE0RJXWf+TJu5+YgFN9GRrDnoONdlK3Z3a5/fuSo2IgiH9Ik67DvrDZsRSgiTwD029FqZpxtRkVcCpnEtFpEw6zOgjhUTvL9OUcFJF+U9nuzhns8Z2di+TzCyE8wYdipJUrtWnFUnHGwLLyl10Dun+2owLaucmW+hZNX65xwAzBopefH4sScylTlO3T94/emM2xW+tBRMZz515hlBq9Za35zmguwTCPkGjh4bQxnv9/vuL3c2msfZ996fN2a/xYRc7pPxAnnkvSKl+C8pOFL1nes1jrvuP0lec6Xs+rIUQHHRPE++Ez1YvA+PtfhjDJgV0JhV/ppJ0N2ZYIIVo+0mf2s14m2u8L0XgcdJDr4XRx5fQiLx17jj64z7B06vK5skWNHxUE2x6B3c19M/MH+EWfOk9XMYzLznKCznnFU8LHIdIYBhMxj/2N4q0ig044KPmdxBm9lRehn2GA5prWeos7BxTs2jLh0FFPVN6CcpZ+iBJWunWtMEb1uADybBBsIxrI9FWWLASSgqnSlZy9oCZl2fg75XLVdPNO3hQJVLJvQIlf2xJ4rPUoeEH061Blh37KJLcuyZEUD6pqcc9CEmRbmRDAHgD/jioNztXbET1O/aWZW2eGu62Sz5QJwEfEN52qB7eVU8l4K3mz5u4PLtk9s3X///gMlX9KS1/ULZ4COJdbXHQBpL7C3ADjcS0lFbxN3okTpMezP4Kf8Bc282agZWwYly+AQCGdRNPw1jASAP0pCgdZsCIwGxl6eyBqLW2aHN98O4Nf6UAa+wcwKexbLmTHKPywLDjT5n3YXS6XZF0Y7A9q9vFqsuztWIlOHWQjkdWZysO+D2nHpSGtZKjh/c/85ToTG1zjDba9Dt4eDHf5Tu353Ntt3KAUHW8PnY86LjYLGDBX7nk4np5tl99x99r4T5hxyB5DRP0oR2bjpqEHmgDnEojn5kznd4LQwpwvkDdYC6ws85un5h2cTGG0tuwD7xNZ9bfc1c1D6uvieC5qkfZznRckF2FSUeQTUQqzF856sB4tlfsS5x54iaYsmj/M5RwEPyJawrBQ2SjeeeolyenRMYH3rrEDPE9HP0kmPPZa8FGcUHGmYGWT/W8qrH0+WdWR7yMpywcnpfBH9W1HKqwcqfjgqNgfzx8e/EgVqJ1IAIAXSlP3ny9uLeV6fLq/Pj5eXp++X/+t/fszBq6EyG2s4LqGmEHzlcchojtTG5JkzbUqHxPUEdtPAuZmcR46Kelg3oMZ310mQAjWAORfgd4hUyOZlHvESjZud5FWXPAVX6MI8ZZymV4ztceo8CF1YRbSGPce99RFhIzMclNEV2L0mbs4+lXdGAfenp6PCU1PpiUcmAQ5gEfzsz3EAVyaftWbk1YQbB6T0nSDwtVDQCIqRVj4ei3JwDQGkKbBsEaHIM09BtyJMgtCkyGwDInpGKRbnyrTHQsURxw94SO+d1wR7W8xjHG7DQVUTvRV+arBHY5SVk4LvXnJU7AmAmRE96BE5g871Ux0V2LA5ixx00GFjrHVnUc1mgQdfkUzx/khXJhiB58eopJk2H4Zh1Rh9T+z6sIiB30uf6RzxZHcgZEP7eFtOqjek14ltsY2RnWKNdY8yuddnvItq3FARjgru0JVRPUb4rWoN7+93mkyPPeGocOdXOSquZlT4I6MEVoD5YwTw6qzNz2akr1GsAbYDmLtj0DVQvJE3g7xuJJPzgVE9kLvzTwGz9e2RQyWdOsMZee3znZTbjEpkaL8TzdwPfgIIyZq3UdZgfwckc6/tu84uvSJYbvt6Q5A90L/L5bzttcek04arKmP3FOe679Z/fN8JXGy4ZX1H132r59rN6luKfc6dOscaNEypLQasyyw29RwcGABn+hzO0uqWlT1yVOCgwU7jUPT8wGdnVkbOyHGV4jwt0GHloD6e0Y1q9+HD6lwTTexQ1aJeUJkhZffMrwIYtB5Cgv50FLM2/6K8qjt3bmhLgDdyIhiAjiPBnnRU8IwfJx9ncJYDZaazPREA3tpRQdt1kMvgroEgYSMMwT550Ub3oD3lb1BbZ32CTeVgdBB7rp6/SdDTAMWoRe70pNrm5XG6jITdiRJArI3P97PxqoFiBA+R+c5MHYzBA0jyZ1gnz07f8VkBan6OkxlY3ifHas+sMocj326z+xY6Dt9BENfmlSWSIoPCo7m9dA/6QGIZcXBX5gj40kD2L9HnwQBku8ejwCV6eVrPxcbzTmuqN3d13d/lZX5eXyPK3npXorcGZbcNkb1GGh6AK52+HikdYLJda4DoeAbmvXZPgO8woai8IGPEz6rYaQ7MR2N2azJtY4XDAA16m9kprIv+KchqUFufgZNehi7ogqblcAi4Y130HjoJfEyvFcmPpugW9FO0yXr+0WfC5s+IdZbZYjbiiFGh2gVWlHR38D5KFmlpnbpGsl2N/lFSe6UrudMhZIY9k30p7L3eyPrlBY6JyNppfQMiq4N03Dkq7B5WoGAZKIxlf8BY1oiWf0KPk2fPrrD1pv5pUffeAyRsUDrtsL/R+4NVO/JMD57MPoQBpqMUmzVoR6N0+9fkWs1Lzw85z+IsT5kl/JaZplFynE3HmzQNfiMvGZfjTCyGT1klm5vYED+6pg9gv2L/mbOGTeThFdBzHyXpSH+jAXtUUJ5rWSYesc0hE8GNdj0wxod4b2TQxR5lg3pdP3c2hhObc/twVGwOtY+PfyUKUNkLyC6sq52j4r/++x/LwY+HAC7qjgqAkER1x0jiI829K8G17yMleqc8aUPNuKlAEr5vbuDXlJEgDza3NRN6c4FuwraUvrgjSQlAzBXHBP7i8Ihr/MBn34rPACdc+Eu5nvqdijyUClcozWstGRtLEohivTfrCIwsgMit9ROHdSo+ERGsKfbMeIjySn6gRdaNGsdeazivDaVBj1kV8qP5kVpG8Q4V/PRYs26hAIf5/khzJj2dN0wxkrTJMqZ77dw8wALM9JYPOYxuvK0Vf/BDKpZkIeePuVGqxkLiPQCL6lDu4FGVPQmVpQH8uH/6GYH6vGA0pHbz0yfGvpK1VfMxX8UILjEgU5HQYQ6Kf1AvXihp5WJK6Qw5AxqcjEBxcTeRQj54O5YPXVYoneoZYySpGt6633NNfGEpKKhJQ+EBX3P1S2ZPPSqcdlL33pHz1Molaj0+G5Qpr9PqEU00LNmUrhSvmd8bNXpaODWu+LeXCLAPK/rl9Olo+9QjtpBiy4jhTItd6utrXt5Cr0svzFHkZHB5yBs0CS/DuJCGmuXIf7eCh3r96XvjbMByzPImHSUiExKsyTWUOehZMfBSlwqQWWcB05Tj8pAj5wWmA57evYOPats+I5pGiRpnb+NfPAEr3fmJRk8bo9BjMkJyXt2YqfGvZco1Guz20MoBNe4I3rtzHOK8PtLXTu/gmy/cO0/2Dp3tPQdTIHBxjRarCVzrkzGqVV2OdnCakZ/79TxX0ujaPjqi64pnVvvrlsXsDondQqwB+KVIjpcTpKGOdI1++zHvdsV4xxldaMklQyBL2TjY2/r3KEFXz5v5Bo9Y03YFzviabom7pscENF9DdLZOqLLH9BJkVKysl4pCnueomiZpVVmN1J/sudQdPBtcda4EuDZ8IDqanhjeqNRtxbfL/YMB0NZjwnSpzTps2UxOlkGP2Z8h5UypE4pANHsBVFAXTQKCjBihBJFllYTSG3fnzn63RDPmOJf5jlU5HpypR+ECBab7CtN+E/r4yWSgYdjemhGRcmwIEiSH2LUGzjLq+JqM4x5aOVtau4gMrsSb6DQyB4CBxnd3cFT058ARpWVbUkbHHlWbEIB2ZPBGzLRKCdeNo7Qq+B6N61luSO1cew/Bbwfu2Zsi7H0PaIoSy+4covNL9SFxnlY5MfAeAfmnl+h/4OW6QHfbN3Q2GMZCfnPng7yf2ArBWs7VgVjFXHyuAHTtczgxnv0zzj0bgEcWgDkfzKnw+++/O52+fvvm4LO/0zMDnjMA1d8b9NRyYU5DNg6PwTGzScdOcJq8ls6A2C/gMbyDc9DnIvjHskxePfsF2JTR9S6aeFeDbdsb5nhgBD8DactBBhCdTbRHTI9/c8zOIzF/n6Jk5bkDhdlICd4jyt/fe3efMpGZUFr5g9lPVobK5mP3GQ2YAeN4meA3fm/YgN5APf4Dr31Cg3fyD7M8bPReYh0yihl89mvZkBFqHQKO/G7XohQZswVzoTKjNbMZImA43x+OZGZLLU9zlvPSfrByYbf5kD1nP3Swsh8t9T7V/8Z1/XBUrFbg47NfjALcgWcdFU/L8Y/p57wIKiM85gZ8Qb+rxrCl+BQguNd110b7zmbm5qRg5buof1WUUoARWgYekjfnakLFBKoJTG865OmIiE4BNipeWv9T1FcB1DPSxYEii4oIRcBTNhfGRqN2CVVkDaxZqTfVKtBzViZDbYwIgknh34BPDiraoUBHRWRL4CCOsiQSCd4P5g4k9fIfMZ8BRAN18bM0pBbNj1OQa0ZPPEiFvPMGUyciyub+Ek2gcv3JH2pMFTVfW+mnPfpRvD7Xlc75ZTOw/pyVo6Kv/oGjYuWAWDV1zVfWfqAChXeNn2/4L0pP+Hzf4agYWD4WPgx3HYco5LXeETWlD1GHpU8jgLawf1+nJVuBk3rROaOdQ6gU2M77ff/K88MIhn5Kh1SNCQEzLGlE4076IsQcsXakB9JFoY9VPViuEW9hfVNEorEZWpQe4bT93Y3AC0bYmZxIa1bvUJb62W+dNaP5voXym45fq78ZhtOGO4ePSdfNy9/jqAjZjzPPrOZ6duMclvMaXn3a2SCg/GquR+BjW73mTIcTbAapofAX4DJk3w2OtRIla7oeORFoZDjvi9NhPMc3TPFTHBWcXZ/lPJexXJSPXYzxcYy75rZbAMjpmhtvUbpsR4W9bB4d4dso1u2j/yw3xex84hAPAbRtwMU12rE3AGTm8RrFCZno3/7ZCT6kz7efLT1A5ahJs0v4a5M49700w515Vns+YKxnZcvy5VnGsPj6nKw+N5W1LLz13h1doTRwjWBjSDmPm16jaxv6TWukffZhqT36DRwTwsbPyV++6T2Oitt5YaStjHHy2hOFnu+pM2rRHHuRUcEIegBsADQNuEM99wCrBn31IFUFJKNDA5RP4I5Zo/apA1RLZ0t7xLTYO7l86KhYsMx+fSpDI28L+rMuPhs+81zbqWi73YLmswABS9eUQI/hRtXydSp+CjLQTcqeHJ1dLeBJROX2HjknclgHjjfI8dq3eAX+Hn08YxqCAYlWT95qyZdeUzOmTNEyfqpbvMR5xFrz9jfoU+VGdTy+DtHDgTX5PZrbwd0uh+mocHA3QV3yalXIcL62dTXswrOxIpNGFo5jYsAOsQDbez+eHqPkaT3b9HjLarESNua08D0a5YRA18oCYmko+36nG1oDbpsjKltYBosB3ujbEm/1dbD9atkE37599dI9zMqwayw6/vvv6JNhPKzjMXuJ1HOMyJpJR8mqa2XDVtLdbJmYIuR48hhs6a9fvnqWj41h7Hlh7/7iPMWm1VV6iVlW1Knp4OF6EKy3OaQDJ5w7eTaI8xay8yX3NcfK52YfBisp9RnOHXcgSqCtOwOiqobdj3JdwMGyDJg5YaKknc8rnpElu4Ll6WRk9GbalLE45hBk9pHNx5xefk+UFFMZOTqPuI/cgcHskmhmr+c/zl7ZJ+yTFU4Sfe5q7fmZPVOdUcysanI/3gN+fEEjde9z8uDZKk5PcwrF51x3YqL6/A9HxdFqfHz3i1AgdvLJHhX/9d+vHRVr0Fz6ALCsTwD0/XAs9QdwyPrH79FoTQeur5tq/RAbD1MB3RQgH4ZA4WHPsrQtEw6eZgvUkOGVdZf2a/AJ4Ro22cFUCPxi1mnwREOoTE8TQMoPxlBSrLzU/qeMbB7Ia8pqKsDwPAVJONYwUinwbD1Yw5FNwKiU1uEFAT8adFjPmIE8HweDkFIVnxWjedR7PmgiSSqmQ/8U6AB4k4IQn0emivUr0CxewYM7cVfhYwHYxuf730PJqxZp3Xgc/GoNwfEzvwOf5snlVyGCJioCnXFU5Bz7evizoplbvT5P4yX7cU+gsVn95J4f5of1no1qt5n6A4YPAjyV58EpqsxTwAqmGHtOrpqNLO5LpXeBARvbv9c9aJSB8sX1g5hZG+tN0bnmqEjn6IBu6B5hnWcBmTUSBU66mq/JFwf6I60XETBWD/ZeeEz25sZbGnEoS/7APuqC26XokThbPMkpGIYWnRNQ6syBvI40nuutzzzEV+H5q0HJZ40ZwjkjjgoozhqB3kv+Oe+vnNoHYODnNwFmFuPTY8z5bBvNCYeVO3k2slBWuq3ASt70bXdlMXM7cD+KnJAzBucGS8WsywGNrLFy9KxA5px3LUcAACAASURBVElOLHimlw2Y55QGEbNHYVnuQe3ba6ss99B7P2QtZKXHDmTavePGbfreof7V7zueN/Q67qUsM3ByVLjvPKVWBi4z7wa1t43gZpB4O+k9NRwkXJSZOeO42ZHrAP87ReHzlMXjbqbTxgVUsrX0Rswl7IBTo28nTIzv7I2rdSrdBEcW6+BrY6v+/CU9/EjeUXbNHzu6JkmW0xrfoX+P3/G9s750q6OCdgnLq9q555mjBgxdALol/cA055QS2oAxV5TkuXOQyJ5t5Wp2pVu2+wNcsfx656jY7eAt7zuph7vEUWER91quEQ66zZh2DtNw4jEzxmXGWy+jq5NEzN+su9Ue8wsyy8b11A0R+z0lAypQcbixhHCj/q5HD3i86MFfvW311oBFQ+/naF7sQKP1gYggziYZskly2HPS6Jy6KQD30DtDL3RavxlP19NQrQGOBXu//XimA3GIHK8rrJD3USGB2RWUow6COhiOuTCa2/pHlJUTkEj0WOB5SIDUI+5thFEqiGWW3PGS0fgWCY/yQ7BZXN2H6RDlDdkLwIOVGHDI4C4vVYZ+HuiVgWh+dyREpgVLPZkTx4B3b06eoG9E/b9dLt8fv0dmCQKtHOS2nha+dtGfwZyebnugBFnu+WHPHOkdqGQScsizscm30fQ8ovOb/sZeEbEmcBagX4L2MvBmzl4iDCXJ7Rnek8IzeoDRPJujJEoYZQntcCbQrrcxWikrrlk5INEoHrwDbMy+Q5+Ll8vrW5SRih0LZyjmyr4WsOPgREAwLLJhEByMai50rjgPstRXzJ3Nzov1weMm5+nccJkcjhY2F6esB/erAxpnqOr51oDbfrxHijhVXDKFMGqyJ/m1yoZxHivR5edR9BlRjNB7DrGMPm/0/hPM3MP+tvHD0YPMJ+JwkJwYpOJeH46KzQHy8fGvRIEQmycdFf/3/4IDar3B5k9p5GRkdToquKkJJOLegLCuE6iBk5t0UW3azL4F0lyuXpLNCErxUGA+LuQB4opnCPP2DBm1VvMsuBZRPO5ssL5Qd0hF9MwKps1RcQiJSTCfzXActAkHwi6dOGXYlCGyXDX5sKt8I1XTHBIFytdL0hJVUYGAhFCko6LGFgCUkB4MQH6Iw1onw3WIf5Wuug4l3LGcBPlHwzqdLRIBOxpY9Y4ONvNASKZtPQIwmtHAb9Q1BsCpEY8A54c6pu6IjCKADRHXy+/4VLIXjO5xUPWMBgUFF8WIF3PgPHIZGo9vtqkYeM2EpsK2cFTU7q9nunK9tEI6zfooes8T0kYVDb1+rTSuaFwz2eFPxwZTjGTgbx1L8y844aMZNKDPZDXYxQC/4eARg1qcDv4ICe0C/0cJpwHgTgXLDAdXhtEMzY2ZMLx3wNSKC3xc6qzN0a84iau/o+D8BhhqZrhUUzdTzrRB3Gpc8xuUl/odNAbn58hTBkcFlmkGVdKIMqCaDs64jo6Ks/T9JI4Krps9v5d7Y9nFI0c+lHimIK+ctjX3mrM6t3S3Nl6OP/ZG2ZCroOc566iLA/momeBKrmP7SM3mhdxqvBB7Y8cfGZDQniOR1bE/r2UnvL3DUaHn1Ebinv74FkfF1nF4ZGmfHsmff+FuGgBVCrQUUbwZdChrw7f77JkQXgtwD/qd6sZjidRBRt2K+N96fQx1BCgJFixl/w7MfM+714fLlnl2J8itQLHqZuPLqH/TkXWNP37etPeOB4xRgHYqsjfsVV56wy0Jak40Wh2DcVGW1Wg3xcrxYM/v2Eh2PlMDQRqCVwgqjdfj3HUQKOKjaIuZHfX6Fo6KzGC9wVGRY4VNY/bdl4evaET8uWrm3yLxMPr1StzqqNi/NwBuvWDITtezp/h+fuI2+8OYP6YBQDPUnw2TIUZso5U3ex78gqyA9a4HnepZlGFXHRXc0I0um7XgNdTposAC7fbVMtr8GNEPB0LX4fM0CQCaNn8GLgY4iVJJ0XzZHR1sTu0GQo3eY8Be3ZZiTwRElzNjwsBxXN6CPKL2fz4tvLSGW1hFCbMPrGyV87mvreigeFiUH0KTZ0wTdCTQ/+YOhuo5YV9bFoRlLxBj8T1rADgdFeFk4Xgd2JYG0smzFhjqjaFfPaIf47USU+BJt29sv/p3d9HgGfu3moKH49dsixg7AlVR/omNk22f2zu+fvni36VzJ3X9WI5Nf7YSd+IMpEgMh5LRgA3E3bFlZaientw+s7HYD/p4GK21rDSi652PvPkyrrfrUFYJFU+QWVIZPv5sd7pY2a3I9GA/jQjSJW8QDE+9KbJfyE9Yn2p2bmtbpZiq5BqDzFx3N0dpNFNnJRIrp0cHCfuTMHtjl+drZHS6fPoEx9Ll0+XhywNwOHOWxH5Ph0tibIMsClHGzA+WEYMNBVt5FEVhqjdbpDC8tWRWRwVtM+6BlWgEi8EhZLY7+5bA2WNjg43spesXr/xwVNxyMn9c+ydRIFj3pKPi//lfd46KBknifB7OS4KmMODGLwNvk8PyiCAUSqgitUhhxbHblPcSpvsnp5E49k2I4ebxT4dLRIKPyhIdFWPpCBP6rsyGx9gOHgfY5ACjF9pBdk8bRqriGL15BEHZMzjWNNKWCp0qeYPCRyGuak8oiz7fOIRL4YcxAOEMwUnlBMpDKUMEWVk6o9F1VBSHcWMp4g7XfXv6aluLA8VXucBrGcacVJFNp4cATJxHrsdYCkfc6jwYZlWaTQJlLmNs0ADe+R05bfxSzw/FJIHwuQSSgt3LrolD5HXuaAXChReuGbR+f9BUr53WmgsxeABGo4WQcq2bfTJSlmn2SteD/b78Kt6ECcQV8p4JgMclW3rkF6hnCfbuUVe11OG5E7AWNOQwpEdFiDc4BWp8zeHhthqiozgXALhrmlDpQh3dcmZ5dE04Hc8cVLc4Kt5dSMbGdwdjiIpsZoQs0CFQYDXxNTGg/127fvx+4aBhRoVfGjRVZ8WNDUzpqNChuaMiSkwAD8C4KF+P9ioNu9OOCn9x340KLihF9u8VN/Mo3xeOCt8voyE9OCPIl5PjQhl2LANXN7nbb/zpbNTXGiBD1VzO8PuIcVztk1sdFTqXESw+sw/n+eDcGc/Im551TfDf9LA/8eKNDPSAAV/4cnQNR+Aw6Dwp83Ncv33BdIoWn/11HRW7ER3y1uC4OZYT++wFfccZp+zRmDZH8JaZbmXZqw7HpTNpf6ZuvpGPj3iFl50rA1a69jXHxszGgiu3L4/0hZXmM+o3XQQfHHiL0k/YG+MKhvLjX81yeb5+dlQY2Gf16pEJjv/9v+y96ZYlSc4cdnOprOoh9RTfJ1LUIfk2+i8efqJIvYmel1J35a5jMBgA93DEjciqnq6hMuf0VOa9sfgCh8PNsMw266H1EoOTKY3h5QrQ7zRB5gPF3q6l9mcRFZTx6R0+llyfmTom569pU9dWCVSJZnfVulwSHVGRgBs9wmGb4jMDDc8SFW0MhgZ/HP0uomIzQwLhp2U36xIjsh4ezHNfpIVSJg/7fSz7ODh7tBTlVJHRACLxt9JIWTFowTr+LyKGDHOA939JqWlRP+b9TlHgd3wxo/LlOpdnOQHk5mh5e2cAPX4MTPU2Rz/eVVsB/9JhES94eny8PHx9MGv4GRET72+XL4gAuLm15xFEf7E22Vg5DmIR8yIuSh7/FKbci0kawtmNBYRVr0DXPj8zLZTqOhhm4YAzrsHvGFMeYR0AAskEzMYIIhIABibDsx7ZNu4JpFstCI8OCafGmbRYrYACkgd85VHPlurJIzU0jkp7pfobrDEBYkFzWIgG1OXwujkvGFuvaQAZwFggbZBFS2BtITXX46PNFQs/e6Hmm1vrs+lOpf72uedRc4y6Eg5FzCuxQ3Oz8zOp6WDUKHFgPcisV9aDVR/RXkR/iAAeIiqgE3w+ahv4fu4VRrhYuiqfW6S2iqwoKfuGuzkBuLEDeCj0qIS3i41jqYvCtTPag0aET/Vcd20bj6jAfbMTGddl0cHvTPcEObbaK4i6KMYqWoJImtDlTvgN+/G//9/+77P20VJ5f374OQJ/3ghoR3P2kMgyN6m3l8u7Cf/z5e3l8fL6/P1ylKiItSTws3g3jkRFGpziG/YOMRVoglKwAKeWqOCoaWM2RWoLtea+riOrzcjxqZqvtOTYlIfxqJQduJmA4sTTHSZzxaliW1FEykMb1V6FdM5eBSQt5LmwAwOdICpGyKmYpLNFWQzCWixJRaL0rw/6PlHh4OsrZ7CFEAcANoqzK4LA57akzRoANGtv55WfG7lIFQFNr1PRb2524+Gq7hUFtwtgU1JNz4Dy48C9FzYhmOFF0Ggd+tXDhicZL0/y79ODIYkKO6ianI/vvkpU6PEV9K4b4/x5o5SilWnxJi05PSPAcyf8htVYSKbxmbKkF8fImkanjny9dNznF73QWq5GRzE+mtNrtxoteMYPapFmx0JkpZ/UhDL3K6JCxbSd45KetAOLbs2Bojj5S/T+JA7Xk0eiwlMieL5QfHavehV+2zXQNIiKGLb1oMW6ym3g+FZnnfJi2pHvdAq7rktvSYJLlravpU26anf9bPyeumCSBNSooPq/XBQNUQ8tt1vJEXmwGowb1bzwtqmJ8owyh4DSrX0jtB5Ma+2c5ZuHFHu15yqOWffu61Pq68xfFYQJBXc4UFfjWy3T/rshJqY5m/Vv6sxRL1eiIuW7n+uBqKjv9HRrqxE8S1TIHpjXG8nGRhHtrKBVRMU13GbzuP9RTjXt8M1ExTVJzr2hEg4sTNtNBp85EmEOkP2JERVnJYbgQ0YpkrzuU8DsKe9PomIcnbo3uyWg3fX4Hhj7sSlN++v/P0TFZDfFxkDbd/zxSEZFGyN3ukeCQ6QDjJzOfN1EVALC1pQOAa6XkR7EouDl9d+kX+yeP0Llk9w0IQH7ajnPtjpv7REVdd+xwtRODHR599uIiojord76vVdPH1HhdRENfFZBYNYEaIkKG5AcFa239+KAU0dWNReHcZT9vLenpkFiv8luzNQ/vEBjBHvd0j+5Vz6+U6TDsKd7yh09ns6KcF58tZoQ+Jt15OidLix9Pqvi/tf3V8vaQGCW6YVwHsSzEBUR6YYKiaHUPBi30ZFPhaLprW1e+FajoqR+UsS3zwHe8fiIwuF39t8f3/9g9AE8+t9Zp1NR4gbOIkWRRRIg1TbAahbeJkjukd5eR89woMmbnfzY++Xl+dVSn7JgedZIQFYMFZ1WUXOOPYkI4S8gwnCt6j5Y9IaiDOChLr8yA8JRtwFp30o6bdn5R0gKE5IsBF3PABhnttfTTsFxzFO24jbVq8B4kkjB0UjnWP5bQW+m63r3OqskvSyNlqe9UnowA+29noN57CtlEkhCr3Vo4yasReSRh63RIZXSr+fgL4yp5gPvwN+McPDUTl6fwxywvEaFzb2lHaMMBFHnxcQpN8VpudRjVDSSLDnTBWjYLaNMQju6wRbE4WQc8xzCNZRZVWQP6Sw1WVk3GT2SJCE+W2tsOf6qBouNGyLHFnuInQPeue7SnsiC8jWKosrTcE77JCp2tPvnV7/ICJwkKv45Q2SHDswhbQLhTGn7lYGoLHxFypodsLYK3NICsIdVIAYbanr/1sVfrhWBYMymGNEeIKrKV4a/2GEabvRsjqI0xYuVCphK1e51GJ6eAAIY+J0iJQiOu7dDDBcPzFIqLAKngwiN8SiWq0LlspQOnUgFFHkBroVS3hqgvumVME+NhfVvqL1A4N0MHXltiDjyPvL6rL/AA0NpfIwrP6Pf00hUGMY9GKUhcAQNp7EYSYa8lsYYjR79aM63nvva8gqIMQCH3t7wxBgxz4HAGEAuTX7KuqY02hRfzZPMtphxMH9l69NpPpEj1UN5ArWLW00D1vaek7EJJn6TqqKuE57wIjJnVIiZumYciYVgl8JoM/pf/LbHQ8vSAywNuzWo4uBSVUBHtHiQBdWApSx30QRad5kyqLTNge/CA7me8JGqQySdWbPbjYp76kF6FXEtUvrMgy1cfHiL+3UNynzQvjepPaRp8gBedM+RMVzpMwtpH3Uko0foIVZW5hqLlfzNC6y0ZywuujIsi64peMXQpUpUbAprp36aQc0RxKyN0ubK+eZ6w3rxmhMgVct4qdWU6a0xHdGJpki1JHkX26S5qlNdajtdCWev0W+DIqiqzn+nuKl/i9VRhH5t5o/+TDNxsprqUbR0ZNHT9zfSOODMe2fnYdqwAjpIzUuhRjV1Hrb98snW6Zoc2v1+7SyJXV5jRWB+hFA5ohLma/bJ0yKvunE5BP7hQBRX4dxvWeo3yKEn1O6GutgsKcudVPs6nL8upOhKX4w6xTVi84q9KIJ6COYS3Wvneox2iYquTe1r1l9c0wmrli3vGezJeldGPA4s1M5wtCBuGcO0M2dbtrx7Z8nWvOYG7niNsuurfBqRYo7V/XNPx1QtE9pT47f8cvs0WkJpX0GsZesvFY6ReQSM6F3PqFMW210Radkxkd7Mgc6I9ZvBVqm2+7rnLDLsDiilgdZdLwwL4NLOE35uW5GS03YXe22SCFM9h3KeiM1ae40bbL7L+0lJtd8UwY2+6fe10KpvKtQMWSKQXFKJboaF9oc1L6Ifc8ead/KVLmDX1qtF+yPuA2AJcBltsvQvsmlmZ4HoXtGuVreAP1l/6lpNjB2dn+wA++1OQ+FEJHOGA+Myw7MNwEcUvmWtCNk85V0CWmO/ogzb+dTwUuIHJCnk2EHvfqwfc8kMx0gg1zx/YPxsELwGAudLtl8WmcYzQSJQzsdUQiqkfHuHefBneqFjnvdpk1ZDlNEJDna75z/WnwH/d3f2HeYTxATIKO0ztzdMPYS+Pr+9XL5YOqespYA+sf7GOE/ER0A83AfRYZEAXmwa42gZLRyzQOQAUlrRnFb6ZPYdxb3xXnOOce98YT+ma50IUDoikQJokcg9ES3qlwirSM1jdS+YcQPRJErnhPbef+G7KbeMUpEzDz4TUSFsCilxiYtwraPNnKf3y8vL0wVjqkgJPFUEBa2MxHGsv47fGFYlosaiNjxNlORIZJxFJCCFMOffIqAuN5e7L/dWZwIkCCPAva6Iny+V0ol1cW5Nfq3otREVqJvo0TQWNaBeac55RjUs0E/61DmmtFyWPEqo1ACxdWjryZV56S91DYkn/E6nYmJZJFUY8YHPEJHCs1M5XxWFXx2EfKvylG8mDWWdkAhRTQ0rRO7RL5WY4uSy78a5eFYBSyXv5Dj3tSz+TjLK9bi3zbr9SVTsKPjPr36REZC0O+NvUt9HVPzv/4wNxM1KFeEs0QBcOVR3dl0lKmqPI1/h1pQOz0YBv65wtNjr5kdwnBujfsdr5PEf4IwX9qUd1Rxy4BQAj4NIoUE2F2xvV7IrruUO4n2nQqDBN8aBVuCh/k4C486VIudCniI0dB0siuHihmm5VX2TJHtdjfTxnoL/uIbTTIYltPDS5FhpzOo4jNEtbtzbIWESbT9UrAT+5sLwV7ZERV15ZQIcafDwSv/e5zRzs29lqT8/+uZTcmcqd24YBDEsCV54w6IrNuZuqBDT8wPXgBAsjoubydhSIdNyGYZPY1NZcl1gRmtsSP5pPeDMREV0rxy+ROwNpuY4g+tyxXnNEiSpIzcN6xmFGDIwjDkjpmKOIpd/Ft9L6SnGi+TJvcZyHLd92eiB0skOkFsXdh5Wz9D1elSTTIV0mGWR0T0x/zK0yvhu11C+ptbQqS8/BipKr7imLouyHAkjE04Fu0ejbJzxsd+LNVM+4rprJGZK2xfz6Yb0cGhekYTDgLhOch3lMXyFGPeIKApdenLWtkIOZxWCdHV+ZJ4Jinh90783FZuMfs5jdS2XlKflw4ty+x+MZerAUuPB36U9bSsnq8Zmu0i41b/Xczc/ZSEFmxsHXRBrudbscHn17wZv2GnwdeDnbP78n7dmsjubJNf/oi3dAtg0vApf7qU/u3c2D02bjumV6y0KAGh6zzXgfPX+Xl/3VsP1Fg7KI0m+sGW55NbtDWh2ek2d0Hly1VbZaeOtKW6671r6oGZdLgrNnxuLsc/j2JfUhoceqroFhy6mZm4Wc7uHFN14/C3nruyIm1YXtH1Im79bHxyDYxptfv+1tXWu172OqPu0/S4wZSnytOlUPNVAJAdsAcCugfA8y9Sx0F43rZzdbqn2Xh3XvXHaHVNfwkrLIzBUm3PI6OLMMGsbXuLOSh+MfDIw/J3FePGDcU2QdW1bJDnGs6/ORd0ZoY6HHMR4VG4KmDv5wfM0vd7xI9BZ4HIdjzFFVup0eILjL0YjIH2Ukx3VY7lsAT1eQE9pYA/0dM+I1GpHoFc8llzfV8Z3rSPuuDRyUcRTffxI2tGaFsEkEHgl1JKZWH+yCZ3wU1+EL6CfWG9cf6xhZwWqbzmWBuB7hDOfqfU42mF4jQpTYx2DNHh+eWb0dsFS6sghLRRS3YSDqDc6cA8vsi3/N0RifP321YBl8y4351ISFADaLUWbozuIugDgD4CdNRSQ1gkRIAlML8evgMZsq0cPeP4lYEpaS0hzNes51lnhujKiwiNsVE9D48soE9aXQF9UI4MjrDogBNcVmRH6yWUCwDrqNIjkwO9YJySKsG5zs8QtaBvAf6WxwnhiDEEcsJ4FoyFIxjjBYWSaky7eF6xX9AtkFdotAsSI5nI4MizP0kLdXl5snUoY3UnXQfnEAjmaXA6+XkL2icXgXeyDargogo73GukmxNIJP4ve8HYhXRaiWSSHNv4qSo5oJBAq/owY72Lj0ZGX/eB5XU8aP4/2O9FwZ2Qsa5+QLFlJ34Xpxt5emaZMl0T2BRaJR/0R6krxKbzSSM1PomI9sJ+f/kojkEgFWfVrRAWUHFc1jT33aF0e60vKi7bLs+FjO8kEauR70oOUDzRl6sRENdJlxBrTqLQrbqgHgTC36eYmcgBKkSv0b4+osPfqEODahIYdNwwrfOQFoCJ8qxQ7IsBFper7SSg1/EKWWOBgabRF4dMj1xSgFUoatdnqbBJGuqY7HpkQHq9Zg09pTKlNxWia0p7M5MNmyC/YJMaCkcRc9cxMn+CqPvKuz+GoLfCwkb1st3kzqFDXNIchYLp/AoNHT2RtRC7PR4iKA8BdvNp/OXzY1OKw3WgF5bGdw4HNptwLOJexaM3rncP/lqTQFmlvXQ7tUkXsAHuDUeX9nYkK6ah8to5OTlREl6ljBtxaB8jc/WOjzyVTjO8WDZmPa/PArQZyfvkWrNoetusIzmtzfMdZomJ7RuZ4xU9uI2VoFsTXzllNRulIJBDgmj9z7d/CyTsjmm2mAPHvaNd0Z8ypQERcqJoffr9ZySQsbFzLI2yOFFER6jrr4Zih2Kyj7lwroiLnf35AT1ToHnpHcb+oY6soGR5Oy1CVIqOj0a2Bmyd2bFMlKrruDtMgfXdA79X21BUwE9h673aP5Dfzc/baudRVBz7siIr2FLIHLu6irF1jpnV7oM2/+iUjKHS8tf8YREXZKzdhklA7XHcpCmubbaOop2HaEyVTYSXHstbK2fHr1il15/F5M+DvpOyfJSrKrn64YR8B9Fdj8hGiouqvABbnaMODPZnbJFDp4O3XL2sJVu3FKQy9WBSiwqMKzTPa0NlMTzbaf2NaFTX0I0RFgq9yTtqPMqryupxf95AnkFVtjYn7nc4gdbBpvuuUpD2tdyfqxlZtCMDbz7CsDUFwf/6J9DC3twZ64sfAux3jRmIw121bqTk8TxE39rs7KBqw7DjE1nYvclRk7qYAq/Ycz42f8hC/Tbp17LX6DKC2pj0W+G4Oju7VrkwKe6QHn17bXN836/m0ToZ5LNGteJdF9Xhh4/7dY3+pSy6XGwPsiWFoHvGM79+/G/D55QsJAJAT93dfzPZFHQLZk7Ee4/GjRcU1QZLHIhZAjJVIhm2rLkaMyJvdij97HQ0NHe3pYtNbhA4jXfA50yKxzgl+bm/vY4HhO6uX4KmecI1qP3BM1iumA6lVrNr0MdJVwekV4LMXI8fnipqwsVC0zOXCaAfz1H/2eiYvLAjtRbTxTvRfxbDRPou6eCMwjRRQeL/SB1nfb29t7uhVz4gRfM6i0EhlRP1J0idlUTUrhjoqiDbw6AUjVBxDAYFSUxdp70C/QYpYmrHAyG6sxoMRF5gfH2OSUXd2bMr0aYWosCPYeo/gudadRZ0kiVoajmkxjV0WaBfpJb1nPXd7B22FXKg+iKW7kiO0OyLjvnpv6hGPRgmioqbZFWmhc5bWBiKthMEkxiobbCWCaqtqUVBPZ2YEkEvfvn4zMgN6yOo4om6FIIZPomKxo31+9IuNQCJMx4mKEcwcgeUZ6Om7G6FZ5RLqR3lF8wsrlpzwpn/Wu0nR0CtFLqcmGFHRNMuKFRWvbIaweQj/6p4ZwfO/TRk78aFNzkCh2ERrQcttzQxyHwKTnKiI9C0eZqvQTn9mHijK4TYMPG98nR4bhOJ5WhA2tXM0/nIWuNlMRTlL8Vbdd42ouL1BGJ9CkZNxHkC40gjChC4XC/BsOa0bYzmPoQwXdONeBzs9xO8bCIkYRh/IUmiSo6nP60DvQ16HALGpDxqf1vhcD0Qh1LaALF6hGY7n7xhoxxDWURa3gPeeOuxHRuuLY54/ubIxEzpU1StmokLfbVODjGfC6WAQslFefpaoKLpgHIVturKxl9t1V+VgDWCPY/lRosLGOx6VY7dRqHGN9AR70KTltO7bIWNA+X1UMiORNoTYF/akZ/5u0PmxfPFL9cDMceJ6SAOSL6X8jGOsg1EW5RyueWPhOJPNWl/CAYk9LHq55Wwqyc66pl83MqrT02hOP2bHhfRkmshM7WW1f9eAnqMkhfqau8xxL+A6Tpqb8YCSK2gFctaDRux9Z4Tr4LV/KVFhAn1otznYm3/MyzqAPeTvJAjej8IY+aa9qrM9FVk6ovZFx7rWG9+3BiL7LvTQ7+qe2KLKoZz6sqZbnXav09EX1MHHfzLl6fF71le2mPlyrPff9hGijcJGSAAAIABJREFUQvq0gh1niYqaWqSmgRn3qWz7ClTZ7JVDTcFeZs6Ov413Jx/NRrg9rVGPRfS7y468euGczGweBOJStkaiIsdB/av9pDz26ygrGoWFsEMi1NoOK1ttJpdSF+QIX1NLSpdFJ7sSCdrcuEtUKDrF9gyBdfQwX/5439PrnnUQQAo0N8TYiqiwiIQdxpLYQNqTPO/ah4OTUQVZtb50Ff4lMOtANc6/fo4e1l0F/FshTwc7DBPAXvwo7U+QTu70Yfn9vQbAar2l9/ikT+cxse66XAtv8FtMFivYv8EGrunBIhWlDoDmdSQtSdDgM5JSSEnhFnyJ6GCEAdNRxdM9owaaX2snhB4UUOzNDXAbUQ9WfBuFq7+wdoSnE475Kya7kSdOmEHOrGD024UFmVHvE46K3ijVrQiHqYOG+TgmbPCswyVvBurbHJH8t2gGS2vkacS9gDfAe4yFCIcgIAkMBXmkOjs15ZTJICIkPBoKxIWiMhSJgWsU+WKOmnbk1KGo7MUFz8K4W7SUUk/5ZYGZWRFoFKi+M+99i7JxQtHebyTFW9QGYSkPPs/qbxhexuLsFkFgxdk9zVn8y+U+j2/VZUpVR4LKyWs71tDBQcSmkQ8Y+6jBc2MkT6Sk8nXEuhyoi8P24xoRPNpvVY+otst+rwJvkpHCSf2g87SclFkAvhKfjF6pyNe4hqV3cB3k2Yg8j2qCqCCdGdN8MTLO5rtM8WdExVkr5vP6v2AEfCUp7NIW117qp0dXap4XVOx7hE1OB46d80dHVFQQbUwZkUwp92M+nDooVRV+t/BEN5JCybtRsmd2b4kKKt5rB6lqrMqOCDDI88ch/I/MM/OG1gOzfheZQfJXqZx0KExQCe9QSJ6BYFKKHXAuyYpIGLf5itIf82HrhgTx+ckK1Evly6Bav9L6sJ+G5NbCS0fwb0N87REVYqt3rPgxz3xuFjLqICuRFzEON+ptI8D145VATSTHxjCdJeqgUVTlfjaIQp7cjhmOXdbeOhejF6NkdkVUdKe17biu1dfYtWJFXtV2Y7qY4fL28OWHFrt4RVQwhzEtCPx3LU1OkRcfsrEoeRX2rkNLAeFZw75a6Uzek910XbeZx+6ds9yOf3cHwpZr8S6MJEV0YBhHeb7lYZuphqw/ewfRLU7A0N3pnhL3dVWCNutOtvhEymZdGhqM4RUWD3DyyGVnbIM/1PX1BnMrul4h+zprEEw52Y0isiKMB70wg9FBbEzrPzX11IC9HXIbeUCQZdWH+uEYrXcE1LsGKLeS743ZIyqGvdcfZBqhAHRnp+XILLZExZGbN8LczFMzFz+ybuqrj8zdR7rz97jniEyd7V/3TOpu6e1iq7Yd7YC6cR2NczHrj7Vhcg3k3A9p8Bzg9uLcv/t+r+VyAGiJLvked3al9Yf2dgfu7IV2CQ2U+VXRlO64emG5YCYMrhMI68YKBJdnq16hApxHZF73rNpwdj1cG4OIep0vnDaRPBMtIlKxpzqQGsS0A0jmvTwRay5pTUooPH8eW7dX2q2wnIPkMHWQqKjdVtsrEBnA5+CQkGuknQ8/u9MWGHORr+akJcTcA7+udnhEI4+9nwY3j8OzLH2M5aR/YaSm12fs5UGDq7G+QlQMc8rzP0HTUQeu+lU/MzDP06DUlCqyZgd700t8NBptIFs4bwC/mTqopnLJtpIg2W7l7wQPK44xaNvgY4KsGc4Nfp/y2BsI7S+xvpeakouXx0f5ep6TFPVARU0Pd4uY8b6m04fbxyAJLQUWSUJiIG73u11K/MNxGwvYYGSB0usYBjPhOWqgzpwCly0CwlJFuV3qB9gkVpys9DoWwpwEMCOiQrJBIumZxIfXGqjpvMZ9t+IcHgU1kbuPj48W9SBgX4QMQO8vD1/tvU9Pjx7hcGtjivocqOOA9ln9A0RIAPT3yIfQ9YhQeOS9llZJxKLjYkpn5Bts3P/98TGiMiArTLf1YtEesQeMIeGBrxkB4Cm/AOYzYsZXi8uFRTh5DQc9H3Y45tZSdr2jRsbL5evXh8vz07MRE0ithLGCTDCtEsgCgOmq70rhG9ShD7+tuWy4/WaRMOFhQdJG5EM9q0BvIAoFc646FbL/o+6tR5PhGuB3lpLKibKaAioItsnOEC6X701dR93vGjUI9UBgjPQxZ2ekHgPBGfUvxhUMAoWRTVkXt+7jkA0QMswOw5ostej4J1FxzWL5/P4XGAGteG0m+0TFf/qnx+J1nTUFuOhmMIzs/i4QMwHZ2MsGoqI8VxvfBtgrymE2/KTICEQrX10PxFQmU+mbuHGup2o+Yul9Aa+5kYBnoKgTjT2Ze7qbY/SmYqilrTQyEjjTcVdPqOmPTMUtvClkcM4KfQuSjofqObe+5jiNvmnO7c8cKCrprVwMhrrtzzDeSlFY2wCn1ERloMO8nSIquuPuGlDXQZSHGuXctPDGFcmQewqbf+1sjX6X9GgrwzT214NIpclNuVZgZz6na5jmtSKcvmG60RiggboWG32TM3YXdM7BqV3LtelW7zAo1wZ0GsH64BaFWRGMK6IiwZfxLdt+8PgxgRhX52+lPGox4qnvw5/yGtMcooXHyZXsz/yOfTB6f2NKPcGhx//5eg1gjkSqfg4TFaWZK6iogi7XwbdtL7gs67zydxEVej4J8hIB4noNRTfZ43LILqmfTP9tNgWGXfMgm/No7Tf9vp6LFgicdWyMueRi0wDOUVnT2Y5ZlsYdZtUyGfOxanyP2o62npV6ad6fOzk7A651z+hSP41qJ8dKAFHKwM83z/4eRMV27GZ5OKlrp2H42cDlR0aZtmD+cCnt67R5Xs9qwBbYa/R/bc4RmXJoazEcbnwsomGU6sBWWAzIPDJ7nuH1dd2IrImK60bQ2JVqT/7I+r42zyt56u7pRGbfal1L7Nl0VJa7upCjs/45ui5CH7unq1LvwBu3FuA8MuYV4ND7PzLee21viYp6k5/7zMZVhHt8z9nJAqXcw1hw1z1xzfYg6LM1FfU511Xfv6mQdaMH657WjXFNN7ynuzT+tU3zM8faC1UHei7fg0RFgIyLySIQ7LaRg5AEd9cza+lEPOWT5Ni8qRtByLOLgDlGwFCnrPenALidoDKdV36nXUabSmtiJcNoF8BGvEd565kb34+rCYkQpG0y0+E7y1Xv+fjtWh8g/CPPbsvIYFEHTfRbef5Ikow2W/QljtlZIF59D4wjMkHwLnxeo3pGrT/VwsD42aMz7ZPvQCQdPI2SngFSDH1EWhz7n8uJCBuRChIdgbeYLCOMbi6W9kn1F6yehARN42kve7+8vniNhrkOhguURWV7rQWdlwHGAwgH2YZ8/t+/PwVAbESFR/LQcx5y7F7nF4Dq9LCHbLPQdUhZplmrWTiqA63jTRVEtmfcsPg1xgHgPdr3gtRLr6/m+Y5xiJRIqnNaJgz3wnueRZYRkXFf0oZzlPEZnq/0ZNaGt7fLb7/9Zvo06lh4IW68N2s4kKAS+ZF1gOicrFTmIFQU3YG34n6LjBCRJSdiXydoy5eHL0ZQfPO0VXj2g3v7MxWVIjZeLCk4FyDXtLSC/AwpoyQ3rdeIkLkB2USyRHpAtTzuPEMJ1wPvVV0SrQ3pDTuv2fyzrgOInG/fvpo+MwLBdA/lxMZHa8zltepOtUPrkCrKz5FObiV+yrM0v1dkHOQeDtPrzC6cZ+prEC+mayxaB7ViSORSpjONVd1TPomKZpP6/PhXGoHclWkIXImo+KdHLlI3hkJvIyeaeb9OHpdlE14acQFIc0x0WOOGE6qpGJx8YH1WzaOonIyz8YnrBRZBCXeHilr4BhstciLyM5m949xtjMgwktJAkJEAhaGQvJUXtYyUUHJiRzbgmg6eDK0bxrw2LwB3fsiiUT6m2gAGo7BEeRjhMXp/bImKrB+RQlEPxSQqnKvxlk2HaPvTQw9FShVAryp3vaNAhBkGqd2n9F9dnAEr2UAKAbStwUMaN4eA7ZnfJzYBz6WX+EGi4sjhkeuinBA0r6OdOqyJHIYxxVj9nBzFePLQscEM3klNDceHPQ+dzQEx75zJlXqY1LwM11wlAUojN6eoJCo4ztQulKN6GmH79nCuCgJlojKJ9PZgNR6OV6e740RFCFx0dZtSRPougYYr4GQDjk9TPq0maWi1vRYGYwHF2m8RFfgsYcU+pqKO0jWSQvO1Htm+Fy1R4aTq0FYjKlxudokKnw9ce7ttkdLfsc2cl+Gg3hEViwM7D1/b/lHH7hAV9g4VWcQp2iztck/4fnMtbFZ/fSefpWa4yT00St+mrh4jCK+BX0f1Ise02grZjFGeylqtiqb0BAdz6b9egn7smz+FqBh0JOyVNZHJbq9BoFWv2nH9CEP4Y8O2uTvAPu+7wLHVa4ZDWd0umjZ1I9TZjJ2s/n2IilHfjGRFfndsylbalDKT+8tR0mOlo+a0eZLH7r3rCbqmOzpZXn++fscRV4D5zmvyMbdbaTG4H+yD4nvLR+s0AOKanmO68Zpe7drxkTHv2nycqHCA1T1FQ0pMSSv9CdPP4IdFaWnhMZc472Cf2JrV+uDe6bvYIIoiMrIne0TC3hjFGc1tIdMxxdCd089W3Vvn197feM3VCFY5WljLF3Y+PxdJU3Kn+/UWre+AI8Fbpkjp9g9Z14NNgHO2Dx37K93h0RbTss/xW2vg2cYd9qfy4tU8iORAMwBYkqjguc+67Dn2VxqpjXPzMxA9uHkWzmgCAp3moOhANmsMwKNZ+fi9SLkfkCOdXkQHbImKsKccqoljvAu4sAb8qZRaApdB5IWBU2SiRi3T0xqkhqdy8rUWw4vnWmofFFL2wulW8Pf18u6pnwLsRS2QFxIXBH79BwQFyB2MixcAlpwAgP/+x3fWLShF4dVGIyqsFgPTkEnnDXqrRDihLgIiE+htTvnLgtSMECDsRWwGwDRkH+0I0gcYUETJJKGG5xHTYbpwAt+8T3+LwKsOsGgIC3nzWpAosN1F9GGh1LoXTFX2Yu+SF7/eE0WebS4MlYusHZof1a4wAqjUXlD/akSG9geREaZXvW/4zgBwr32iebVrnNhEe6wfcgqOKDcSCIik+P790QgZ6mymKWK6Mq40jAvm49VJCFtbop2NKPNU6BY5x/bAcjcMx8cuHMNc9qytwvFKqvEqP5o39peyIVzo+fmJqbiwx9xmhoAQ6WJg5ZmH39o7AjN1vE7z4H2XHnK1zFRpXmfC+reTgr6e+avsQR7w3MfHJ88YcmMEVsiWjrafNSpyg//87VcdgQTsjhAV/+mfvnPJBQjuIJ/VhACLSaWlzcoWTjEYN0bju8DuBNBNXTlowEO34hOURN8VxcJzYm+UpYSPHovSKB2JkXiOwluLkUAjSQbg1rBbp1dKgmb09r12KJQXs6zBNPBs/Au7v+lzWI51xFZgUhr7vLIcWn2jDaO3gGjheRDAHDfR8Wc2AQWmyVysVq67tuwBrJOXpWS0HgJMN7uMch59xD1MNXfEcVzUx/i0RArZnE9THeCkxrn0fiV/VaZWMixnyvGgZdvadHkdY4Gi+mz6bu/W8tQw/DW+/m/nLZWebuO6GYGb7fhSZ2julf+1Ad1Eqnr0kYzNFDHoiq0Hgh1IPeuEHSxiDOrYrHLfeg7JmdCYiJTt/Jg5tpyjIPA2k5sTk8+TR37mH9ZDA7Qrb2GO5pHsHQ7ZsY4kI9f2Jx3a+UytnZxTGW95YnyLSClfZQEqNp5lpQkR72SHQQe4InLA95yjirzKcmwz49oIIKPqqFqjIsZLRdjTHI21DlLWHjufwOu7VofwdUfq4SvWIOb1dgbmZ9261bOsrTGtJXtt3pszd00Wlhpq+JAyua1/tKfn6iiExjpDVO5v/h/p1E+/J/3Cpp0w6nLl3O0ln7Gxwj04zPg+xgPR6g1ljS+88o94gscBdrHj1J6sQCLdu5SaYwh63Fp1WoT3X2nTasWtds7Qp82sXwOi17d1b19fvSYIqXuX9UUae+jksHpjtOfOe/C5ZXD+3R9Q5E2TzgLq3fUrNX5tFLpeVL16tn3dO3/Wc6716dr3Z9vB41FjOTa6HsCRpawA6OWg7+3NXZLpk04z2Gqx7AS0KyXw6GHO2dvK7kggXbPTNV5rsDxtMnvOTq3ECspbWhaPLAHQ1HnG780Vzyhb4NsiSW/gDc3xFGgogNXAyUilIrvLa1RKa+wseHk94xyP5xOAk37Ztpj7Wt8TAYssCEzv/r01Ms6Dn2VruuNCVGgswp52tZs5EKY9O/LGl/1VqrptFnUsUrGwEPjt5fnl+XJrACJy5t8zHc/z86ZbOcw8b4pUUN55kynVWZR8FYaOkQpK35OybnUOHDhnaqdbq40gUzgJBv6GzBAEfm8L6Hlj5KCRFYUcNI/+11f39Pa1BID/5ZWgu3uKax5HsJjgswB3tA33WZFo72sF3ldygP7S4x31Ke7tErtHxaQvdwY8m9i9vXMu7m4vXywd0VMSFuaNzrYwkuFiBIilDSr4j2x2FeKu8hf2vEUlZLoo3l69DnOczIZ+e7VID4tkuWUUEImeO48iQ8YPzgfAadZZ8DPT7S1TSOF+L85tURuuS62WhDvxWrowH1eNpdqsovVV/3W6H59Lf9SxNogkzo7u0Gw4VUZsol+oPQL5fn1/tQLcRmo41neP9fLMMceawdhYf3xPMTla6KPAaDjTISpK7VXrpI5gzrgvdA5cImpMXzqZkw7HOa5yhJZMq36KqY1od2czunKZBF3Ob7P8i5ire4k2OZsLI9/eLp8RFXs75+d3v8gI+KI9WKMCqZ+4EYUq8zzi/JvghJQBD9GzIg89YeuOBkcY846bJNjJDxia6TnrBCpf9fzMIa6H5SPHotkgVWHrALdLLYhZEUSIez1EBiiU41ZaN/Sk84obBMaeNwJPFdiwNtV6FPVmgXWmycaaEzFO9h3Zas63bmJIHT8k022zrc+iVokUfAXptiLP+0xtjl+6a9QIbruibvT48HE59ETbIlUU++wtY3qyQQhLU+pDJThuaMcrSs2ktMHrjfEmHzc3UmIejqmCeP0h8G4beTSO8YoAWK8MylKRrp9KVJTDT0RicJ5t7pu+ysMm5s29YnKd4xnpYZ4y4PN+415NU0SRjJgtqVKIigDMx0WVa2VebD1RkVpzLXMrosK07IYgGRcFD3SVKMrUd6kbFkqhEUUaPQlkrYiKjKjg/DHPZ+mh/mgOtgEE1num9gx6/Igin+7vIipcXaYe8jYE7NsQFSQpXH84ob4xZhVdVUiBsVnrjlSioupYHQYHvTw8e1Ja9ucsg9s0cPY8l63TAFQx/hPUbvaWHXU3v3cP5L6mNQd1rYsP6c5rT/7497tERWnbHklhssBd1/ZiemNpzf05REUOX7P5qk3N2u7m8bScFfL1H4OoOCcrjSb4uxMV1D2StH7OV707O6db3XRkzNZtOv/u5l0Cdhdfd9tON0q6/oxuW/dju8cfGak/85q98f5pc+HepUZYWGFRpKTZ2kCSVrz3zYj5aZd1ec6znczLOZqlnkdqNFEZ/w6cL59XORFxwnMHD7xmTzUxCvbdG73icQ2L5jKFR5/Cp5NlRkjau8NZRF79tO0BcsJeS89jtoyplegRL/tMZyfTETRMehFT/URPr4l7AcTzWfN9GOsdXePHP6U0sSWqFECrdap2DXNC72SAvZa6RVElnmUhSQoZgO8Xq8yx6GKN0pj3t072NQe4HqC4RViYg58TQkgx5OlaZvtPca5s2S1TVZmzAjMrWG2QKKLrZ0wQBSZn8K7W2JZi615LAuA7POsNBLeCyPiXgPzw8470MveWmghDgtRI9Ny+v7y8vdCz3dMDmWi8svgwUv7cXu4uViMB0QpODKBPKm6OKBcDzSP1db4ZYmvpbTBeAxCcXvUrITTg2FNuaTxv4GDpKY8sbZUXiMfcPL8+X75AxzjYbrJqNTdIYjx8ebg8fH24PH4nDob6DngYyADVZogIkiltU4D+KnaMvt4xCiBqYdzeesSPpxcqaawiIwjm9O3N6l8ohZSdt4ycoNf80wv6cR+EDMZdP0i7lKmn6GFf5TXMUNUYwbOjDkymT+9WqpGpkCGkggIRghe7fNp7SrSP0ohJpyhtkyJwlHZKNWW+fnmwdWsRJp7aCrKF/uEzzMOwVn3t672zjFh6RK//gX8xhqoJUqTPZBzfI6JiTolOFShMjOPDVO+sHcI+UH6VWpzkIucssnns6dGdTZw6czsbQVQ4MWc6quB0kqdPouLPtJA+n/2TRsAX2EGi4j//sxReRVnTO0QHbIY3MlqiAgZkkkvTS42KwLECRHSg7d2JikC9BAy5sXflHLU6JF/DuMT8JjhnZkEYb6acomAWnzYYgUtPt9rQ8Xc+Ib1eras5Neu5Lp0IYCPsqzSIh9DOmDZd6KC9vbDO6cLzyb4uRAWZEGe7PdAmjCE1eX9yqODnOgh+CFHBrgiD0xxcmT2XkzTLfCNRFITImSC8kikjuz8M7GLs+7orOQ8UfIWvuoDEsxRLMpJSJlXLuY41tAO0DXK+NPgLITNEuuRBZvXy4TBVxraPqKDX1NZ459NXfc4x1wH0OFHBAxMOdrWoL2Z/S1QoxL+mfrKVQmsqCZJFO0OXDXNAKZMhMvZvT0UXObNDd7m2/H6UqKj6h4ZTjajwo40/DAYexyFfdAS/zWcyei4BGI5dEhXsiwL/hzWhxi2GZiYq9NTQJJtGXlH8i3fU1RVzHhad9F/e2BEVeUWSFIr8WxEVI4E2Nmxl+Jqm9YP03A2rZVTFJXS3xqOOS63JUu/aEhU8pI9rYE+C63fqc5IUnD2t6y6ScPX8vOf8/I5t4l/DU44I+tFOf+C6lqioRM/i0LEcJycqmNeXVyitxHh96qiVq3G3m3ZgS0s67KztHyGchjktjhN1f/+IpHT97p51zWb8gDhsblm/o7MbbcCb155vbSUm8kw77hOj3lm/WvV+jo9HZ0nsPWE9S2fB8VaWDQzft8Xm1nXP6oDlI2ti7M+2z2f7e3xOfuzKAIBPPKYdDwfgAPJYQVYHDrtznXnut9URfFoLsMQmrkBzpY1anO+6fi1kxu52G3Wly9a6vWQndTLa0sw4cbG8pyVPCGjHSpbXvffaUqu4d62A/5ruxSxpeG8DuC73iqioBEi3TwkExHNRlHZNVKCd5RxaHkagkR7liiSwWdshKoaIlcnzCONh0R3y8gYRY8VrPfrX3y0yqU2FWcENtbdEbKx0hBFplmqKaRpNjo2cYH1EZA99vdBD3rZ4mmThzGhawGSChXEFClv0wmI8eLRJh1EDS/1HgDf+VcFjFaim/T7XryAxgLHDPFb9wx4xBZudey1FDsiggAkYEeFplSx64/bG3gsyA88zguTlxSN8AO4yxVO2Gc/L5LtKqbRnq2S9C0ZTKDUmPoc+ATAN4uXrt68kTayYM1JF0UZWmjCSh+9Gunz/zvRUTI92uTw7SYT2ZD261CkVG8IzVdA4ozw4dubY6wC2yabXQZAzpa1jr3eCNEpGOFwujCp4fWUaKYDqnv5PEQ2qf4F7RajgPgDqrMNA7TCbx2kTUGBItjB9VmsnOUGDscHcoi0cF861pTECIYM0Wf5mA/dB3j0/B6FKgo1jor1Y+Ay+QUqrp2fUycBZlJFCJidVlV8hKqA/IvrEI0vQT6VHErmk/eyaVSU5VConES3SH7UeisgXq+nhuiycZheKdCSTcvQ7ncmHFoI6sDofV69b8UlUdJv55+e/0Aj40jtIVPzLvwFRQc+HBPdMhTFfn7PEDFeVF6+UHD7ixhVe9GXla0MzENH0pmATkgJiWQmIEbS2TaiQISvDYG087U9BJSp45ZaooBJwrwZrrue7hJfCJlf57OE+qnkzmRKNnhonE7NYRVJAQS4sbqnkiT/cnHtnVDQeW3LfC2jcnFMzigIbRPwojHnavQRS7oIhgQ+KMCgPQZomD+9lDsc5XVTpdwhQAadmrx+Beils8YBoaxxi9NXk39r0kTu5ZN0LIjVzaltFPGcCFlebVJnLleRugNDFgKd8pue0t9Znu5mlMq7DuxtLZbw8rOyp2ZP8O2HFdadiUh0M47rHZVNEnLwycmBXOfsdFJlSH41w5vb0oSWjQ2eOWxIveRa6Zs5IUDxCYSYIK2gZw5RjsvKesCeWqBe0gPOgGjEpw9KZId0jkrtUjLgkD5cl3UywqZ6GbnhWGYeqc5oDtVIEcnRG+ViDGOfhSd9WckPSorU25fP0vsgsMEVU5NgxKo0nXIxB7YVfVUnBDYG4o8+aNY+QaM13TlaNkBr1CUmpWZGPhu5mfI+IcFW9paYUnzzPzf5czQe5pRCe/HCzdf3FJAWav0dUVJkPfbMzD5GqM9I/6Tw33+QzYqp4Ow9Hpro7JM1TsgIMjgCyR6e2gmLzznJWG3T9bg/gRxv5A9et21RbNLdub/aOzGw2diQqOLod9kn9s+7oWfA8nFVOjdv65Wff3RIVAMPaWgDbhlprmgGpRMVH1kJ14jg1RNXT8+yNP3j9zyUqKMcGcn/x4rc7oo0deLELJ5nrREfs4avtquxfyWlQ5tLOXAzSvGBcJrgDbxu9B/LT0zpz/NOjfFs7Tq3Yk30B/TEIfna1HSnqKBDks/RaXjBWe6jVJUC6mELpaAXasxvZV58z9VOt8LYaD7elpqFNAFDODx7hHP3o52J4i5EdjBpA2xDRINkKsNYfpTk7q1PoP7AW0Po5ZBnAPdpiNRlUGFjFnadaU7TpaUEATEc/rO3uva7IAILgHOcgC1CIOorS1wLyTC2E9//xx3fzSLc0awDrS0H6aDec/NwpDIWIlZYV7eCYjvVOgBbIs/7tFYWfWZdB18vXsaYEY60OXgMQHSC8gekGtHrEhXvV46zYEcG5Lvxs5FErmBoByYgEkRc95wARIIzsUD0IPofRSBbVhIgLFL/2YsWWAssJhDg3xFjz7mrfKoKkpodSTYKSSSyaAAAgAElEQVR6XkMb4fGPqARER5gTitrlMoPUSHgOIj0AUT0/Ptu/Ni6eyk39EIFi5IFSMAUJsC7cLuxFgD0LOqugdL8HG/EAosJTS9n9hRRggXmvDeNrRX20FH+WRYVaHPdZBJSiYzz6CevnEbUjLA3cjRclfzlFVAjIV8o7kZs1ekWyX4nZWdts8UKSObY2LYIMBC1lX+tQuAVTr/Fa4R+r7be3wXci0QohH/54TvjG/vdZo2I13J+f/Voj4BvqUaLi32buxPFgDWY2wwDJgDvoSOsulGPdw7f7uRUQoHIHM+xpn1ixPtNsUGlww7U8mItBXR0KgiG9MgmmMKAAI3xPRAUNOZEU2sR8O/Kngqjg5jZ+jr86QKkDdjqDx5DDzeMHsF3eIUpTBU01vGZ+ZyEhwrDO9/PZ5R43pOKQZkWNqndcRr5sx4Gf6Hp7dqmBoJBAI8VkuJlhJtBtnMA6StFCGc++SbrF4CDoRIqUBwyz5g+rsj4fOAZQNV+eolGMeNssRt8YNcv+bYGBhU0gWY4NZwCD84ZKYuRmx7nmdw5KtN6ZOdaDNF5FhuoF27UwgpOZqoj5Rz0qYG+d+ilKRbKYaqi8s9SoyM8ln5oFkqn1Ph6y12cv68VM9HkblYokvCe0PJvoquTDRpBf3m/jq/yaAnbOhovWoc1mqnX7PcOpRe6u5qMf7EoGYXIYRr5OHxSCf1U+Pr4TyqA//QS1qa5JTyko8a+y0BEVeXsdBxIV25+9cYI89YfaeQ8zQ9eJCsoH16/2ya2eVfTMai/iYHBu9Vtok1NDGxEVcVemGpvbFHuwC+lq/dWXj3pi26zVPm+61C/NiB6XzD309VSvz1/cERVjf8fnds1dERXcQ2Z58nk2xXBiUU5syVpKx7Z2T+/uPdEae5EO65RW30u9kOMSLNuZ65/VpiPjclRS1s8SMb8yAnbsw6Mvjet+Vo2KcyPyM4mKs13uAEWO9LYfu6qjAydDD022wxU9VN+egLa37E/SYadB2Z0B/1nPQvoYK1jr/zKSva6FcV2QqNjuwwnUOIhr+q2CttIqI7Aoh4+6b7V6q85LdbSbiIpre5p2YxIVrBsQOeSbMd+roUOiIodNxEV8pJz97igUnuwAqwE63t9nSpSyb5uMXmEzAaorasPSncx2eukPHCBXj5P8cw48/34Ux230zfQgXUWvdILVitAw4H/yKOeQrdM+qcnDWbDWvuhYXK+r8fT0ZKl7rF8gn9yx04azpGoZ1pD3p7q2aPxFFikHfkRWutDjuiiEjBoUiCJ4YX5/jCmKRysdEIkBAN6LugnW8Rtbi1iCr6/EdcwzHwD/7e3lHuSP5skHnYC1R4+gRsfd3eXx6cmOEA8PX2xfD3IsosEv5mH/8PXr5fnpyckFRlTgWWgv1gUjjVapjDlL1dGRESiMzsF4gNwxssrPgIgmQcSECBg5yKId+Bxe8FagG2MksuAJ393bs9AmFu5e17ZRqh9Gz1wYXWSpgQTEv0ZaLXyHaxiFxOgEDKeIDp3pVG/CdArk6f7u8vSIsaUNDgJAc4v7bdy8zgXmmlEcnM/wO5Njq9etQPswNorexZh3drfkDG1WZALl008qaJc5oL7Z9xYNYnOJVEmYFxKmRiSiwDnSkilCBAXp8RlqqmBMvK6Loi9QZP1MREUeB/mb2mRt8cgnfK731/ofVQ1XMkPXhy1u60SRQeyz9jNMmRyw0W7N7UrF13eMeMVaZ9Zn8IzlGWiwf6pGCqLKPomKs2bj5/V//xFIRCsOvgbUgZV/ubwjpO31+fL28nh5ff5++RcnKmjj+TI3jz4oFIZ5QcGaslG+a9M6cwQGe7ohLcw6SG8AhXpBgYDBt5DCeG6mflqZKlzMaZ3RdvDcjVcG2oA4RUg4Oy7wcvBML7UqEjyrRMVo0kbhVd/w0+DRbwSerKUiYJZ2mBc+sxAJ9tG750reRpdRHviCaV03jq4JUpl6Hcx/GmEzhEVQix4bnnIigN5qhOKqTEkxAiS5I2oDi5A3N+7NiLDNmwY65JEeI9mmYaPwP2K0q6FYiAqTCQ+pzQErT5rOQAPIVeahGqh13LdgSc7/AIBKLpHmzHPYz+thI6JFlLYHnRINUwwOypHLUyluqxy/a6JiPgiOLYlh6Izxjfc2ZZE/YRpU564AeGWwxaY6yH4OQP24FqgaolSKwEd+VlvEKUP0ANoeO3Uwmg/bpp40nils1rMwlt0zSvMZ6aZiGPd1ArPi8oBU22a6o4CHAj3RRhWXoywWw6XkQZZ+YkRFHcH22J0t9ktSB+IDESzjgcY1O/X7FT2793V3mM/PP/DwtExdGvkBD3xztNkqPoKyE/PCELUrDZkPUfX6mq6sPsYLnQ0kpxvTZVQrSZpAxfz8qjPrd0X2bQDW6yu/6fu5ISqU3zY2eO1p3gdLfcA3hn6aDndVd3EtraWpOzBFf6redE+tD0jOT7nlHFFBRX6VqLAxzL32ZxEVw2FIymxnTUv3bAZKgM9iBK+tnPmWeRcxyd4jKkq7u2fNn3+0TT9DQBoJH1VM2N1tQpIPKt5zREWPT57V+ueu/5kY/T5R0c3our17hX252RQb3Rxw9lNe7Y3KzxyD2sufRS60I/eBhr8bOOWAHlIUOTDZPcoS1txkahLtM7jeAEiLGgC4Sm9683AtDwv7os4RzriqQeVA8tIRTc/xQ4Fp8HC6yTQc14gKEQtquwAsnX9X47tHVGj/jPd6YV59bs45JW2QeTF7rnnTrw46ytYOWQ7baS2tKHj7jPQsDsLhF4Loay1rgOPyUWEtRO0EpfDZCe0ahml+rKV/8r2DUdxaj7nv7hEVM0lRU01NwRDRjpdnALOoC/Bm/z49PUcqHoDHctAisOgAchmQ6gTFlEQ3BvQaoSUCSE6hAHeR6eKNNQiMJLq8XR4evhopALn/7du3y+9//G7tg+c9alVYZAGepzov9dxr4C3/s6L0Ni10SGUKIf7Q2YtFrO3vy+Xy9eGrperBd/jd6lV8IRBNj/N7W5cGbrstDlLg27dvJkMsFs26B/pBBAiiUsz7fiU3XrjbUmXdY7176jBPZxbRDQDK7x/sXIT2sWAzC1aDSPnjjz/slRhrvP9f/e1vFoHC2i2Um1ibDsgzvRfGgCSEIlFIPhC4xrixcLrqhnjaJrfpSKjwWoD5eIa900nbtNlZwBrjZkW/3a5W1BDqa7CRWcgbdTZ++9tv1jbWZfBLNGEO3FuKppuLyyovEjnElVJbQbAfY6gi2EZs2Vrj55YazPc+9AXz/vT0GGQA2gM9AyILqblMLznxRXIK6blYowPyAf1qtS082uMMUVH3YJ3fNf9KT4X+isAI+7OcVer5RdE5tn7dsVbjYfilr020HWm67Eeq8B1rEGRXpmarCqzuzWGbG7a10pnCWzk745mZUWWh8z+JimGf+PzjlxwBX3oHIyr+j3+LRUSlys0IGxZD5rhRzAbIbJyVvNWzh35uc9ruNp4zwSrGBmiuEdP1uTjDmHAkir29aR0LlwaUp0vSQcTy/21AnVKrwd5BhlqkinaB/iCgQuGrMQx0rbyX4H2OdkZLmLeDnLciHUwtaq6BNpiogKFuVNhEmjWf7wuwW6Bec1gzTyY80+fAnz/mLZbxIt+QmhuRbZrnOTvUp0qZPWdjF5i8p/V5GqFFkZts+/j4vzVKpQfLOOAs0aFxzPNPJQs4uhkCbZtaledN/Qhdr3kbo3JEwI0yyfyiozStQMoSmaTrI09rlQeNEU0T88CwzhYJ9IH7kcNujhPXkAoHRx5GCz2mJ0oYpko7VoLrB4Df836G1Gte49/sg9re9sHIwzTPJqfjpYaP+ZWHHR16BtJV7iz0GMbc1RB5Sew43pX0uQ6WF4sSOUbtPZQO4+58HvPgJkLXZagD4+3wX4kS10PuFVWJZbyNath1R4mgwuNl8M/AczsXLguh6yTtRefVCdFBwboS7yY5W/PY1ntsFkIPFL1Q1d8wNup/HmNlnG4AdSeZ8yhXV+u8j+bfNneLdbcUPk+VV8Pph8g4E+VR/sXl6nkmq+5YGOBAUuN22QoylZNBSO+sWJcNbvaVIjMutaHe68GktoP5iD1NZBnOCPP2wxyj+SiXHfjViv8emrjoXxfQcBa/q9EU1RNUROJqaMchpA7j9bOspZyvvpF50Ci77cd7REXz7tz/y+OuEoLrFTBMan3GycneB7V9PL0JseZXMlBIt5GILsqm6cr8MTNUb61uXQczrM7hvrh23zby0Q732ZoTa4Qp94qVt2zTptWc2tSkPXRsaM/1uRKKg4/MXPMskA62ou6H11VJM04TGVz7l/bJeO+efbOnO+bv9kaptwOv97S+Z1c3ypRwWxS63QiJQoIT5JojJ8aeqB8z6NadcqoT10Dwxw3zyPiZah7AHYf9jsyQt7y+N3DfvcPXc9ftqeuVEHvLSnfJ8UXOafI6bnRzWsokhzA35lGss0LRl7vrci+woXRv3v+tWLVHhQDsxfeRrijscXrXK4ODrcsqdI4dbKZuiqAw5yqP/veD4HIvlAc9vkRbPLZ92X2TW9fxWVuBALqBpx6tQl2SMh4R0E5ImcNfEDHTq7xwtOo9GCgOkN7IKe4wBNW9/kSzICGPJEVY+0DkgdafFB6nizYsgt6VHgd/A7QHngRgHZEZrGNxZ3MDkuOL1ah5s+9/++03ps5ScW2vUQCnWas/YYD2S9ZncVuXumC2e9wKV10Ey9/P9OX4Mc//e5AUaJ8X43Y5VqootAvXkIwjGRH7sDuSUK64KkjK8exkOssLKyNKhWmu6fymVE3d+hChpRRYRlR42qTcZEQoEAeSdtI7bW2CxsJYGglFUgcEAGp3IArFokq+fGEdjMCDMiOBdKwivyx1lY8RZTh1otJmYe5tvp+dlHAgH5/j3SDNjEBwG1LEAp6m1FnKcGLufS6b0juXcDJ2B2fpG/9XZ79Y74El5Dm16mH0RyQJo0WIf6oAN1OmUcKNeCyOUfaOAhjEvCEy58uXaPu8b2r9bM7F6ou1gynWpAeGMxGhvCDp7EyubCg4+nwSFbtbz+eXv8QI+C5/kKj4l39DZhYbl3KrYf3RY1n/ZccMkJXyiPzzteMLU7ejxsOw1ybj6g+K/tq5wp+pY93SdGvP685Cl5RUdH2IbYgKYnhohqce8j4hepYDY7/mO1JJ6TqMazkQFkMx8lPqcW6QRaaoeI2epU0k359KlZ/lLVk4fSu+eE7pt8uDbRqxQY93VSCQ37BNdtCvb742v+NU+J1ufDREBeeMm8d4KCge00Pn1ws2CSzBhzmuE6ToaVbMXA6gmK/wfvuGPhNmGcrO6wQyV4HJe2B0cBMd544py7iRjimPOA4pwPVZkm2OURpZFRxvwa5pyFbTOK/FYs7Qq8cu8Hd7OieLrokbCyjs7wtw2X/JXJsuZSETW00Qxs7i8JXHTY7hnO5pJSGpF7Jn8LKR8cZn6DtfQ/Jm0gPDc38eQf/73Nm/JEZYExXiYkicJJEx94+HI9pfowxQd1USQ0oyPY+KlJvHUdUd+aZrREXi3/P+M41VFBarMlCv2UrnWDejCFdV9mG0e7RN+U7TQnW+lv7x01Da7cqpqdPrmC/HyR43giTXiArogVm/oEu2z8/71ELv5kc1/L3I/hXA+SrROevzunQqaRJ2h0cVesPCi0oE8XT/ag13Td4F0dbbxdJWOfscabxKUkhPN6/1KC0u1tBbfXrx7jH76aNWA/WBiIph3YRAHTUCpqafHdxmsveIiqp+6/7R7XciMjbL58ramCdFRMWwz5eL/hqiotuMznyeqVY3NEzYA1sRXb/BldfgatmL9/VvFm+peenLfmDg5ah+ffPhP/akxX6xbsPCSWc4+ByxrmjzdvZab0Y03+zYHX82URFj64SzDaWBlm73i4iW9+tZPVAdGOqEmNc11ODU+d25WAkBBaAbQvaP31aMy9KueFpkypDL9w3BzfnnaqTPrC67FtXoXE/FolROHcMvMNacdcIWpwNByL+/P+RlFuNhgMYvE2DUeprnhE5VeDeiQsy6Ri2FyPzLBco0QEmIbmS3lfMxTSyJCjlxDULj8+hpfqz+iHvLmx2yTl3UERU27t5mpakRUQFHRciHRSjAW/71xQD9G3mcz/NdomusXoan1mEBdUYrqOh3JUNmOUvg1QF+2V9OUIUga75Nrmlhq4YJ3odoC3mVC+hWMXctMZAXiPj5/ff/1+79ghoN5lnPtEsGHLvDJMbCfnRUsqWoCt9b+1/vEKEmIFzzpVoDNY0TPOHxWEU1ZHSOv9ozW2A+rVC3QGUjKpA1gjKICJG3FxBQSBH0wr+diFmubSeZ8J3qnGCub+9nWWY/lYJINRjwGbA7jDMxCV7HuXTd8/Z+ebEIoC8RifPN0nERC6QjHn+w3u39KKRutU641tHvF08vZcC7PxtjYamfvA4Fo3Jw7+3l7UWRQDwXmpwLs/HIHsijEX2ItBNRUW0oJ65FjA1j6CSrxgJjALmAXNm6w7oo51qMB6PjsL5Y9N3a5ZFnKWSekl7OiBWbm9ce3uNEhYgmXDJjEPhbxAwjXDimJJZcp1iqtslpjDAF59XJM9Y68r0Cc/dJVKyW1udnv9YI+A58kKj4r/8rlB1Yaio4SzkQOa7LbhCbESBWpLfxxeILRrh1TXsT9lEU05Yl78rTQ2/5FuXVhvI4cIAdDgNNQbIN2FZmqnhA0wEzi9TKMB7ndQLd1MbWWCbZUqMCMDZ5YM+aCux7ISrKwciUXGlIwF7YeMoXCUQp5ydBvur9wMs19mPv+gOh5zqMw8M+eJgQ82QwxDiNdTX6A9bYoiG6YAa2Sr9CDmN+MnpheNceWBsAaEYdiJipz6hzK1BWspyb3HYNmQFQZnUkrXSnjDEV92X6oBhVBxgDk/PhCoLGHrOaVT9QhAeK/ka0Qxo1kg580h68rGuLtVq8GMb2Qnco56TLkYgK8whIhDHeWR7fgbjz53OT9g7ynIv8OUJUwMOnHjh4KGE4LFe8SCM+14zcIew6VvE0fqWzJw/hisVS3zOigsZqeGT5wKqf8941EBXhme79KOcBeXBsDrRFd+ngf5T02nS5gugNMcq59V7Eu8v4Th1cRQrYA/TyHd272eebfcpj6RZau66q/DoJ5+bQPr+4pDpLHVRlJ38PA/nWLVx/lr3zJxEVVAP9nn2GqNg8qygfrqNtarcNUbGZqO0HXXNPLjuu7wPmyrUmTeLnemP/LoEMpkmHVFHr+9op2uvAyYHawTmtUcNQHbHzVl1pgOB2Gn6wD0eIitrMH+nja1PfRh/bXNc1sbM/X5O5o9+fB6hXUjBHSc+KeT17vV3aAMVHOxXX7RQYn8jrYZuZG7aqwXVFmZCmmIHYyW7e9Ge8fs8Jw3RTOx7NN9cW8OJ55+Wjn6TUg7JLfX7CvlU6HZFV5yZ8mU7p70RUsKUpbzqzMVe8avoxInpvY9k5cq4HoyOW3cnJQP8CvF5NYVY2K4GaNq4iYUorlvbWIGPbdT+TFT5qkToJ3yvHvIF7Do5XgJX2ef4cISpWR3p7DmqICRyPR7LdBL+ZwojFpwkwA5xeb13riIrwnkchdNQP8PROiooAWIyiz1YDweoy4Ly2nm4QN/DoNsLmlQXr8TwDZo1E4Bkc7QURoBRV89PkjQ+QWTgCnmf7+GJP1VzgvSroDpPt4euD1ViAeFi0gjvGwp57enm2lD82x54+FNdlXQimZ1LUytsbwGQpA18mthXsExUE0knoWjQJUlK9vNiYWEF7TyOHsUGUBcH3N0uPZHU/PLVcOJR4/ylXJCWy7iqGF1EglA1ZPYwoQF84F5186DjCrCb0lp9Tj41bE0kIrQu7x19rxJSIUGRN8aiSu1ukK2OECOYKJMW9iL1CVBgh4cXdLQW86yqLjPlyf/n+x3c7PoFYwpghOoMEBF069Q4r6O7vs3f6ey1lmdXHYDuUFgq/G0mCKJYqa4uIChtJrfcSEQYCCvfiHSSHOOIiuoKUNZnY1gyCXKBtA7FU6sOqpoh0t6Xyiqw0JHVqxIUvnCK0+nW2AQoZQeXH9eF9I0nrOK0cVcsjPomKtV78/PSXGgFJdfHM2KlR8V//HTd6ecoaCDf0ZwJPbjLU0uAvbOBvDsBbeYWMhvBsQdwgWNbCVxw3SgNB/WXG0hbmcanEm3HubetmJ7cXc3yiD8XuDRBueF/VBNeRibii1CuoBBDzo+aGPx9aujcMoGxpX/WqFWAqokJKziIbKlhQLLP2QDhFVAgYy+sn+VjOkYDAJCkqyN/PNd8yX1vzgm8iBXR9Se9VPQvGIJfmcEzbwze0PDCFd0JEGvn9Jugrw3QLmOoZrxYhYb4G0f0x6mLKlW8Lxd+RyGx4P8yGj81zdeqJCWObYCdVgMsMtZKrv45Mt77smh2iIp4R14iosDd73/X7NBf2Z1Izs2HcH9AzNd0sV0vj2t8iOzeu6ZXK5RZF0cJAyBU1HrJr+rMZkGjAiOGdOw1YLJhK7lY5yggIynT8vbNn2ajXeS2yI0OdHlPlgDDoIql5X78HAcnhAD6RDtIEm2Y7eJ2fc2zlcTJfvzzcafL94lb2D/Zjq1XmT/xv6xQ9h7qD36a/vi5ybemK8o4p9RM9cKYnOWnuo7WdvQVgSjJfwlDGeUeWcu+ZLtoZS6VESMDG5cnHaSCtuZGvf0ZO/Eorz38tmez3zvPP5B00UK6RJhhCAUSVqDj/VurgUz/XGjeL22JtHUpvt9eoCYxqe/CDRMVihQ2tqvO/3fNOjSq9COetsJqedaW66J/bKc61p12/9pjuzavP94iKGs18oH12mHAj7cDl7MOuIC2/DM917UVVn8zPWxEVemrz8p9BVFztfrMo+vHYy8mzftvPJCpirbnxamDPkBIy7fEhLGFuWtPBNVFBEOjPjqhgE0dtAdGi1zht6XFvW09eG1HRKcArRIXqoe2v9Vmhc3cWyQHwNXo2EBYLqmJYO00f6/yV61W3QcC5HIY0r6vIjrlf3TClc490i+ydFSkgOaR8oj2WbsrrHqB2xeqnOjjV1E+DaHjBZbRH3tYCS6tNVJ3d6rsy9ZIXWr4nKO0zFqSY1fTw6JRlWz3tleYY/zI91ZqEIdfG6AeMoGovJACNFEZcAzbW7oNnYDpqaDjBYqnHPSqERIIKP+P9AK4JJoVTntLAGcI/zq7NpL9TNo4c10QISD5MtszGZWFneebjX9ROkLMXro/2Iz3Uw8MFxdTxA1Lj+/fvdr5GVAaue3lh2i38WOHol+cxFdlmadWodpJgL69ek2K4lvIhwgnXEXBnOiOd/5PYI5mGcQNRgTaDVLNC6CAYkErN151GUYQf/sb3KHZt44Z5uUdB8BfH8srm6Edi3AsSzLAFjxRQmi2Rehp7yZhSk+EmRGxEnQrvt7VvaqOOAMN3ESH2lvrVnyG5IXGHej0s4E4iSzVUhSN4hElJOau1KDLLztReI0L9Ud2NOo72+pKebtBhpQ6NPJDte3VOR0YnpIyUFXlq4+tK8jOi4qpJ9HnBLzECLrAHIyr+8/+MHH1e1NW9rDPn4nxi4kKzDXLwblyHOVKhx7l7Gh2tPEZQqOzzVe/LAiqZwnTTbx0FceUIJzDaH8TQMO9LAGXSbltDLT5ZHITN7tycYEuDyz22AYIAclOvjnoH0MZ27xeviApGx/CnHuvy+QRTZ++T7GkabGqugHXO09bkI2DKjod9MF03API2JD3SlAf/2qqhBzlBflgM8knEF1KflDYUfmZnxdKLRB2Rkefw/uQZCrkpYHQuwZGIKHOeqZ8KEaOnTrLBsVQ4eDY5SCMDzTNkk7NGIyHujQmRgc3nqNg1fl/J3+Bt/hH9VteGLQjmX2ThZv2LBpc5Le6j43mzyttmcYWkBwHp797VKbomdJWnqNhBNqyeTx2L+GNeDzKmDX5arBfTEptVxCuv6K5ZHTVAo0iHMLK9GVVfjF3he+dWRftd/+bakCfTVjjS+6h8twNQr2dUCo5jNf70eiMV0HRLeUTcrT7VS2fZ6dbkYk1U7bT9epFicKtGh0i41ciSSa26gHJLnZtfmOwHUTFFI9jFuna7tma9PMqECq/vK4U9gDAM8dBN0kml/Yt1MIA56t8poH294/Cti8nY6eLPqlGhV+ThuXrertsEj6/BUyyWyvr6fi62OmiaksOavxs9AUnD9weJv2FZctNKDzpr6BVdefY99XnFDrxqm9ZJPDxi44VvK11QurfRgBNZs1BhwwuuDdW62evx3RuP7ZD7jjbonA8Oks4fJ27f7fdKaM2Iko5tNMM0LINW0Vqca1qUNssbd+xG3aCmhtmf9aX5+6p/5yyIK4PZki3NfSUX/3zFWtvwqnBN8XOYRdGJqDDbhWPCz3fUddP57qzR7QgzMa++8PrFSw4MenaD568xRYj2wH4v6opsdzNITq9vWAXMqF4VHbx4op8z5DmMKxKk4ztog+R8bp9SU5p0i29usj9boCBSJXmxaYH/BRoIR6z6bo1At0fhc1yj+QggfDnX1cYqqXWQVslS5JTxLmNvp0T/SqSKagyQACgYhJ9fE2jWO/mMlVe+yAJ40SMCIwv5EmfJ2qP0YL/zNEFLUfY1DBAX95mH+qzPAp9mrQQr2u0prEE4iAhJTCllw4BWK+r8yPoUqFXh6YdY3NuBc8jjC6JEGE0iOzdGI9L0zTObWSsGENrG2XW64xXCM4QpGSFjoL6nKNJ0avL8Ps7BuxXkBuiPQt3ow8vre9RjACGAMyMLTd+R9GjE3iJfPMIA0RdRjNyEc9JS74wEAPFxg9RZIHSMeKIM417ImEUcecF0rAfIBepmKPIF16JdeC91SyGSHEDn2kKEgUd/2TpB5AbIEtSkeDaiCamtWJeEEQX2r0cAkYzIFGnoktJJGXnkRb2FR2JMK1FBveJEujlFp7OzUo6xLyzi/vL8nNEa7ggt/cZH8QEiaqAOOm4AACAASURBVPBnjazgumOWGZJ6rvOdsJN8Rj+jSLiTa54mq0ab1QiLwdmypG+NtNZ5oosUvRZVMe99sQ+6TH+mfjphGX5e+heNQFgICW7uRFT8l/8F+eegVBiOJiZZIX6bg/sdQXXz6vA0DATB/Gdxcmch5vozbvKz8mihgmKYGhjtF6IpKzOMhsZ6R6jGCBURQw+Za9BN6XJIrW84YItekGlj3Iy8LSrwWQ4ytvlXoNuHao+koC2ozdaNW/fOjxQ0hagotqNdfO3ZMZ1ejLpGLsizoicq8m2+7w2DEc/yMegODzOhoV7W8a/tckdUzp+zzfSe8DtDFPhLV4zsFuNYCo9v7fzi+eSHR8q4kxW5BEl8+d91zAeiohAiNQwiJTfz/WtefOYZDujhoZl3FE3JlF2cDS0SHfQ0JiRk0AQU9TXZiJdogo5I/ELdaf3EA0XmOGBa6jSkY7zrFR+0VYSsDlbzG+fP63i3oIrrCJEb1eOh8/il0U2SR5FgJVzMcypTWdHwXRyR4qPRi05zdRpbywW7mQh5X6gwIL2BOt04rpX5kCsVnOtr660vW34wxEbBXQgLP9qMlIqEjZJZ7k/ZzN8GWnJ4l21P3sDcs+YaNnV/isXrLVAoYE+wam1uOymSYtyTNh7Uu5MvHZNERZJO+0SF0jqO7VrLAQ3/cd3PREU2s92x12DORr+UsZTzQOjQRRtsDl1eLMx9ev8BdXVoz2mlNL/4mURFnXYCQVxb816tt9shz7wRaw0Spl1Y/nRg1U7qpwNDObyqa2vYW/Xqs0rO7Ra+gzZoXcPtdJ19T0G8TLICHD2QbmawGdd26Z5YWX9cTVi2tis/FfiaL+26fZ6sWDfk70NUNINwuhPrCCWO0fqMMGBShbzv+q20GrNe7MdpeWopaSymdtXIuAH87IHos2XQdzX5yTGf87qnfF7fL+Qwxn2IqVkErAVI3tTmsFHt2tosipq6tbYzweC5zbT3Nz97ASnDIzI9aJLN8/P6OgcrtdA6fNV6K9ONmQYlvet5Hu7XvFLlCPQedT7vy9tXrTpGVPA5xarzdDzmLOl5/gEOY/ky8qbsy1Ox9dqKjiiTLlXqK46N7zWbueZkMrXNjYHSOhdXEmcaDFIe3qdKVMBbXeme5GBG0Flgs8Y18+W3hB/A/8cnS6mktrCeB21GwzoK8Nova9rFdsY0G4NEh37PrVFnykw/pOgSAubpqW9zGumHAKy/eIHt28vj0xPTLCH1FWooIIWWR3AgrQ7SC9H6pW0aRJKVTdXJZDAwhsh3GwONPbzorfYCZT11N2VLn6v/JAQQKcJ50NgLQwibC1EE9h7WEmG9CgD295HBA8QFyILVD97xgDRKtyxErrRN6XFazjvvjDDB8x8evpnD8e+//8FIjmLWswg4U17h+Wwf347fEQGCcU955nfqe/03Cl6LcHhBTQrIPqNegEVYwe6vXyN6Q1EchCAyi4mNsRFbBPZxH8gFpC3DO42ogC1b9Waxi2NJluwGFn0TxdiZHsmIEtMPPnc0qu3duBYRMVZU3SJS7izSBGPJdQKZ9poRliLqxnASFg1nNAv+EzFT5SZIOj6obCtchHTUKsrS17rJqPz/yvHTdIeinHSGdzKx6uDP1E/LpfX54a81AnHCP0RUIPVTwofsCc9pMpLG7RBbxJuCDqix6cEZee0mEIY7kzSfoPVg5pcHhQBMHfK5gpcOaU/iUGkv9v7QS4GgohdO8zblAqdmD3Bt491+7sAUo1d2DAMt9ZhNiGLk4rFrFO4YG+lk4Bi5VItv+/Y5+kJv0wfVXgweI92h+FSBOXrlK1xTDL+liSnhmTS+/DOXvg154cpaIZPY9PEM/r0y4EvNj3IYwaxWUmBYq+pzEVkSYCQXzPRxsoeHJW10Du5HjRVIVS127VaCDOvFQZhh5uk9I68gI0l8Lse5Wh2nPdzYwxKZZxahps++wU+T6jLXEXidCJAIKfBrAW7M66CGIXrrl8avF/Xl4Q8j7ZFcXoGdBgGBIVuppojWh7UOEKsGluZ6CZgXQVBliVhCZb6sTemSTqOleuPEuKR3M4kfCZVQ1fAVDB2YhxYVw+W19BSTFEgcyvgvNhwBEiO5VxXOdFNHVMwTN6Kno7GVAxzFC2sI7Ojxn4usJ41WO2k9LDokPxh440HWdHj6S20eGAfWMm/c8wqkU1IwdGsiZWXb5vUBchuWrhl+RQ7kQh6b7Hh4dX16ALSmnGTB6ilezN0+dvmr++ZmQVb5rGC4Dp2uzwZdWvf2chIKLHcFQI0AoR5HA730bg+7WonFcOuBm9dNo30QJO6Oh27Xhg4Nnj+Xg0Li3lvZnM4ys/6ab+gABhymVj/dulNUncDAOjXdsLXP8rSC3Nuo1yzfcEkXcWC2rsz49uvhwMfFlBedBFh3X17zNxfv267mTy82zRwd6Pkx0G0E+epi6/bOHlDvZmy7gGnj8nA//tR9vH9eBTjz/nRK4vdmjS1HSiAr2vBjIuDFNz2FRBiEEq3V69X3cOLSWWo9qQIdxm+r0qaOFVDEPu3uSFudosLT/s0eucRlkzaD2TGlAHWAfE6ECiyuRYtrA84RNNy3+KNzm/8lwEhEpa7gQXUtB806umZ7tMTf6ry21rIBmupsW88+jSQ0+rrTEd1ZdF7zw2wc0Cxauz05PnjkW/N4Lmp1iuz44e1roiLmxovbGvCP/PgABD2dkGRUcmpjG0vGQVCXeZ2p2Eq3a3xf+v790YBweXyTKKC3vn6qfMcZwjysSZzpM/afHvP43cBgP5/bCvb6FXsTgOufngnUB7DrZ347Y7keUpv4LHVc68TPp6i54MSC7EiD9wHA3zPag2dpFn1Op021kM8lYM/5xX/w8Efbnp9JgjDlECMJQCwIrM0VXD2PRmwFz0MNB1M3JcpE85s4iWcK8DmFrXx/D1Ac40xQGzgD0ivVH83F6wudT0UiyWMenvrvXm9DxFfc46molEpJHiN4xh/f/zAigWdTpkMCNmHRI+9vUXha2LTmTu/49u2bERCUEY7/t29fDRwnudPsjTfvdp+RT0hXhPc+M7rBCo3f3Pr4S3ci/RPTPCkqQPOOz+SILLBde4zAdY2l1VsBmeD/6W/NOa6DHHxB7Q0nBEy23ObDO0Fk6Dr0AcSAEVAWMXEXBLRUv6IjAipzHRL7oNcVAYmD9QLCAWNAUsztDMirryWRCSgYbuvHyTJbqyAakQrLClozSkTnAdow4/7rKy3WtPY+pvTy/mDtINWa68Uu3TJIGYwF1wIjcPAZZAeRToTAHAcRYrKw7e262DrfP4tpH9rpPi/6i0fAl/fB1E8zUUEGcgQuQnViIWPhFIwivTnHTW4wkUoecT5rBjymISvs+GyHLg/OHhFBfCcNEtmxUhjJghMkVjvsHb7SuQFlB9N0PndAYFyGv8MNOntN7OJjTxxfooHgih4blxR+HSEBodsQ4DIxxTirHoFitDUNY5umebAm7oHd81xapa4ISTUFbMYOcjXmk+T5z75WgDDfb/PghI1trNh0AW3PYbVVnnycaexk29beUoMI+FNcOs16Ug2RTJ9F734YwwTYcwaxJjInaV0TNGYnqQ0vexn4HB2KnozP7T1b2Xfjz+WVJAvHygzM3bnbPq2TcH2eekBt5BsIjNXnNfnVjTeDTPg6tXbfesEMeuvYGtbjw61g0fOVItjolvXBbT5UMTLJHzg913SHERUumxVhHchZFbHHdTCMqz6kvslx9E5uDuCSA0/XE4/IRnXd3hAVMYjNrErHXVNrw7T6xRW8do9vGI0quicP78ybybU4DGG3S246WGVtIirSrT6i+2yFRrDBSsZLhxdgsiYu95Gd7byZjO1ho1nTLq84fIVMag87QlSU90MnpbfX6IWUAPTcYP3Nf+u6sAKSWn9L4qfU1rHbO8mci4dWHV/GduhLu7h3JmP71QCjLh7ZgaKnXrLX1LIGBbDy4LN+Q8XTj4GsHVi7fkGH1wcR6xcM49YMRg/4Eeh0rNYLd9baJr2knBr36WKq5bJT/RwRGt/itmHVYwFgdZPadOpo81YzrHVOy2INbThcMTmWO5DVtLUHlvu1nd2TDvkxokLPCx62fXUv+wLW0ga8tsktdIdHWDP1BPdlbTc8LywmNogK3iLMv1OPKvA6Pik7nPagUp3p3HJupaip0eRrAL+nGKE96R7YBSyqBIY8kT/WosVd3shqZlmvQyAo80EuH11IIViN7i0Tupla+2B+URe/QDmxtamJl8dvqyPW8tnp61aahY4uu7gaqG0fdO7q96jZjuXcrJ/OcdjqlT6iwtauA6xW2+BdADjODeWMRYQ70j9lrSa2BGdnAxGLIrFl67X4FLUAcNGNH6CUsWjt3b6nwLtdERv4vRIVeKbZuV6Qlyl2VA+CcsP0O+9MC+RA5DxFVsTZgEsWjk6HH74bwCff7Sk+zcatmSwmW8qjDYPQQUtATEQaHgDbjFxQOqXRyYne2/hRaiqB/Ep1A5CX6aAuRrKwUHSe51PfaP3kGZfgLPppgzwAwkwhRTnTmZYql4Y9CA6CuQSXbU597iyCQXaMeb4jBRZIhHcDgSOawD3R7RkWXUHQX6STIgdEaAiTgZe/geOObURkj0UkeOFpr2Sd4P4XkwESB7fmvS9HTYsUeXgYSK7V8r29o1wjlReIor/97V+RbHBdbsXVvZC7ao8gNxJ+B6GBsf5yj4LXXFOvAPutKDOjcm1urXi3UrmxkDc+R6QL5tmiQnCvpQLjuZhzxJ9K9Fj0iqfPsvH39GFGTDiQH+suCHI5DXHuc9/KupPa263gvK9dzJucYkEiPT49RpSMpc/ywvG4DjU1LCWW0mLLpvNNXc/3pR9TYYSBkxgk7ShTisqojiozvqAaLXq29IqNYdFRkepsUPzVrtJa2UqIkaHQOyAoP1M/rTf5z09/pRFIS4/GHP8zlvLt5fKO8KzX58vby+Pl9fn7pRIVhGRz8/Mlkhu54fm+gbh2SlDWP5+KaQP/35pDxazxYtPxyeQBpJGlcdxZpeVzB3qqcSRwXgrEFIby8MUeymeI1JgN0y6MufMkkZrNfhUyBKNcC8T5V5XVHnL8VW9EtyCXADg1fzG5xxFzrrjuD+cFd/DK1+DlY1QYFm82DxXb7Lg56fAhosU2rJKiSK0174eShy+8INxrBUWWxh8f5cApQjhdZpqDwGKk8nChw4bRIyEbxXwq4Daer6ghXy7lnipLlBdQJ7x+lB9tSjWPfR3juR9ZkD3tcRbT4pivC3yn7Ezr6cihb3GC0ZjJaFyf4n3GDICVShEI4OcJs5L80OOH/t5jbt3YesDdE+7QBXZRtoNzkndWICrBRp8HvzBA7ZgegZFCNGh2hXgOERqSl0Q2qIM0XoMWbrs0HBWPgGaVbd4ZqGEs6noZhn/0qlP7eXYYdfNVhbOZVq1t19iTRzNRgUxDaGutApbTC9s6LAOVUuZ/q+IOdIH7aPxsgI6xk8s0cJWoKAS8+9gMSNnGWWCctNC9W0nSnsdOjmKTxTGrTsxOVTJub5BWupfrYuZw+/396pAvLxicYGe5atGej71rvmsGWv8MouLIMq/t6oCvDQg3gTunRkT22w7SfGSbOfXOsC1GD2u956dN9URUoI06dLbsU9ORM2Mwt/8MUWFtnB5whCg7Nv71wbJdBExubZV85qr34/W1zUk4cMRtGnYayD2bz8s0NuekQOuV+5fv41W8lmqN6SQqD7DDCbRsB5vvEJB1VPpyDQjvzdUOnL68zV7nYK6ICsmQnmXnRAMM09vzmLz4Vb0i4l4VY5uDbCZjWX8fXXebxeBNWjt91V4d3ECKF6zOOTpvjmezQTOv969GZLs5dRfczbMgwqtzagXlUsauz+SWnG0ck5oTSOH81tNhxZK52ATQK0JgJj10XpcnuAHLbwSMSUZMDmAOqj88fI1US5af38kWKw5sufOrIwbXtSsUjzpSxMHt5e3V8YRSVwWfyCMfbQQJ0WMFfDSAV+T4DwdFX1+4n8D5DfPve0SH1RngihnWjZ3DAujPK9AmrVkA9OijPL+pK2cZZ2qhCqhq3RnB8fZqIDvuUpoeqq4iuMX2tc9LMWGLHDcuiWNLoNsLLxcbXkXHeT88+J8Jyvu8mWOUp3tmCiIvGO0pjsxr3tIcgZxhEWm0ncA7ZQ1twd9sB4pEw7MdjqJjiiZ7tkfOqAi9pXjCeCK64ZXyI8yA4+oRpd5/vZNOhW92392XL0akdDJixbRvmGJMgDnGxcY9UpcjioAppiwlFJyNPJWq4QEidFRfwsfMIgFKiqXAKEreZYHzTB1Fggt9xLqDTH5//G5to5rO4tKR/sgjMr59+81ILSucjkgcjyIZdJoT5S7Vo09ApGPyM/Iba24YofKdbWBqrXurFfL164O1CTKA9QOiB3rBonw9mkLGBPVh6j8tB4qIo2cevcAonhemrnJZlL6i/gCJ5noD84xrS2RUHU/tPdYe8/Wlo1nuv8VhoNk7cQvxtssnUXF9C/u84q8fAV9pJyMqpFC5ydVejN6Z9r0ZEtzYaE5PYX1+u2C60dmadzg/UXw1E2AXmDRvni2Q4d4Vcb1AzhgKeq7Tu2BFnLAP1q4JPUly41y2V40TCAmZEukB4dpuOklH0Z4SOqfUR2pXbiJAAdcpkNJQKCOmQlqaG3/3x8ChQFE34v7s+fqY409eaALEuB3J8OC45M6wBDVdzuSpYSmxNspaYOaIMufz1ha/3p0EibqTQFolyKI7Id8xiOOhMw6X2a65b2ZEeOqnlLGySRYwOz5t+m05QD2k0UgeL2K1JteqjE+GaXf630HEtiSFpL3ThGMKLR6Q8iAOL5B8nUnLKZVKQ5q3zEZfNaDrd++XNEbnrua64zNlLNdGtR70AjhMWdILxc2PYEMSzyMRK0OfIpQTcg3YCgij3rOX+alGkdTOpOPoRJaUENRoTCowO0gq36sXIUOeVk7EJNetaCzRn9Cf3GwyrZYdoFyD5HhdJyqy+WV8yx4yDMe1gd/0ZUGol8PaZkCc/F88puH7RDd7pE+Mb22oZKlM5hLak16uJIWeQ6/AFCd/ZuigOWpob5lqXsfBnPXvLCuHF34H6IxDMj5u3aTDr0ydvL5l1htHHrw6JO3e95MQ54LrblKptOLfvFsgSVHDS9E+Mh5nr1lOqTWoEZCTL+hEhlr9J/4sXlR7MNjHO+47nIMRxJq2laHR54eptoojwOG2XWwakL3FuJKWtBnHffwMUTHuFedmaAQ4udeU5bEQKQOkzMGmMBpXB3U7TrxFZwSBFO5Veq4To5PYQGCv10Q4S7nHbL1FgEoAKObRXt2fDjbu6phMZIV7pGNcTRZ8Te+u6gPvqK39aUSF24gC0PUOtbU7iaxGruvCzyQqCNDXtbnVF7Vtub5peOjvvq0LM8YHgf/kOud7MnKi5n0nqEuP4fojm17gPr23mbc/z1VjaiqakR7BAGDXiAR4yhM4xVlKnt9c94rgEdCu1E/MFlABTp2HDFj2GgCR0mUG8UtHREaAqFAdAda/yHMMrolc+5ZWkcCwxm0YlwVRYd97gWX8ymiAle7NJzEdlmM9DuoTk/Dc/w7c40EA928drLanCksJLMrtd98drCboHdMKUWX6WbAAw9Q1chREJMDL5eaOzoMG9t6BcGHKHNb0YN0DCKbqrUJk/vjjd0tPhHnF+P7tb3+zIt4kJCgfTGtEkJ2EFVIY3bnSJ1lk/VbtEKtpwLRSeIbVWDD84/by9QH1QZgWCc8UGaDrVddAc4q2AmBXhMqsD26Q7uqF8kB5fb6AbCMpwXaqzoOW89sbSROsCYD0z09Mj8SIEJ250UYSFeY+6WnBqtxxPJhOmvffO+CPlF8kHFDnYiYq1FZhErgWqa8QoaF2RJ+qveDKhE7OSXwRv+O+bGm/gliifPzx+x+Xb799M1l4+Pr18vj46HNKGTNiBFEYvqkpCodkZlpx223S08W7czPaZaSUorEuFxtTS2flKZ+MqCipQeW0K5nksku5GFJwlTmY5WD194yhfUZUHBm1z2v+4hFIK+BoRAXLlZH5jc3d88hHKoywZRYHkOEwuDiyzQ7icRDzw82AZHnBpglo3AXUK8h0JKJiOkTls0eiYgAzNzl396fZo//CSkt7IGspcNfJ59jW4V4UKnBuRoEzs2JkZWRkHRE9oxp9Y30K35bGSBLbjfzew2f5/QMnzBpLBeR6X4WxwECPm0FJB6FHToBmAFnWf+Xu97oGm+GvXt2TtDR5fa8BQzpvcoOUsSpCTWY22qMInTKgMroKFRdNtsLVL77m0hBLoozPEfjKuRtczfxRHDCGb8qgZAigeVDcTORaeNGvoZVOBGqx2vlAUoHM8JIeMfZhpmIdeF2NjFZR8V6Bo6EkPgADjTpIhuR6xWI+aeiMfeHVOgiJIDSZEHcSgzEL8Hzww00MV873yPj2ufaC5mZAVqDjYO9Ng3sHDuARg8fPPC7D6+NhCr8ddU29N8eIpIVSPw2rMYR5MRvLdeo6zXUlCWfVYyAgJmnm++t3272oetlv2qUm1YXARbgUnTVgsCIq5vvHv9mmafXNt8TXE+QR19W9VGO2R1QslO7QT+RulY7La0fCvB+bccC2hwAdQGIO1kO8XrIbgV1fdjWiYtpvOAuHN0JXEM27I4NkStlah+f91/ajzZt+NlEh/XFk1Lt3xxriOK5G80emeq9pw652RAke6We5pu5IRZG7HJyUm5X6m7f4MlD16WeIilRpPh99Wv8P8DkbRVmIirmDe3bjvLekXiGIpL9LH3bmTkRJtY+rk8KZaZft8BGiwra6XcB8vToSPMQTEgzmRndOzuL909ru2jUTFUppIW/s6gTC82U/mruA+uq2Zs1qr4j1/ScTFXnuqynr2g150xOd4UxqvU/Trj3dsx7EvzdREcfoUn+h2d0KsOy7ZiMHtNDW3ZV1kVsG17pS1xjAr/QufqbU2NazuaXYcdDa0jTB27vUqRjmwdOtqHC1eeX72ZLe8+8R0SBQOuwCN4zlmIkzaRAaIlBivgla4sdSujj5YREMje63wr5fvhhgjfoZKgpMmzedLMMGU5H5eF7uUIzsKpHG6DecB0U6eF5//K1+12YZgF5SeulZNhalWDGBfYL8j49PRiJUudXvdj9f7n1xcPiWdUHIgbhEGNmgGoWl3p+TohYcYCQAoxHMk93HH33Rc5RCCv22tFoG0F+MoPj6lYC2yYan38EYMzpCkRVZ24JEEgt6G1Hhci3SAi23elyqpeEEhd4p50FFe9icIhIFURROeKAt8qqfReTp5cnAd6WkMkIBBAWiGyyNE8+Tz09PbAP2CXP6S/Ct1m8KPMPBdOJMHH+NJea1Fk7PdYSxYESFSJ6arqzbW+Jax7iECUWK4FlNKJWi45OWJ8zmmTVh0LXEPZJAAvkBPWARKiW1kkXKvHDOlfrJSBRvD0VJNVm46u3/fVlpeyIZRTljLdkkFJUKTLU3bFx8/VcsQQSVjcntrUV5VN1G2yE041oN108DP/hM/XR9sD6v+AVGwKX7YETF//nveOwxiMdCJR3kKLvpCNh73PVw4GkOIXrwfOCK/bRCRZkHnl46aeTpqs7wzUiF4kVdIiew4GMTmY1rb9sYUWEqmZvYlVN1a/DDsLqlV9T2mgoS+e/apP1wIwVo9R0QohmhYyr6g7DJMSyRwjd7EFZipB5xAwqnMj4F0EQMwiTvN2yrM8vogxWZCsPRWyhjTpq4OM1XidC4KX+ibUroTtNvQXWO8BcOZh0NExuQroy55mYoL488KLP9NKpcQsIwzQVTia/wEhk2lUpUJDlYN0XO5LYY+jjgbDDrdnAWcQ+JChIow48TFXN/dM3Wq8znSwWqFt6ZdY3YeFbjeKEN43DrBdU99jdCK0EbBOBtkQhNREV7QNa6zTXm59rpyJQL++19TnuT341AiYe1Il/o5hQpcBivqUqD0RRW3ScMcdO2OTryJtJhRAb9ZIiE8K3GtYzTTB6tN6WpDbrIxnVQ/uX2uo5CcdJY9TBiebxYWHnxfhvW9a6u0aYxia7rNoNuKlFheVip9uzQopR6vodIy+WWk+2ONVZe5aZpDkFM5XYjOERUTEU4fUUtluW8VivIkXu6+xjl/dGdqkS1h3dEBQGwlS4hMIYxXREVTKWQfbiyOS4ET7I5i9kPuaQ3uuAoUUE9y66d2wcbJF79VpoypTsQcNkgUC1RYcO8GOtdEHRn8KevIhVfbbdU3Nl31A3BVEmsqHjrealZa7DdT68Zbh945Ebnx+HwAw9bjKuJ4CzLMg8HHZVSuqBFR90QqqPdMK82vheB+sy0l9c2cZ31WQJq8e0xuiv3XzaTbZm9wKe9gobI6Hj1oTRF22gG2SbxxmGrHCMqXKW0ET3748RNzd6nKPeSJvXqpPkFlagYrJJmUgVsvSIti+fX55GCnrsWpVuA03m513alPak9ve5j2x4YsZSD5qeSLOZrd2jNuW0xPTlub89lzcAZKFvJHPvdaxPwxbPWdIGcnL0imj/PsOpSulTUPXRnx6nRrcNWk0/iavBh08EkRiHbvFKHxI5VgHrsXgcecg2y/TpHdGOttu1qntJHPzqwBoEV4f3C9CpOVrJ789pOkNui+D2FUs2Lz54Vm97Odkj1w+LQ+Or+HgW7meZI4CLuqFFE6RRDxzm2i4DpbM+Y57+D6Hi7eZ47uLkUQY+EV+oaRFbovgA/AWgHsJrn93n8DXz1mgA4P2nukSIHwDh+FAkSuiXOdimPICRQkNjaYemBksjBvKgY+dPTs6WRYlok2Z6+PLTkKWwbouLt/eVyd891jxRaCXinwA9k3/vbBaA9QHQjDV4RZcH0Q7iOKalY1wTg/QtSIFm0N9eyYQnCI7woNcYHdRws2sHrLSrKQyA0i0e/WjFreOqLaGCX8F7KKYsyq0j5q6XyQr9UdNwKX3uBcrwPq0XpvgAAIABJREFUY4e6JCjsjfmpXvqDnPg5R+m2QAoZKeMZKoys88LzjI4A4ebphtwBWbUlULdBco4N1epv3N16NAgBeK1tESsiDa3WhkdRvL9xrkHuYPxZTPuVqaiU2tWuyL2MtUzuI0qJY8dIlRGGoWOorXbfc5BykOuM0S06U7I+B6NrkApL9WdIYPHMqhRyGAO8X9eydWMKQ6XWqiQPoRiRYjzLo6+KwhEJIx2mMVAdC8mw2jPrAJr4SjGXqZ421y2PAUlI2rh81qhYqtjPD3+pEUhj8EhExX/791io6Y2tw3rNsVe7Z6RAGJNurQTiO8c91HoJVwYpLCkWYtTP6PV68ogbzxlDwDEuNf1QbZkMN3528n3Vg0Z1MKJfelZntimEsLRmImw2I9idIAertE6WDNybMCjCi9+aNfbX5GLjwTUaIhWUn4crCa4CcE3A3RLHmzo6ez53mXqrwTZQYOaN430rYzMAQzHftsUbuBxroExd3pMHc+Yxm2Vl72CO5pQ15/01A3NRj6SXxexlOvQQuhjkuDRFHgOr1YjDKaVAN9B4iHnczF3Kso/GVU24EDN/ZyUkFmukzsFcX6a0mceY+WckO4b+FYNqBPhpwsxrogKtMi7syqagIFsismJeYzwMV22n31sZL7lyU0fu6Koil6OIzu++OnV5IIZMaJvZ+T3I3miodIcfdKfPjeSo8heDXTcESRpk/M08h6ThUkRqCN+4LrdRaNf6/U7vpAWwP+52+fZOw49yl+8dUrRRqEJsKD6lmLt9TS+0+WckNnf2rk19ku21Fjbuak3PpSfhKHUpr1UXTM9rmiKCK/pxfrsdx2kaEHZz9dDGE7jUP5nHtgVbjmxgw8PWGsouadu6kr/p+iFUqGntFYIkTZUyZh5qT9wuQ+9rlF3t3pyaI6VlPbntuLp868BcuKQG+J3Ddsv6apb4R8Vt9bjajx957gw66bnzM00leHagaxqsfi9iowLY8uSrBSE7+Y89L4jg7dtb4FKK2u1kAgGnqUGqxFaW1xJVna2OjpfAhwDKHMSsz6rzAuAi1bfvU/6BAFa+uwxE05ihe9ElAm6rH+ZpT52gtdwBztECOZZoR9lRHf28Mjd2bJH6vQpv+T3JJlFOkgG5nCmlMK3YqlNyKNxSWAyHXRO2BFOfGBgmj4YYwOxsr9/nlc33Ctyy9DU3twZ04/FwEqKALgiM+BD7tylUc2Ch44XfFJHb/LsZwuXn+eLUuj4US1u2Xk8SQGl4WCx2qed6hb28Ht7HAGJJAli8fQKd0xp2dXBB2qRwfDEgFgDkk53ZmXaIpJn0AKfVGyZwwus0zBMhazGoHpN/rslco6s15t7cKGjtU2U1FrzXLo0xj0xDpELUKt7LdmdRav4uPTgMYFERAmxrqzRfhuF6cWB+RmAePyASANwaqG5pujvbg+cjRXsom0PcB2DYoyiY4pXPA9grIgnOct//YOodjBCiQszZ0lLufLFxQsqfu1sRCi9gSy7394h2YBQArrN2OLmQ45GrwPYqA6nSUxbndJ6dQXCpbiNqWNxfXt9fI3c/CBE68jG9FybIsj+gbsnTs8k8iJxvX7960WqQFyBEvti1IDNEHqcDIuUH8glSQv02B1MH8ZFGCn1jKjPqB6V+oiygngSLfcO7HuP69Px8+frwYDMGQgL9oAOoO7y5cxt0G+ou4EKsM/QP77u74xyAzEGaJFyH1Ff//f/579YfPFPkCeYOc+CeOja0FgXw/maFqTFnjJoBwfHmaaBIemEcLDrF17f2TM2ddL10DQgdOK9CX4K0eHmm8ynGHO3GuGAcrQ/3d6zl+fZ+ATZhRAVIFRBuT5RrEkM8qIBMe3p8JDlk43zLNFXPz5cnmwOmx+IcgjwiMcnt2BdcbuA5HtpW5cgEYvOOawvvRBvwOwp543lWZF57Dubaa0egXgZTgFEOOvhuVqTzXi6dIYLsBSSXp1q37z6JiuVe9PnhLzUC2rDdzHEvi66Y9n/7D8WNqwJDy0MzOpopS4bDawvryyDbGaSyA9tGAuNtoFcL0Hx2rG04ClFBJqY1+Af8Z7AMrh8/6wFmPH5tjpmLXnATnQ3TWfEPNx4iKuodbj0PxdWU0kjKulxvKY36aIQBwI4uZl9zPEr/Z2CnxxeiIaMs8HCz/BmYh0U7BkJhDOsenniDTS6Lp8W73D7S32P/5jbVv7ftJfjJn0Fuwltp1cftO2TPar+NfJ4LMF/v2jvkR6sKwZYc4vj+oQ91Tq4vlSpk01Q2a2W20osHhq9we87aFC+F8SoJ429ODxI+KX/qaZNfjQeTBAZ2iQqba62jWS7WcnKMjKtD1wz6zyQqTs1rnZUQdM7RTOpU9mfoUtUb9WDCz0H25eGrW3/j/jNT6WtFMurMlPNuTU/vbg7zHViWoGFohKHu04Yk+VGigoPXkmRmObxzbO0M4IzFHlExgiplPPZkZsaArk/G+ooOPIHn2slnds3tgayzi6IBC1p7a9p0Bj3b7KtdepgjJ6O5HYWoINjh9mLX3u4dJwmdaj+Fnal3d3N68h0nRWP38p8mykfmqNORBztkNkNxLpJX5SGiopwRujWxsi8q2C875B+BqKhtlRdqS3pY3bG0IeoSScCmWhCzvaEJFAjrfzd27bBLyW5kg9kKAKVTTv/cYSgDZuGUAretc5YX2N6KGOtErX56nXlOKyMdZgW8qugu30slFV/R25tpYgKXHtbAgsOIqejbyqM1gS55y+M97SbVpu2SFc871b9zo9RFA/bpqwR2BxnsaXuZrpf57eefs+oJxA3BVJIPlkffC10PZ+Rqaqv2SaRBvjWwEYCggb0lVYuKRq/bOu+dPr4c5eMyi8eY9zgbqZQ447khH4ercI2lPwX588r0SLi3RgzUAuHdOVuOo6t5qJ7vtNlqRALeecdxu2dNie4dkFnVnaj1OQC+so1UJvyHuiVqVygPv0XI8x0A/fHz7es3axMICnncs+YD60hgTJ5eWLQaMsdi2oxsMvtzmKIRGRn1KfEdpmECjsKZArFl2QUsHdW7gcl4KEF4pE4SWcHCypamyUkLttP7azURkqSoeBL6+fL2bOsF0RaM1EFBZ9a+YEF1yC0jOWxMAbqX+hZIR4S2GvHlpJKlL/JxsPorpVA1328a3mSL51KmMLJaDF4knEQF+sR2WHqu799J0FjUByNgQPSg/fjNSF0jfNRGgeqKqOP8SKZUfD72FU+dpPWVc8g1gL5iXIzY9fTyjOjA3x55hOgmT5FG2QAhwXHE+7SG6l4VUUdKF4VnuyBY3Sj0DWC+pXmjTGdtlJUqqMQlx9oIUidzbT49qgq1QliLhDLL/nmhdruLJBrkwoiKO1SQJyG3/5P7uPYFPBvzY3PlJI2ILls7n0TFlTH9/PoXGQFX6AdTP/1f/2E8tMQhpjuIIjw3ovgmIGk5AjMgMl3kj6gA0tsM4voB9KyRFG9yj1QejBwoazyTBqaAFIc/Zg1I1AOfqxU3gwRI5H3zYW0cCXnC81Mbfo1zI1lnDVk+eATGx4PJ3EeYHR6Wt2pDRCnkOEUpj3hUyTEZXkTlYb7hbh8/FU2sotYRFfNj60PjPfmgOPDUdtnXTlTowOfv0ya0IWDsnnVh85TBsYcV5Od8r+VruGsz4fQk4JqVMcnn9BEVbSaCAeSvh5dhHZUGqQ8D+HugG7PcSy7HlEm6yju989xKZHFO54vr3yt9VI3g2rp6evoZREUVYim+tX48S8a1AIO0V1mP2cNzk9XhgP1TyjexliZv2OHzuoClTeUJ5nqxzC2jktIbU3f7kUo9H8TtTI8lFZuIimEdHn/iLlFRh8r1ET3HUp5JGIg8npWB+0q3+nTSsAeICstxG+zc7Cyw3Su4WoaONDuXfzwtu/39sdeRvafvntJYfPchA2P9jvZRJ3PMrwGVYTNc6LsGLLtGLlRSs06RgXG+z9jm8oFCBydJhM7PfnebPPmOfeE8921djcc1wvYdH7LpzjXV7YVxTneJ9gLrjaD2WjrretSa1phEKpWaq/xk+ymCf/5IKdIti7nS61z5rTfNDqIid6JsK9ubOm6v09m36ObemivjcVT2iOUnUWGtoRF5ajY4D40z06kn9RfbK5YpdBuwmZ3zVBr0AAfwRo/mtKyqg0Db9V6RW4NZPF1pk9PTf7myD9TKqyuqtQGboSLxtLUL8vJxbgX22rE4wH8CYOalfeKnGyakcQJ4Zrn1AZAWr3I65hW8wh8Sdpe3SZ77BsKpXqPW0kciuzqawpwzFj9GVOSaJoCs1E/r9YK0OwAkCSyCJEPb8beD6ZGSyQtzAxxevX0nHaXmz6LwzfkSESdZ+BgtBuBtqYWM/FnPqXmvIwJAResXznNVX0hXyCMff+N3FEpGNExt15f7B+u/pSUqhcepB0mdWJbiSNvEtMVVv1ewO50lCjHn3vBGRno/0CYrAu3EAGs5cBLN69zTeikNlMBf6gqSPJxjkhlJKrkc+HmbmoaZJ6ALcA8KaYOosLoDNpYk2uzdFhHkILUIBiMiUHiD69AIBNzzSi99PNdSGjlRx/tVuJntQdSRnQycrBHxgcmgdz+vj/d4iuWoZSIHMos4yH3AyByXB40fSS2S4CZXXlvF0j75Wk8iKTUaVjvWBX5YF8WdTmMtMYqDssF0WkpXhnFBdIQR757azCJBSiSMjY+9H9EWWV/E5NrrSDCtPDKq8LxEe2Rc9do+RP6JGIo+RSpEjg2JKaa0otz62VVnW2sTr1XhciMOD9W9rba+9mubkSA8bMzukLqOY/sZUSFd/fnvLzwCZeOn5qNBCiWKnHWvL5e31+fL28vj5fX5+8WICu+NoCGCnM2PhalmwVduN8UNZHPbKi3OeNEIbhTjpR6cB0N1C5JsW5vXRP+cqJDiXfVw8OQbRuGIAV+vmWIqSl/Wh6wkKog1+bP2DmTXgIe5g6b/537Uv1fg03wI6e7n5xGm7Zdp08kD0Hj/EhAX/DgDWa3v1tTRCXCZ51RbSQ6tj32U81BqFXWCByVuXNwk8hUeYbRcLlkEbf7aQhrLTwdiDuDdxoouRAWDpcOLgGvYb4ghn3Mfxkh4Wg9P61bknkb5AXVXpnXPa30XS1p8CSPQeoYBD2XTEzFWjHqlg+KzsXB26q68L5fedHD/oYiKaRCHVGTbNXVtyLfy0umn+qS9tX59jj9EVBQiQm+gF6J2m3wvW1rmoZISc15y45xZMG748fWZC3TSN9cGdhoG9Hn/ltWYru/o1kVSLXURFU9I1FDRWNglq9RPRVfVfevdDx5NvZrs7rh3sddKi+DzMgjAlf3wyHbZ6L8OhNwlelbiu4dqn9072+Wx7ujPIypsV503uGnRzG04SVT0T0/bbi6CeYRYr8/tHI3b54wHyDqe/S2N0P20ue51ZKdlr2vVefCbPjQC9RFuxlJGFfJpJWFzu0VkcB923dS0aSAjyoNsRv0eeY7+7NRPp8d75wa2lTZA2kEEGpfqZrLpNDwJSPA5Aoa7V1dgzubmyJ516KJJbZyJqJhJaH+UpV+MnObTVtzJ7NlJMrDW10V5ZgXD6iOLeREFgQFw3QPosiKw/PkxooLPiBzkquNWgKppNNpC6Nv9zs9SJ8fpPFHBAsEEd5N/JtjYKex1o7o9m97MBKLTY5yA/ThnBP4NrvACtFon8kS2UXFPaAPqHFTulsdZMjNSCk1dNC0QGH8WTKbcL/S1Qx4EjulJbrUakcIGnuIuw0o/vYefpLPKLE2ZV19EBYDbIU8/UhKpfsTL6+UWtSAWP1lkOddFpCCeIikMSPeIaKT+gewAQEbUBMFxAupIv8PUOpfL77//fvmf/vW/NqIAn+k8Z57gbmdmfVTW/cgUyJzdWPZuj9tRMOoOKbUWr7N6DRYJ4hEsHlHBSAO0gUA2BdP/0bUgN7zwtsYFTazrId/rBMsbAXXuESye/Mfv3y2aAZ9ZrQyPIjJCBp736LmnAbNrjFQBuXHHKJCbW0uNhHG06Iq7rL+B9zNKg6mMOFaMaLG91+aIWIwRSL99M72H2hqI+lAheUYxkGARcaB3g/TCOsT9FqVhqe18L7RC1S/WDxULf3hgEXjKwFjzQfYrzzkk7fBj5NANU2SJYNHasHRKz890uLSoD4/G8sgW1iEhQcBUUc9eDwTPFInC/Rsyh/aHzveILeolOlcZfTEoktRHuk77Te55JEMgJxhbOTCgXVHHw1JBUdfN+2S/ZW+tSbQTMoS2YqwteqboEpsvjxb6JCpObpyfl/8VI+BCfjSi4j8mIEJDgH93oIAxgU5U6NBy/bDRoxYzSWELuh7Mg1yoBWzn561MlUQVpRBqnw6DRmHVNkV95xAMV362X/h38d54VicXGZo8F6X6YUnaYqGDt+6wa8fLlJ998XYBgr7bi3CwTXPI9Y0X9wDpLlFRXlvn68i5rRIyNwPKoYdKnrJ9FDVP/hzAXr45D0a1T51shwW0RDrniIq1AZnPXm9qdVRYkIweR/S6juNOJW5WdaDdYHuPqJARML2C1Kaxd8Abrwe79c5xPM0jqxIVGigJwWb4le+3jmi5yBtQzxcdCFa9I2TU1iUsfRlGSLtIV4C6y5BOX3HvsUPqeaKCz00SptfJXTfauWuRQ3/nMBXTflO+q/T4xjN/gQSuiYqy7jRpVY8cUh55Q0dUZPtWuu3cSzZEhY9nHAwGUovG/hK8jqZUef8oUQFhqWDCtYiKQVm7rLksXwHRZlk+S1S08loF/ugG2rW1BbvX66jvQy8b3TfdSiXA4cp70B8LfbPjK70E2VNRpH+do1nnpNsbdpaoqMRadnRnFncYxf8BiIpd0O2sKidjQDttmud+C+OsHyEqhq25yEztwz8CURH7epGfvbPRTSEqqhpJciYjKpSSaSWaWxWUYN01fjDuzUPPekqLJ7rsGGvn6cVNMGj108nsR14Rlah0vL2mE2IPJbFEj26AOXkaqe3bqNGwM/u+EZiU17WfDz9MVOQi1hw3Wbt2lihB5PHHLZWNnclpo0+7O16VlEv9+b8Tp26c4JKFQrf35iGOd7LQtSP/xaCOlE7mec7MDZb2BoV+AbSrULN7VQuIvqaz5u87+euICtMDqH3gdQFE6pBsWSnf98vNHdPYKK2Spa0BaAygGHUGvA/0aNeZefusPaICOgQe5CoUTYDeiaHbm8vD/YOB39Jj3fGMc0NSQdEMkGtLZxMRID6KPngC3AGOqwg009sI0FYB8S9WkBsRBUZcXJjmx3Ckt7fLw9cHA+QNqPb6EQShWUug6pYEihNkkRpgAWn55RJkJhDP8UDqMRAIkmv8C3BbRaJRz0Nrx9Y0QH6XUdR2ECGg5ZXLzNf/LTzrCa5DTlF7AYCyvcdqSDDlFHok8g7/WtFl9/K3wtpfUA/iloSFpT96ZwF0B9Rt3xQp6jUb1F6Tt7c3i+hQijSMu5Edb2+Xp0eC+kYQWfFu1qExj/x4JolCi065u7VnYd0aQSXZ8mgKzQ9EGUsTgLzW6FZ9gnDgHQGyQxa8ZgkJX/4XbbEC66hlQtvOiADXH0yXlXU2QKhYJJiN/xiRozoqaBPWi1J/sY18J35Sd+Z+m+QCZdHWhREsjKTQD+eOkUt4P4gL1anA3sVUUSzkbaTXUENn0lA1k0o502UaLEa8MQUWbTjTKZ6C8JOoaHeEzy9+nRGQJedAuTOsbUTFf8yCdlLi+0RFepAHULcLRDggd22AigUub/MRDDp7GtsypUeIiqGZwyvXRMVmrIrhNXxXn9VYSiSAuD/rILd7QL02pvP3k7FqLHKUYljNEwgrb9CsS92yHw1aec3Ui+dx+9g8xhNFJiz6HgdCfecyRaJCFha+3IKLOW1OcE39TuPUfBf4hg7t5pd+yVr+Kxm3EodhlP4/9t6tV9MjSxOKfd6ZTjsz7bTr1F12zVAHV82I7q7p6Z4ZrrnjAiE0TM90w81oNAgEQvwBbrrgN3DFFeICJITEBQgJIdEDNH2YaYY+VNlpu8suO+082c59PqBnPeuJWBFvxPu933a67Gpyq1y59/e9bxxWrFixYj3roEtXx7NWl6V0SYXVjtN8eeJBvPTScWHe13FaHHueZmOpHtaomOHLzwpUSCbkfREIRc+IXsbk8BC808PhbxRy+TX9vLmIXDWiQp7/k8kr2qx3QRkQsTFArF7b6QWYc15/H35moKIywDdXPI/cobSpFpWEqKxf/oylQerLp6kBV1t2BDj36Z3BkHbymVlqOs4ZkkaFhqdnjrepOVvqwnCwbOKL3iXZzw/fx6XdGaAsCtb8u/ISS2F3Gq+KqIjL1hj3RiKhx79fGFAxp8c8NaBiLBy73Xux+N5bZQ8v5cGRMak9zmplxW3a2XCwAncabKSB0jOga+GLcmmkHFjbzNmJIvUhXqWtkVgOn68vWWcOzDzUGfqt0SH1A/4fjR58WZ+NRlKJ3yWAVXB2MiNHQ+tfBKAi61YCaKIXfodQAiqiEat+THncZfSJukj9ZE2uuParFrvZL3OsFXQJW1LPub2aG9sn1tuT695pzI7kYx3TpaE0vO39PRimlBYjaheVDj6cwnhu5A8aHi2ZTM6tP9qr86JxpJcuXY+pJzPe9HuINdLwjqsV5uWeawzQwLxar2z5tT9nyBczIjo4Yf1YrnkWW479iC/kmUxDv9cOCKmWVNAZI7Ai6UMHqf6YhrEi3dRZTjeljPaUTbbuXjC7tz4wysr4asWuLUrA60Z4gWsYVg0MgOHSDI7rHZ1KO4bpy5tehnmMbW9/n17p7n2eC73HbmD49XFkIzzGCTDB7sCFhsrJj2HCiG8G9Wyc37QxsIh4iRpDWikYcFFLATYogBb4OTv1+gibBBHwY+mxsuE1Fht2mSYgIshjO7vccZZ9l+LkVqMDtVG8+DEKQwOUwRjgiY/Ni7E9OTgwAz6esznmOZT0OihuzfoX9SXQdKMt8PiJFauGAZ0pgEhkM2yfCXjx4uohush42OoWEODJxuyzMxunwAGkTLLbuNc6YZYUAHrbudaGAXfnFxZNYfT0sx1/m8HfCpYzqoyprvAM0y1VTgQepcF0bR79gHRKMPI7sGI03d41g7xAJXwmWVLC1gqzUW1gBIf6xh5BxAjALtBJe0XRJJDRoI+BV1bXIo6ZabX0o/2o9EqstaMIC0bZgCYCnQRc5z3jdqL+GWOaEyO+3CEhRrOUCArup8PDQ+Mtyid+Bjmoz+bse73zMdpmad9R/RMBdEr7tfEs9dPSA/PZc18kBSQhFwIVk9RPjQG2UQOK17XPUadr3N124NbGwcUU6TrGyYA/Osl5XNXpRMqz5ZLVMYC1AxvppY7mFiHCByMSzVnr4lfC37IyFmxNXXoMQsqX0K6n8Nl4osGo0xCNEBpYS18Vq+WLdRSKHZtigtwylf9I8ZA6KPBFplOb0iWMkemLvI8cojd2+ioG57D2ukSENCZsk+F+pf04F0SS9KiuOctLKaQjmhg9nA8yheoGR0ZfA7fUdfB4rBOJ6QHlkwTJYxoofC/lo2bouQtIN6JiDqiowJ+WPwJ7tHlWY8RNNF4biFDz1GViREVtux7ULQjG7loChbWogAo9NTIEtMKg8KI8Ugvjz+Rtz3uiYargKZ8VEUs3Sw+rwgaRn8uYllwmW9qpzWzkHIjUHvej597j43GsaLwB+sj5g3cq0R3/6K/RRIzbB+PxjOYw2Xcuw+J6uXBMAAsZhbCe4SbSOvJ/ATYcQPQpqDZHtUZKD2W3gapFV7DpxZN5ysFWykzSvb4oN+CG06+IuYaWk9pHpa91gYeeHB+dgdGY2D5zpVVY11rQ3xEzPDC3JxYauPJjq6I8PztFKrXOh16Ai9GqTD8fgXQylE9G2iPFFYGFSXTqFdvhPu+s30ye9MneVrqd5aSzJ4e8vIb8zl3KktHMRbpHpdP6pThrdFnfX2UfDOdhhz7tsNfdq61MiRf5NUk7fLyVLXOyhovUM4H2HUXIgnOzBoViOgq/bwzk0wgcGbK6DP+1mkZaVMNad2Wi3F8vfdDoDsNUM3RAiUZqGpjISXmPE9Vo9KeQklbDy9dk/jKi0xJQpbpHDHar9+K9i/vL+mJZVQhYQ1TKkJZBaWDz9DZBJll+/UsYIVlHBb1Y+YIMGvaExfSeumrO7fk897ytxmRf1PnZR/sqGuREAxj+ULwWXuFM4TMWgHy/cxYx0cv07qd6Eu7BbUV+3Tu7YHq1Ls5tnKVjTqGVNp2u5SuP5ik1AJRex+jnemVfGHm9xvyMG0wdWIH3vRUpvrhM165dswgFM2R6weSy/gR2jDfc6AwjMY3k2kuMEmKh32kdI2O34H0ucAKfg1b4Uh7sMuRaRLx57G/YM/So9/up1XaoF0lLCo/14+MjAwAMhNj01EZuJxGgYMW5BWTJ/uKENEN/LpqN/lGnhmAKPeMJpOX0Z16EOa634/LlOb+Pqh3WlGB7GAeN0awJgbnv7AgEYcSLzdc88j1qwqIISBur5+GRC1WUhxvHATyp9gULfiMyBDVGCBqhXyv4jNoUSEHkXvzaK6zhgLFhzqybQsCrSCisqdWBsNoi9No3UMRBpHIP9HRVALUsAod0VdQMo4WY4knF1EUrAR6aq4HJGLvVc+E6g46oeYIfASoAvJjWi5yYP7e+WKRb47DIljPKCYApraxgRMJWevLkiaXHsn6dNxSdBGAHP4yAZCotpBAUDbi3NkONCkZUsG2vUeN7Tp+pj5HiIaBYtUDi/sW73fuRRVX43v4b//Z/cfVT+2lpT8/aeUaBWQpkDYzepgYBjmtU/NO/ycaq416SORrLvM8KqKiUhCZsuPpuTS/W7i1m2Y2sPBWf77y7rLlMaeTSUxhmBCsg6Ho/Vcjmor5oLLrKTyuA8/jcuK82u8bxnApn2r8h7ZN6JRpjj75e7NUPPRuXs2CwvjeAR5hxbNKN2+sAFVlhDIU/TZmxSAO/6OE3KXzZSOcpk3h7GmOfAAAgAElEQVT0JRoC2x/Rxy9GtmmCp3P3pqNczjVgZLrtaKmj0mvbRtEbvaOHjfCVMK5815S3UasIaj8WlcPamfBfM8h1IyrKfYzjzMBGAXo0aiosAioITOC7fMkJQ+FqljlFsIkeD41Mg2IrY0knoqLzxtC7aSosC5/0jHrh24ahfG9o3RyUMs+jKwEVfYYa212n4M+c7OkCZd74WGqtkGdXACqm0RbtvvA90U6mknPLpWw17zydkrO8UhozUEFuX/rTv2zHGhU0Ooj3VLyvat+ACqtKOOWzBrSkXJbskAwgUMGx+CW7qmvRA0Ci7L7a2dWjUVTMV9HwiwYqBPgVss/TYZVhZTrfWCfEv83yvrfW4r0e/y3nyVV0X9eLdWQIXBsXKgfe6iFqy8i7Wm9cFaiYMYqNLJ1FFysgfOWMsHgW/QdnA+Picjdnca81GQlYtNY97N0rFM9X3KY7wmccf16SNdvpXdYxvmnqmzUbvsLjeSwDmT/P4/N7sgU0hoD6gKdXARWzZ34e2lXlxlXfK1GuGJ8MT/hdXrEWvSBQwgyhJZrYgI2W6L25hOH1HYFkoLoCUzSvmGk834sMWTFgS8Z0jDdjgOEO0OtZOfyZPkg2bhr/cWOzQrG58HSdy79tr9aka7qPZr0WUOFG2QmYMVMkOvYb36NRGUCFp69xY6CMne14lV6td6ZWnOmEB92yAdJAMRob56I2ZCBnH0XIIvWTfSf7v0dkFHtB0O9WaosR0Cr6GfjcxpxrDhEsUD2FzNPOTwB4LI2Q38VAz4sz3vGNzu4oZrwIUMBqKeSkawS8bJolf7CZb7NVn1l6FHlRaBLvmTwHrW278/WdAmFgR5qs4+MTM1hbBITiiB2Es/HY7zQM21hRy9SXQUkRaDgmiGA8dMroAoEmcUqci+7/Qe+2mgo0bAsEsggVbxMprERbpG86D9FpuNMx7Rm94AVMiXbUYVknQoXHDbT0NcB4rBC2F7G2gvSWlosROjy3CQApAgL9Xbv2nPULsMFSX3l6JwJRSEPE1FRavxhZQcCBxoXpfbrYHWxc3i6ibFAjRXIafQtsybLa7xgE0QhkoAcVmxdrYb05BjrtGQiDwuiWMozrSGBiJ9efwAnw5OBTAzIBxCj90v7+tbz+AhwEJmAMx0fHFn0kMMfuQcHGoHGy/gvrZsiJAO1gDBgv054517tMEa17snQiE/0hARlKo6a/ufPHPwasIr3YM6Disx/Yz1r4vCmwPlAxuYC4gMojHYEOI6CiMWBNojBWkGBy+fKLeRlnfUGvjZZqPBrilhtRhoYEKyLOI97/R9VkwU17Nt96GG4/bU3HU93fmXjy+DTLxUkn9hzBRRv829JJKEMUvlMDlw56EqRcFkWbrEhlQ3QZj7XWnIT5kJickN7BYDo6WHPuZRV1ynWz4vx6Rh7Ri/n+ajRh+q7NLypFk3F5vRcRJnx/Ocs3JSVD2YPB0B8/DEBFayyLgFqlRM8ZXKo5RN7oE117r8vjkWSuq1ZLmiMrmDKMnO58GIGK0E6MxClbR4vgSnvkZJtrSG+XebwzuIHDbGdZu8QoSkr8WupFVNbxvafQ0wXBL9qm5AegYgRCTuVOX8YN2Szs9TpSarTOcaPWhBpL1/43FSVcMyVf4JIxfSd/0gVGWrq6fDIh3el/rag1KqQu/YJ4DAUVLVDB/7YHFbmw3EizLlCBkHzuu4FM6hygBPycytoTvi9o7Qhc4CHaU7V4Tn7OnTGf33dPFai4giG6twazp22mfftU3/uTXo0tL69ah+W89/mtTNvyet7VGaDvDLB/wVsw52C1td2zQHerj8MZPXJkKDaxWdIsSReaaWmtJXmaQEXWrqJM7kWAFIvqWmOde3jB6lWvj4CK5pSqUlo8tcE2DT1toKJmpZoyTw2oGBKjrVOxemVGBpf16a1d4TctJ4TlS4cF1MCJUpy5GIkdqFDNCDfgt1qY/s70beTBrFLXk0P9F7o8R6OkuLMuyJxrL/j3rDHHVDi9Hxb5DZ618iJHmsCQdsdSCvnZbu1M0leaxtUE0ORb7mD56ggMrBjBwSmf8FM5OGhNY7N93qr4v/H+EZhKT3HWOlB6lcmJOpTJsd8iiSHWWo9l0BoGVxl5e0Shob/Y78GXW/L+1xe+/rY+9nt9Akijm7YvvYD6ngy5qnNghZrPmB8fBuyjwyNPxcOW6pmyVosZwFGjYGuboIF9xvot5gXvg2DtDHqM8xiT/lhG2QKp+EYe+krDhGcYoREc0byA8sj0CqM3U0ZxvJZSaBNRC4ryIP0skuqSwIf9HVL/ks5y9KA3POsKeNokc2CobqQhmmSaAllRJ3glplBSBIEVN7a6CwQctF6402F8Kn4tlmDxbHr6W8FnS/VUABUCXaztQP5AlMRWrp0BAIQ86ynFkGZrl6m1APBce+56Ojk5tnVV3zDgay21rlwbRnRlOgb2bLZgWHzyEWpZCHiIfCJwxQztqk1h0Rteb8KBZwN+DEziWhiYA/AF9RwuBPBg3mcZkAH9T08YUaU7ANrB8ygYLp7Ddygoz01X6oNoP6NPtAUZfHR0bHVFFAljN3EDnJhSDPKGaew8ZZvztIpncxwkT7F9YQ29Hs9EQPVFrABIi5CzYudc557tw/oLa/UMqBgcW88+/rJRwHfK0mLaHlFRp01qPCuCgWgcUVHoUB/Bbihcg0y9FNtjo3F7HPesjR3j19AoMbhCCiFdOI9Qizm8IaNlrxEvUt7/qt9rR9+yg7o6WVxwdnP382gvgrWZu7VTQkLjCldgiL3m75oRLf644TAoBNVlq1EmR0bTutXxGlVeHzw1zeZR1JF4AiN6wkcOTwyaShNrL0gx1LwUHVIUtzxLBpJ0fmLB7sgGMef8Uobq2F2JpngDmldLGz0TL4Ht73OX0TVMKvU90729yvvWS9NcdfjafMSPnJbyQbYpumI4eRtRUdal8DbvUjrVSx9DJWwxmBPXr38B6kVsVISwYfkFxjy5yLPtz5xRdmh0G7AXA9/DYrRr17yXr69dsGDQyeCinfcoBU/x2pkDEdp+dWObUqn5xCemY9Hztk5eG26BIguqsAY1cOFGfhsP+XXDakhMf0YGnRFQ4RugbHzxpMnYtkZFkOM9pN8unRpTkRX+Vhms9SFjRDuPyDH1Rp6VIIO9tNTAFZX+dfaEGbYWiteWMu1rs+xhD8dzdOyZyrn0ZOoIqKAUrH/i+/221pz28PF1DaPjfkcUHH0+jsJdG6gYCvmRcByMad0zIXojZgNitlg+lSVaG6gA981v1pIGYgakMCkxMAReZWLr7tMhUNEBUXj0r9vD8ll8PkCFdJVm5w/UsfH01py3Pd7Kovk2xrRdQ3ecOZBluIHchBHUwArdx9y4lSMqbPgzaTjNGsvOqlkNjdojPhid8b1UR6U/0ipGT5QCxnFUtK+O6SeQxrQ4GVztcS9Kq1NGOlVr0crT+vyACi6FzmDXIGuid4lbLUVnXdAEPcLhTV6Ak8mZPVzTem9ltcrTp9hpvrGZ89nTi3rmZMupyTwlk+XTVzoi1o8wGRRT7q0FVBQgRMZQ06Ftvbkn6NWOws0oMjziG0aWw0hr3uMWjSDwj2l0LM2P1/4wozbqX8Q6RkVld4IUylB00EueNCxGZAOTlJ5Ye9fOl4EDgxdSN6jL6pqoVgKAlOhUE425HincXm+RXipE7ON3pmdikeh2P17AOF79FJ1N4IGBKCi4bXT0FOCeisuARAcnWHOB2Tg0agNyNkoaLhAMhdZhYFckga2zG8lhGN/cYvFvrBkM7wbSeT0O/s16FqK51UzY3THjO963GXjNBvIOaMp5ZVniQF1cO+7hsMZhI2xtlDRaFnkEkMWKkCMV1RYBTI/eQBQUgQTKb6YeA8DE/QsABhRiAfGULjF+rNGlFyI38AfRGwInz6wWh8DcnFbpkpEnoFWsbyMQpGwNMon2EYbKtHKIjmBBdN5TPbuDy1EAP6BnjOJi/Qmm/3oaQAU3j2f58POqTm3YOq0WuNmAr2cRFTPS+tlXXxIKFC3MVBAXFrPFtH3k8XiLB3Oxb2AjRuPW9ECMzxaCrKewTu0sC2tUUMLmQ3K+//XGZAJ9jVfarBl+dHc9T/TdNPVOZ2Eil2mRfFzZ6JulpVp2odzl0EivZoK07oa39L0L8UohyoPIPjoxomK4Fn4xomwubeTnQ/fZi3igiGVDrl9U7DJtDSuAteENNy7KcFQOZM47G2nsrEJETUNwO+mIUiwCKuK41zV6lGwthZQToELz47jWvKJ6u+1bM8W0Yw+BByl3/LD1g34sHCPP9TZYGE+g2SxQEZ6TMp91rZwCKJCxvdeuuzYTZq35rH+RD3M1Wgmo8Py9DSlGxtp1AYp6H3b2m/F0f7VySHX8eggYYE4DY2MwJMQQ26H8c7nePVsml9GWh/xvCgIrI9H9GW6WyH96M64dw8Pp/fI5ABXo0sEQHW+2vyZbJY6p/VJyvFzQayNI7/mORbM6ACcMOt7ia34T90vk794+mgPv5vO3rTmoEdsEmqwaK9fPuKXT2tMEKvqb+OqyYjrc9UC3sfFuKGx6SO3skrW6Si3f885doMMNi95f5VwoN9eSVk0Gq6fAgk8VqAiynGpZIxQbsHgsMtfXPNZ9YylQoXbngIrPCsZ9PkAFmaNmuazRTjjnaQMVveUfHZxPCwOaYkyFK8ww5Pyp9B25lkqr73eACm37zNflmsxpPUWgYiTTsO0L31Ific+WYbPo+ih1kbURriL0jKZOgO9kRKMhkt9Rpg3OnbiwTofxflweUUGyPj2gQjPAuptns+f0X3f/VjfahiSo2ZCNymakR1/naXN7pMs68aRmOv1ZR8A9952xq/Wv1oKGxj7N+xEV4XQzA7Rqk1g6I48umAgQPyyYHooRDuAXpbfC7/AOL2lxzolq+74z/rQIhhE4xM9rYy15vABKBC901IyACjwDoz0AAY5ry6IEzMDuaY4wP44dxm/WeejxOKYt737QCYZo1PIADxWHRIkBzWHqCCSvfwMBrP4D6x9gn6kOg3S8DdQN8XRVNOIjqkDggIVL5VRUZsA/O7OURZYiyvVEM9pbuinYnujZz1RPKHZOYMoiBk4ZaaD0SFZfwguXM21eSoeHR5YyTSCVwKcS9cL56l4d9dQ6tVrh0o1LT2PlgqsAHoxwUfFoAU0AYzCfLJ+2FMXDehQGujnvGnixrVRLpe6DgAoW5OaeBJ/YOoCvtkAHRqkoQoTgj9uXXOQiYgd9EJg4YWH4zS0DIcAfrE1BXtB5gxbOTk/S1s52jpAR6JPrczh5qvt6t3bV2Hki9leNW5s+n13lEKCs4V5+BlQ8BcX6WROfNwWKBnZloCIan5rLWQnlnGjRtRrUM2IvnPqVgYoMUkgJzNfTTs+jG+tUXeAn4fklF1ahse1QTHubDofO5CuUofa1OKQwvqjyRINUXxGaFjDO3XhtEx2cpEGPbqHmgWFK4TALKDPb5ftRkPdBnTDZSjCPoxGksCnVAm955uPs9SRC/5255MusaVr0TqABOSeCHdtVuhedaDxs9suIh+Lnsc0hUFHzeLnsKeS6s15d1s9X+obLFgAV3l4dHVG8AtoLWd1BHEz/IuUMU16z/NnFE6eKqKh4rKYNcTfx30AYLdnbC+TY2GhZ5pg9MPJFm98pzDePvgJo6r21YCijiQpJyt9n0GBwS83RR2Vg/G1wyUddn95PvAj6hEu4+YD+FWeM9khz+asYxv8YGvbGVremGY1kw/LhijezB9TTjqgw60PNs1OgQrfkIt9quhvjVx+NgAo+pVzE1ZW+aaLZqzP7Zn2jtp+4re7R4bOnDlSM5jEyZOW1qekxP+eBwWgJD67k8ZEcn0l1NBQic+BJ/6Wx0WiU+mk06fXqmpE5B6aeCoiOtSL6Y/r/LVAhGTlzqIy05viKrcKa1uuxYbQ/mCFQER7PO2FuLE0dt/L6ct6XY8bINWRepKyaeSP716Xr6CwfntliAj8JVg1vhlfmwKHea8NjPbFAL/Z3LDCanTvCXDLvNUQX3/L7mj/n+HU0h6uSRSl7lHaFW4WyS0CFimovASoMrLFrDtuglzxTnJTUT64X9CItP8fUTxIDpcpBFAtjCpblrNOQcdnAAzRORzNFV89cAT5NQUC0D89opTqCYRhGyXOr/THXhxlG3fBvBYNDWiF9Bw/z+mzhfdrmMfYPKrxhy+iWVicN1lle5TRUhlRYsoe4zgAjMFM+eZ0Fj8KQgdn4z/vIjmCGc5UoHTNwWwqdeA8RZaKRH0OF/q9i2SXTA2upsV3th5a2MLha+qL9ffOOlwF5y6II3PBvQNKW3QWREqrnBGIxGxbBUE4uAxq2ua5lz/ndy/eRTdIiJNwYb8XCGRkB4GoLfOHRXSiujALmAC8kLwD4wBiuewHmB3ABf6P/WMCahaRpOFchaTynOh7WBu4VWwSJxJMGcFxcpt2d3XR8cpx2d5DyiFEe+Hdnb8/lJiOQUC9Cq4bZYnzxvFO9C37m0UFu/I6f6Xc4UGkPlmgOyhoBpqCzaCJDur4TmEB6AKw5t/mDniyYvVFHVJwjeoW8yx+CVvobfWHrHhwckM93trO2HEEUvK5i4rmY9j5pV4pzsw/wu2pUAOA7Q2HwbcofAXp4joWsNba6HhkL1Ux/hmeLwOKgt7Z8GsUReNKAMK/l8Qyo6JL72YdfLgr4Jp5J/fTk8b108Oh+Ovz0YfrP/o3v1sNfYKirQu8mhutgvCl2wboPHABKl9Ptry3cKeB7fE0C4lx55EdPxyZvYd/YnkWxi8A45M4VZAGd1ueLkdEWa7rE4BzV8WAQdeWjhhA0OleWinmqGrbl5xO44Ab7rOzruKB248cbDzkdJMVpKBj4wlQok+VL3Rq/Wu0NfDMTEO1Fk3PfNiwV6xrRdmQ0KqG1aq+O+Ag86t4OzUYqNKhWj6BH33u8HYsrpSKiqoN1GatNy1LCECcMHXTu6nLo6+ZX45oP4rLm5fZ93NkxOljLWsS5qLHAo0X/7m+b3uuB/2yHmB43XU+7eGR5GIC5vF2cIIGPV+3dVV5c7ffdaBztadsEDqb5ftDzvX60ZyYywcefSdWwT16m6JD3ucgxX/Vc12dAzYrebhjJu6bIC3ILvydoqIlF02TgJXu0v9/HQEVzES2IXxFC9lndbgExddgxr2/vp8IdJ2xaz7e838jxfKY2dQt02x0xbhhT7FpUtdcaYFRRUVZk0dvt8/Gq3XK17/t7qCev12x/lufXNEENQ3Si92w95jV7CExe8i1zRRqecSRxmE5hTTLNPt6bxNzSZAPAkEHDF4XbVg85Pjui7Ghg/eftktzreI5vekaxODRbLpdbM+U6Jk4m3sZKo28oxivHABnFsoxai/GKztnz9a3kXkMrec/GFCRqLQ6hSPHxKq+a96oooer9Sn+qbzHTEUSgIurf5lacpaG7sVOHnaHvyF96FX/HtZPXdUvDto1Kvq8JbFRtyWCiD9fin7koqvVluBkV3VhIPc/1hca7O9w8BmdwmET/14YEc4va+a7SG6bQKd6QF27sSGAFP9Om73NHjlj2R7WPmFKFKXxomJOgUeHxDpc7HfOwXQ8w/d081KVncK7RsNzyZmaTkDIF7Ux438mWI+Qr82mz77Iup/69/oNSfsGYeQEDJ4oJX6Ttze10rnm7Ll1oGnXMsKfNFkEvdBlctQSW3iakJ4q0r9dBEdElnYxWn1T01KBef4RXaa4z/hUQ0uU2p2FPFtCYzvRSZiCGSdsLL1uxZzfmKm3OBVLpuOe87kWWk98KaDNFEMlmnJp/N36y+ByvFWPe/YzewLsWdWJ1ZMi9tgZmaPUICm/SCn1vsOg3zkMCkDDi17UmYPQ/Oj4iL6M2w/aORR2ABlsGMpQC02bUR1RFZ2/ZuC0KA0Zv1kqwlEr2CwGYtiZAyZYGYAfRC57qx6KDWIMCPwAJthHZsJHSiafcEr/LgA7gUDUaLBLoFCmLkLZs2wAYtA0AwYz1Xly67FKm0cI+BDiHaAuQFcW6DYwA2HB6lvb39w0oQYopi6oAAIEIC4sOYBSKpbo6O7c2LErF5k16GP28ELdlXtHphmfSRQI41ONLoykcBl0Gox3M6+j4OO2oUHe6TEeHx2lvbzed2RoVexK7IVeJl8QXR0dHxh+sQ8NdIufEOD5FhKilE/DMFscBsOjo6NBBqVofzzIYa3d8bOCI8aHXx2AqJ46rgMiUNSYHwX9npCX43kApK+p+bmtqIBLACwOmsN7k95L+zVPB+YYzwNnrdOoIEE+DRFpXpZHLd7OqzgejSJ4BFf1z89mnXyoKZC2AxwyEyPl5evLoXnry6IN0+PijdHz4aR7x7/79X8u/z5iA8zN24LoeZf/IeJPz8VKJr+50k8tWX9XOl46LURGxPqHzkZo9CAJCYn1P2xtdKiqDmLrLpQakWJRxzOnuJVVKdXXo+2Z4Q+XJ4MW/hL/ypViqBhWXPAVH5adN8bmRkbenVPeGkyMkJl/Wl5KpJ++S248YLqvkfYpkQ2JNb5JheoWhjl7Uxdn7QeXVrPb1Lw5gFT1lm+Wn//vUFFLTiePSKZbVxyEnTC/sBCpyq3lDhvDOwhz8TZfadvN2PAJ0f2A9j0LF7B4UpEo1aLsfFB5t7nV99lzB/y2H9Rop93Xfw3mOlB799Rp3vMpAEt+sPeDDaPMlbNrPdN+1/FEvWQVsRDk4mEK+jPSe7RnkqkvfEoHkOTY7wx4a7KutEuSXZzCU+1NV3K+tOVGJkz7NVo1+Gg1TGo1eWzQu9CLS+jJtuKZZNE3Pl95YtePid1n+jgxTs4npO710Ab+m/pG/NhvVsIrYq/Z24MXhSTFc5vH693UdmQKXDhqt9HWVOQPrkhOvlpmUlySFnzOtfDXAhPOlLOj1Mup5hk7D/bteW9kU4/mR43HDqRQ6Fn5aNYe498ah9FP+nF+BnM8YFA35uUc4BW06gzbX3HfRW7Ac2WNDY2QDyQD7V8aDzrDWWzlWKev9DOlBG1VdrDwYvSUHszbnnqS9PqLnbk/eLduptYk/a3w+gaFnY19TH3Y5KE1UeR9Xc5gZvM5nGfrMG9vqp6mWWv1yZLNK+x3w5WjHj3hjFjAavLQKZFq2di7zekfUMAVNewEtL8dI3Nhkz8GFMmpIkfnh+2vRSL+ctvPyaYw9jd8bRYkJIBGfmaE1gxfBC94LlddARdnjVvDVTx3b34E6FI8hle4sXUMth96aa08G+lq9Ci8yvLuz40ZDvNy/N41kivZclk+SD24VFDDRAkV+6PIf0W6iFvjZnNP+hUh1f6972mW9u96xommPCQ2UgEe/pyWC0RxpdwwMmPwwxVjWPJ1kcobKFMyDo84Lj3QDDxwUOYWhfAtGZRq68R6KIV+eI9USUjht04AbDOR4DsZzPJyLG5unuhvbbRt7Gh9P64S2bGXt85LHv+wJ9k6DrkcFDHYqI454xpuBWsZl96IXAGOe6l4gG+O3+hSeEsgKLCtCwvsh25Q7LtMZsbalOX46eKE+CWRwDFZjxOtxxJRLO7u7lkoK74LXlQpPvJqjL0ItD7Ea2mNkABfR1AMDzAjWk04hbZcZDsSfZR41Gd0QH1ItmYPCBeptoEj4loNfm+no8NDAFKS7Ymq1UpeHKchYa0Jpr0gX8kGRvxifDHEEiew9q3VBMMuKmaNeyzYLzFukyfFx2rQC6r434XTl+9oiYi4RjaM6GB7x4m0zfZtjtVW9LtJKvG+RHyqYbcBSSYnFtSYQaE053SMtWQydgAZpQV5Q3Q3wF4AXgFJMSaXUbXLOpOeh+OYZUDHY8M8+/jJRgBv4/PTUwImDh++nJ48+TKfHB91BCqioLu6z9p0SXVAMOr4J7bQYAxVZWPSOy3jrGQAVQyqHtDh56FWekvWAij4tAlHiWDtao870CVAhJWBwAWqNJ/p7Xm2NdnE3becxBWOfnVC9liJtnoJhb7JIpc0pSDG+UMijo6BiasdUtD4rrAQq1Ib/q2aCEZ8N99qPtGnaUXHb6jV/Jo+pHXJfaSxPSXX0vTU0Po1TeujylXsKF/Oq9xYtWEQPGsTqSKbAb27Ency6BUH8geGFcAVLTubRZQ0VOrZNUBtQrP/ieWZPrDBgrANSkJvEs6O91k5yzH+0QcXn5fXk5VI4AZvVHOliD5PnvnCgIqR387kaf8hDy8Lq3SPqcwYq6E0jBb/e9wIqIs8s1wR68mR+zdR2C3JOgZVmFNbVylOkfqkBKkZ7YtVemaPHaB/1ZIEZm0eNDRl9vANGThkT788VC7oUqChA/ngdxjYxXRr93Y1oOtZZJqBCM5j2M2toH8yz+07PSza/36d58RkVjyviT2YNl1mV7F3Ns+vI4pqvZtYBF1X3BC1kmR/LcO3WBSqCMaGQdA6oEP0o8Ct6wDjYGfZqqvbkx3LJlou5Bb0i68TB+9LV4dmz6osEKkYzHsmIEVBxFYM9DSQ07uK/CFTEcbXrO9EkvkCgYnTmjA3tY4r3vpFxrfvWQNj9vIGKov/N33XinlzNL/0dPAuOj4juNQWK0ZcGPaSpgSHXPIRRZBn55D2/fC1zy71stB5U1dYAKoZjbaIznAwqJg3DHrztMU4Z2nu8MZIp3HLU97Tv9Jl5QweQJDo0VvIgL01fh5fxeWI76VWpmNQgrE+jWYDVz+icFkopkCqC+N1S+q3bbvJ8KoS6zAePG63BIxeXLC4MgAF/X55bsWeMbWd3hzUU9DfqEIQ6KngHIIHJN/CaFQWHgXsz16cAGALARXyI7wx02dwwQzQ8+k9OjnmGqFbLQqBCUQyxdgONw4z0ACCBqAfMEc/gB8Zw2bjMy/0CaXdYdJw/9d1MxnYW7qY0sAgNp1eOZkEhdERYeKQJxmA6r7XP1EixdeNPgRIeXSHvf7snbW3nPvAsAR5GVhiPK3WyOzWAv7Ge+I5rQccY8E82wjebyTpF/z0AACAASURBVFJo7ZTC0jCin58xwsbGjGiUzY10gnlZSieCiAIWJWOwhjTM87udHdLaxuIAgGgXbRoEVWWs972bLqzuxLGicdwOIUCmOIAyOsz4z/dGjkB1uqquTwQmMaazcxTqvkjPPfec0RV0A821liwIznoRoCVAGkQHCUwoNYQYjaOoJANxkNoOUSS+3aw2y8mxgYIAKvA30o4pbRcjTsivNg7YN54V015DWX326M+dAmenxwQmHnyQPn10L52fUoDP/QCo6Bnmh0YEdx6rv1d4FFHjWmD3Cn/yiakByN8cpFMYXwaDkS5PNh4YHaBiRJSRBW9UP2LQzkRNKfrcNBTWPdK7xmPP9zdcw/BSBjay8lkb1p4GUNEapqZ8ssoAH45b047rmRU9r8pPUx6ym1lL3dbo1zQ6ua23Y/S/7Z94fQ5jy4Y79O38lJvpeeLKWNzvq2NGoiKSL/ctbdY1LzQRFT0GGlmuKpVoLD0smgL/ma2k4bVBG1HWVNjkoMDo0LjWGuIz3boTDR/2PKBL4bSVRt/WU5SLJoHWJVa5yPSN01PzdM/IOHqX5M+XlgUghcneRko7880sdnlrUeSds2+Pa0citlL24z7gYeH+P1642hvppl3ungHjqcVvpvKsXFyDELJfTZEVvWf3Utu3jLJiG8kKLcoqfiq8sMxQO44UGBrswyKN9sSyvuc93Xur8sUCFe0Z0DsPymdj+hUCtnQaS/KeVRl9qT//fgVQUUcQVtw92ATrni3jAILRLtuw9Ijxst2kJpwAyDNUmgCHy/Y2xciSudqB1gGs58Y0GMOaQMWwqO/MsLNkjGqMREmPpRaBlpViuZzA+dwv3o/1EJhqwwwtztekNn/a/TSadk/LjOdaPeCrRVSM5Nswr/pgsMt4rh3xXwWgos8269OjT1gzuK3JmcO+Bw2N6kSYBtV7JzJm+L5SkZsx58dcNunvdenE59ejCI1xkneU6zLUm6HQjccy3sbaGq3eJM9kM7DKgtjIXH13NVClASo0gOAUJbtrdDBpWWSOQhGoqN5rgIr4XQQwyud95ihe8rUE60dBzuj8s84CYQ3d0caM7mennd0So2Sld2bCZnaaHpt14WyT3TC6em3HaAg347/AVgAbqNXgHuMGinlxdDPSWtRFAYx0DhuYYWmmeH9jTv5QTDsDYeTlJREV1i8KURvgwrRfFi3hBvNcnJrxENXdnN70LKjtFugJbTleP9UccDZjttf5oPxyAM8N3RZN4Dcd/c57Bgks/ol1RpC6COCHed17fYrszBadE30MGVB0mhmnhnoh/J71Geq6FYEvOC2bew2+8VxXxIetuwGHaDBEDViqI3I96G0AlUdcIA0T5sG6D6oXw740L1tfRX/ldOAb6fTsxNJFkZdUaD2adYpdxXh0gzLOIh2yXkkAwc5/Ocq5XHVYIx0fHacbz99IhweHBsidoNC7r6u9Z/Mm8IA0WIzsQKFvpPli8XOm3iIYtblNHkQ3ltrMAR1L33V8kvb29z29GVPxqXh3rBlj6d/wv2dAxZpawbPHP3cKnJ4cpoMHH6QnDz9Inz54P10A3V3j50d//4d8WpecFQaXeNVUNwxpoyBxicomcxr/6aGdlZlmrLbJhxEV03byJ9W5315j1gQq8uvxsja6GvWJ3Y6rREcMFNyR4ZUuCBP/aGu/yjternpFCZRBTN6oSh8Rx1zmNQp/5loumL8fylOKBG/YHOnSuVXHF+0UCkbg3H1PGS9zr5g5M2jLN+1cIigAXukkO6gsovH5aESK/biBqaXJ3I1lkjKqvfUsuIS0Bt6WpraYcT8MaDO4cFXNGVBRPolGhomc6BSxjiw1urgMAVNpzo1hXrlgax7UGuHTOsVI32Oeby8a04J90b1OD4rwgqDxwtl6r+kSGalOybuAN+bOhVXzcPme1zjKyI7xb1gLorlK12K7I2/VkICKEJJsCnW7lSsyTGXWIjnmdOIZNZUFPO/UUSt75tZB8riRv5XYCGOeQ+ZXrVe11lfhjQXyfg09Y51HRw4MczzVb388hz7AoHNK8kLvx/O3/n3Uw2gOozCnoQeoTbqcMVx2rif3vI8gp34qdSx65/AKbWXxMi2y94fWAFToYso92NYhm93Ii8f1NB5s1+4qBsAyjvX3XvXGCkL3Wo+UXAcnQdIOl1A2fKouwZN4KXEtl3d9KrXqROyHhpn1OJMlg6c/fWo/XaCipxdwW6631rPGWm/PAB0Z+TzfeqVzNV1OqLLumEbrMNfOetNeCBbGgQxW9QpAxRAIHPCT0sP0yNLjwJ4eVrx5V/B4A1SMttuYb8Z0Gm7dEFGhHOpF/pGlYWDDzxmKGlt6nymrC8jAd2bcDHpTHO8SoGI0VqXIyd/r6DMjI1PFxDQrc5ETc7SNOnYeuwy+rZ4dSF6vy/ydM26nPkjhErhJqV3viv56ywAKloZBE+Pa2901A+lUh+oAFRTd/L9qfuyd9GHbBBBgtKdnvdUgcG9/GJlhbIbX+d7evvUvb3o0gM+Zloj6NN7LhnE3QudrnpGDRm945gNAVNQDBkkDvQZeAxUxD3m7dwSUMHUSokBQO4J1HXACWn/b21bYm7y9SY92i+rwVEGhroNTqLAoIhLOYZNDxAL5E3O0/WTpuDh39A0DNeoeZMO/efvz/GUB8XOLhADIY2Yyq31Qal3Y7ycnud6ERVUEAAZ0sjXrOAlLk4y6j9JeslZCXTuGJilGPKDGhq2n00hgksAUzNUAX4+mYSQIi5L7suY0T5ZSDOO2ejG1vSrisJktfeBGqdzuqfMSDfqRp2jJL3zMMbHOBgEGjjWDQ825QJ0oGVCBKBvUBtnb3bMC3gAsEBWxt79n68a6IQQkDIywYuoAx1CbhNEWAuAYnVPGof2gOiN7u/slsuWCEZaMoCgRGaLzM6BieNo9++LnSYHToycGTDx58H769OEHXWPK0vH87j9woKLjzTRuo6hoEujlkKhTP+nCEtuSsair8Bu60c/7PFQuKuVBVyD+SyWgA1SMDD1Rg6gsqX5mTwyjM5R2MtVGkRmTYmP74nt+UexZacxQHNaCYj9cBHigxZ9p706vgB63z3dTYbV2OhfgrJLe+PW0Yy9uL0vZtAFq2iid6mreaTMG6lac6H/IGCRgpBSUKk9HOmth9dkq4+TgGl59XNIT5Ut8bclfTav4fMO7WfFEK4785wYbo7+zUelvEO1g6+wndz1D/dW/yrH9aKoY+4Et8/guQ+3fp6f8kWWQCYl6H6m1VUDFcqO3ireNzDHt5+CnaBAVudyryOVC0bmuYEyqBXK15ENuDnTisrtc7RjzjayD6Y5EbIlMCamf8mK4gAnpTT5PoKKcUTVQkY2sWdlvzrt8Wept1zovMZ8IwnIirAcrIUPvaonwdJ+4ktweD2HWvhV4Z1UEz/hEHe23qed2XotBzYnuLNz4vi6R17Tr+UaiTFgGVNhVtHsO9sc6otPaIx3aannklFh9u4BXzc+cFc2gR04uo3VY9/l4WRdIMTgi1l36xc9XtJkzEvvlumo4nNfdlR3JZfMwDOeyg8Ijr/JZrglGZJ4VHj8Rcj3buuj8XUWZSWeNxiFD4ohW0cqR51gAlVXdV8flCCQZnIOjtq8KVPToPpZ0g94HdJo9+9drakjSuXn3XxrLoVFbV5lHr++YJ77+fqzc2JiafUSQdgQkxJZXy9x16Wcnx+y+8P79fC+57HmX5FTi7wIqylhhaEOKF/wgh35rdDNtVjJA41mTB+ml7/IpXzHoyMdURFuWPkcG0s8CVFBkcc5Gg3bPe/8VXePSrYrib/wV+7yhu//UhtGzq4iLNGYZO22MKoxeMTEnwTngd8W46U5k35ZzWkCapQbbMqM6DKkwzqrANWiG+gD8DGlqSmFhtKZoOjSKmgRIaQNDLgy6xWjPqGnqCARCjJ84Wjf00+hu6rOfW+Z971PJHvdhHctc2RKAAoIjpZizoiBgWJaHvM0VKZ+Q8goe8gaUMAIDHvL2uxu7Iwtg7qABDNMaPzzlUbsDjRGo2bJURWhDqZ+UworrSPPVzhaAJo/GQESJGeB5d7Bi8jYHpAzycXthZwOqrIA1UytFvm7TWwpYwjNK+QQaoe6LzmnJEhvWlqfs8hocFsmCOXskA2hr+3ETdTxIa6U50t5SWjlwn6JBQFMCSIpKCI54vm+UYiqzs60j90uJKgGQs1NHRTQ1Ki4sJRf1nny9yYvIPaEffg++I5iEFFVI+6Xi6lgrzJORDaANIyoEaIn/BMAQcCJNmCYKz3M9UR9DTgqg4c7uXi6MDqDM1ii/z37k0PRXGqiwBTg7SRdnp+nizNHD7Z20ub2btrZ2cj60viLx7NPPlwKX6eDxfSuEffDxR+nJg3uDegPrj2IEVIyUKhnPy+blZi46R7Ox/XCJIxsBFfnzCykjy9TvSq5ItFQhW1cAKhqj0djna4bmPvxpOPtAGa0UHTtSpgpS6C4aAgPVwxO1oKW4b/uuQxrb2eS0AnnBs77AX7LCWB6YzK51Ss75xkcGlXYUgQ/s1+kcyhsjg0dejPKoNTOZQKgpUAzqWUE26/Coj96422c1js4cqvVnaOQwrZDG0LP65vGp79CwzrOWjLGvasjmYlBPLMy/1GHxR+w0j3SNjGNqTliqrO0PaGqqT3eDxQtCtRxtJip728NHnWHbFVl9Nezv8SVABS+t0iHqS1ZPZkbv6SJjCz2tPdE3yJeSmazDV1129ecawKi3u3qzr8+BPgXnLl/1kOL+dv6pFrU+U7QXnyZQoUvddK713CJQYbQyxbfm8bEhoV7/4toT9k4cwMi4cBWgoiuz1vQCHgEV6wAYeRzRQ6uheu/cHI3fpjAs99vduGPgAx2v4SRhx1cj0/qiovp0XXlDGah+Akif+aMed+2hGXfaqOeRnrXuSMdO5YqoMEmGiKSJoIl7vI4qi8SLMjfus/H+XbAgzSPT/UtenWHBxpFCDZJ+q99tz8vy3srR95ZuKVARAkPtWLF95LsjR665N2Rni67mDsX8uNwLsUBsrqOftGtRmdDCl53FmAekHCQjA040gdaVZS5Ccew8MZJD/VVcCVRo7rFGRV9UTu8J2mBryv3ZNR0ZlocvDfSC1YzT4YL1aJhp285/DvTrdDFO/TTYmU2Uh3Gan4++qycvliEtI8ycAb6v6s1D+S0f6m8Z0SSzMY1CD8ko/ivPbswVRjZ617MwrOlpPms7MlugIq7RTJRMF6jwdgVUyNMdNB2laJuTqRirDId4Lqef8VRLle0i3qWa86zNFM1rQHQoIsBSVrwfi0NPdlgfpnrJ3KpClstIip4tDc0APMme68GgQJ4suk3kTLVrRndETeTi3ac2R6WuQR59GI/NUO0RCOJd1mBgmiMYYukRT8M3Dd6KWmYkAujO3P/8kTFX54jSBum+VTtXFufN+t5Y0hIpUohgAT/nZzQ4A6woqaIIvuguxogHb8vHp9RXGQQJcod7A4DHbjCqs41ioC9/U3xw/gA+MDeME3tOvGq08T4M5HGaY79Z3RZ9p3H6nd6M4W4kt7oHlykh9ZJqm8DwbvvZeLAATbZPLIqppM1CP3hfdOIzl2lvbzdHR1gRcqvzEc9+3qEEYmgPlugtt1uFtHTn5yUCwkju36FGilJ54WNEIqCmiaKxeH122jrAxLIgTMGE8WHu4DMCB7SPFXMLgVu0A/ojagKAHdZSgBXGD5432iAyBACTr60KZ8txI+8HpfXyxq2OiUX5oNj3hUUkodYL2mH6KNbzoGwlkMp98guW+unk8JMEz3sUVb44P7F/zwFC5N+PDZTAZ+enJytTBqFyOgCLLYAXO7tpE7+Hf+07/L29k7Z39tLO/g37+9nP1ShwcvBxOnj8kYETKIZ9dnp0tYZWvPWjf/C31m5XMleIH1MG6QiJqVWklFCBX2LYo8CIhqvi/TgxmmvkXWVcBtOgTczfNFfQoYyJZzjnO5pTDSLU6mNXwZAAdTdpO2grBW6qgkrxCFd8B41E76ZeSDcPAN8uiGyfDJOUL1Hz1OFMrbw0kFHeqOC60K9u7yNDyWBJZh/vfNmuuwx9dqGPvOa0cAWtamlSe6UZW9tt1uziF7IM2JFfGsinYEzsPzPJii+kUHpzAwNvPdqodi6gfXu5q6bUvr8CqIg8GNody4b++JbeN0mO+YLxy66HY/EwlAE+SOOymplccQli05YeDzlvzHlk2YAbmTJYxtHqrskB08kv4DMLQc8D4C+tMak2PIZu8ovlvWoQSC9iReyb1av+HLzbWcr2sl7GVbc/BSrYWLnArj5OW14YOFqOLaNV+Z4F+3duSJ/pTFw916GLfRt1F5d+4LG8oLcVQnl1C7yOTWlab1/9JePnmhJkrSVT2FoxGnTJE1JERUPW5728qykq5aA972YYYCIvext2HIW3eEyDB+cMyKO2x2cAC7tyHbxAZgWs1TJqDLr1e24NSNZL1s06JvXg2W2cbp62rLdDI4+PR92ZPu5rl3NBc4FGhYlz9IQ17AZN7aoeQ84c5vK25biK0tkcpxVxekBCGUVNx9ZpKq/jzJZee40G81ulN7QrbsYTWjzzj9a6jDvMFI/6+k7aWqpAxRfXfGf8+HryshhNl+1sGch0LmdpPTP+0YiCpC+dy9N5TXqY97cbgOP1Z115kw3/oUD1LEVXzVvzCXJ39MqI96nX2YafRG/k+3Kx9lWRVMWOULS5qtivy5F1xzSiq52knca0h1h/gMZoGISR4sV46hzFupm2xwrfwrt/VLvSazJZm+71v7HBIrnVWgX52HMitM/smTplrQzFy3YEn4Jnvfou0w8ZGJoQaDwf5bf6Ag/kVDvmwc/MDSoG3BuTijPnCAuv34B3DajwyAaeQzR2EwyIujV5a2dv12pL8Bq/wegN1ZnAC/6Ozlz0LXBFAIOiBwwE8vR6opLNzwzHrJlxcsJIIUvP40Z2AHCW+ufkJJ1bHQIWOMaQVHPDXtrYsO8wR9Ae0RioKbFhKZ9Yn8E+OyHwYKsEg7l9DuM3oyDARCjcjX7RPgzkjKa4SPt7e1Z/xHhRVnR56PvdxPjQwTtLR3SB6AzSGONDO2aYT8kiKI4wRjeu29rAQG4psI49hRUiBRisoL2BUSqtlegXzzik1LK0XQ6IsH/XLfysorFfhn6m3rVi2w7Wqwi5tkWsmQNAYmubbSKSBDxhRv2zcy82DWAHEREEfJTyaapPl+jPHF2mmhq2cYIekovD8y4qPqPIwjyY/ky0xljIS4yAQaFsATKUL4isEBhilgMDJAyowJo7L9T/EpRFyizr68tao+L400fp6MnjdIR/P32Y8Hdh8HVE2dN91gCLa8+nvWs30s61G2k3//f8swiNhtRnJ0cGTBw8upcOHt5LJ8dPnu5iDFqLERXxkaHhUJEKlYDXYVcu+Vkn8SNyyWTU5wVQzOqFVl1svr0CULFEVa7swdHbIKgai8CX1qg4sExRLEkWtdEUPetG8FQJhr2ihIVoCV+HaU53b9cE8MjaWT4Puiaf1ut5vYL3goSqI+vhcQIqC8GrLu/EoXaMk1320WAdqKjo1HRy6QVLy7XdO/QDfzKmCencAOBjaz08AFTYV5VhoNTymFy2c97naL/k5V1KZ2sUHu+5ctAGdhvaFIs3Rn66OSfD5KtaFLUXkCm+HDHfXwBUkA7LvZzjRarQYxVQMS3qvkRetc/MGh7KxtYGD/OPlgf8Djq1EqplsMFebQY1eqrDAeHNvnQsn2pXzNOtrEWUHzE1XQB6dYnnpij7ohLC9WwI1PbpFIHXJTI6Xlzr5+v2C1DR7O88zplIgQ5gNXs8jqzMOWpoGQ80m7XmkKEle8kJuWCXtAaB0N/QI3AwpnXy7c/OeThsyN8+TSfgktpYM92LjsQFlAtygnI+83qPEKFGBYGKmN93FZ9cZa1XSZb2QC3Gbu5wvD/Ij70EqIjSal2D4QrijwxcS+RI23QcWgQ/p9tC8mS9teDT/v/eaGSP6SoVcJcGGj+KYSAqHFemocK4E+1wnG6w9BlHN78jR7O23PMbNIRRRZVmVM6eiRNN5q+4GqMeRPfWuWe8DusalpfvdalFY1/p7ho1ulTFc+sCFcNpj2vrja4NXyRQkdfIjWwyUI7WYkRx8XJFFs8pv95O9Z6bFFBMbzPSt/qf4x2B0bSDb/A2Id2pO8lpW3ZK5GLavj9dIIxBgeFO7c7DjMTeR9GdnNrelORQAaQCCKo0tXORFqPUo0O6joGKuBby8AZlVBQ4SjHlme+R20CBEImOqW4CqKjOrfhXLxqLMpbTqO/ytnZrzLuVxFE/jqBFLTHp+V+OmHLO4DcULWbEAcB4Gve51v2fnE5JfIfIhWDctZuP2yFKceMyb4wZHv77+3uMrriE4X/bjPws+q5aqeJlnhkw8FMfYmQqwYlNAxlgMBZYQXAKT5ybcbuuneH1I8zjnvd0RhEhdRDBDqU8QgsCQvg5Ig1ogJchG79bzZDLS2tHqZsM+Dg/tygEGOjhRU/PfAIlmgP6xXtoA+0jYoU1CxR5whRZWBeLurAzlHJDdEbKKfRnQASiR6ygN9vDv5Izkp1MAcX1BWCxu7eXI0vsUweWAEQAkLD+Ly4MwMEcAKYA3AHIhIgY1qJgfZnKMddlJHnUwSmv/6D5ZVuhRUFcpC3sLczPbQyKNOEaMq0UACEMH4CGdAqzkzf7SHUuWSeDvIQ1Nzllt3MWvbZdqUgJk3OsH2IpqDw6I0ajEFzkc8YHW5tWp8NSRTW2sCxbvBbM7u6epRDTzdtf4D8OiqBNKzL/RQMVmKABEU8epaNPHqejJw/T0aePO5f1oaz40nyxs3c97e7fSLvXb9i/O9efz39/aQb5OQ7k5OATW8vDTx6mw0cfpqMDrOPP/+ezAxWeViWfT3UqDAq2+vCSkBkZh0pR5/aaFduJxi9t10i/+YiKJUpmD6hoFdoll9fW6Dy+hvj442UsT6l/5awFnLw3OLuINpfLRDvzaHCbN2jM2M04Sjtg6rzDFPpSTGsFFSOJ9Ft8AZxji86t6TKDAf6ie8FkA/wkqgLj9ItrBjeCsbvHPBPS1YbMEhfkpArNxcNnBDLVKWYiv/fXc16SGOULZ8lYMdwU+qJ+p/t4lQqnBRhkJAk7IB/4/RFvpFq5XyUhpbzXoE1cnHqheAdYZchb1et8tFi5JATZKOBJAGE1Bii+MxJq/arC8xNo5z+64IXnlsi93n6WYlfJrch/VuNGilsj1zuVs0fh7Lo8DMHXhiIFjJsVLi6vaGR1kZe9pUuTi06XMIJ1+W/d53vnYzlr+syxZA6r98UE/fxSAxVjL/1oZJ5GDS6gQ6OaLH9j/YiKlfrF8s6f4pOFn6I+NDKIXUUkP2W84qnNnV6hrWcom18oeheOxWk8Yyyiu6k7CWRPUhkTF3az+LE1ZEhftbe7g7yWmeBABieBFtLpgoaVP4pycsaA1nGYKOfHdLKL9dTFdKofNMPQ6F1bu/KlZpjfaV5cO6Ji1PHc5hocR18UUAHqmMHTN15OP6SN2KHtMFLAn63I8jSAiqiCD2g+Bk+KAVtGrmjQXnqe2808pokztcb1mqEM6Q9WOfgnO85TshRZJ72pRF6wSzI2l6iO4pKiNWbN/jdDQ/5MRIXACfNMThtp/xo8mZGJhM5D4mkYI2mM7qd7g/5O7/si9y3VkTcQs1DYZ7N7CPNbnvpplK5Md1qMqQ9O1KsXbTcthVkXwqMMzlhDArVJ5oAKq6sg/oIc39xkFIKlgQr6tIN3EUwp9wbSSl72LFDNdF0V8G4DhmGYcyVAUHiPAAsM6ox2gEy1ehuergr/7qAA+dmZRyl4aiKkpUKf5pUPgACGZo4HwIHqIxgtPArj8PDQvrNUQSfHZsAH4ALDOcaFQt30/me6H9AJBn140AvAODw6sec5B4Kb6o+0YfFpfK/aHbuIyLi8cEAGYAijRLAGAA0M6DhjWiKlScO7GLvobefgJlNNYT/gHfxthbA9XRMoLZAnpk1DZACAAEv/ZIWnT9MuAJhzRm+wKDqN9piVQBS0B3py/3If7e3tORizRXohtZIXkxaIx7YuEu095AmelYwgAQCDeZkx3wFsK3TeASoiUMb9EiNvouwqdWxsva2gN1PGWf+u92lf5AhWby/WQlEqL9UqofBIBlYB1MFewdpkYRHvUiG67ucOVBw/eWwe9kefIGLiYTo++OSKqs8v1muKwGijMQBu/OL9XBqYZFEvnxJYwloOw6Z/zhNcG6gww7MP0gzq5YCJh3I5eYsHV/192fztlC9ni2lHDa+E1E/JtiL10wLlOl4iceBNvNwX2osWAxXZoK7ZxA6mnRksEAeZ3eOa96tXW5Ujrl9/QnNGg7Y1Oi+4ikP3BEJVyuk440G0mPUnw/QPZPRtGipAhfhWRYDDg42hmJBL4fPaONUZ6WBM2Rumagshk6Rc20cJed4s6Hl1OS0dZS/Dji9k+W6eqosMQpO6D3OMH7/rKdclWmBom4jLsiZQUXkeZ+qOx2vGj/ksJCvZcmy0n1zbqplF0135wlQ2wX2DvhcKnprD2l0h5q7GxD8GF7+8HUL/FW+uJFVW+PKToSle3vhBDTT50xGoMEADRcpNunTm0JOhq8c3faKmRS+ioly0x7Sr17ftZZ31rKTGfLOxm9EtfygAxoa9tajYXRoH1Gcu6L0+Pv+IiqsAFWtRYyluVvNzTq3pxFwRUVEMDPVe+mIN+Q3wP5FN7R6Y4b8Zg2NvNT5vw/I8B6gIbe0ZOnrnKmOtKRU833v2L8eBefGWLGG6ick5lhlmtDYjuSWZvI5c66y3v2752fPvTkc582RPR8qUNrqi6N5jfpJuSkPX2MN9zZ1+5cdngYqmVVE4GnmqQ2G4RDNn/NgiPJ3TzBJ/kUBF63iQ7x+D825toMLvOesuMl8rxu2rRlQIxKAnsu5X6+w36io0kk+TpY1rc/SZ8QKc4QAAIABJREFUw4x/wSgvHjb10I3GNCgWw7GNIBjYvmigwsYDQ64bQDE2K9BtqX+KR36cx3j9aaTFT6m3oFpTBSjIwIU92b+bD8+KwRergIrpvhTfNPcVuxeV2j7F7EMgCYZT8+IPtQN6VwfpzOalH9IsQa2BwTuCqQSpODEBFbWNI9HYv7VlKYtk6Obz0zRR9rkDXwCKZNTXgQLjPcAF/GCt6XkPozCLJOs7bjJeTwxoOFNEAw39lk4I3vveDus0MGWUpSRy478VRoaB3iNQ8L0ZtP0nGsRjH5cJNQ8INBiw4O8QgGExcBQxx3fGs94nmrXoEKuxwXFa6qhjgiB4FgZyREiopoKll3JaUG4yVRFrJpALAOIg/ZTGgXbwHmpHYH6gHyNtKO8AShwdHdm/iqAQ4OOSyNtijRt+RlsB1wT1PE6t/AD/ZRon7DGsB+QK66BsWToq/I3vCYKwVgR+8Hs55xX11LtDFj2DkSYOPNh+nuoIOl9AQ62pWT5NnhDYEuijouf2PYBOr80SdQ+AZqCfrfX5Rdrb3zfAycNKyS0NUIF+Ln8eqZ9QUwJpf54g/c/jjz63ugQjwfdl/xwI7N7+82nHozBiNAbSTH3RP9g0xwYqPUrHGZR49EUPa7b/H/3WqEZFX+kpiocfCqZ5RGtVMTZl4Svv9CVWUWuvHOg6gOp9qVuL/9vViJ8uUBFTQsTL0JKL5VKgYmrwjGvQWY+sXzTPxQtm/srXaHLnbNduAbu6ttmqVfjblCQHJaTLS4jr0PMgi8pDZWgc7enFE1JEPpjSqQYqyqU3Am45bNpet5nUh0G0Zq8cU7tusTaF6B0Ox7wvygHIA9XXokqLUw+rZf24xWad4Coy6Y9VxslsLeAgqsc7c86sVNpXSq3oae36X5fx1o2oKEBFlBE5OfAkgYUBFYP0CKOd0F6Cs5xzgpd93Cj+/qCijHhBLM8Ucua4pGYIK+TBgq37mR4ZdT9rBPcv9Y/SoHf4j3ww6MTe1z7X2l6my82m8wFPFo+tVTyu/cU+WgNGDVTEsPxI2Y6sHhF+DiUbnZdxCkvO1MleDYNZY6ifiXfal2f6HbLTsqX7TMMcBSv1xeUVEM616d2LqOgQIqR+4rf8/yXngQ1pzXGNzpYx7hXGrA6H58eYYVt9awwSX50Nluh0y1svZ3oxWJWUAUvbmR1TVH+cdFqH/rLGizn1kVzkMXrbNudZvearNmM51ed4cCy+OHJ5wYpOMDYxFzdpaMYnGUgjaBF4mmfK/Hh7hu2la/PzfK6qPxM61tqAnrFGSVvTYuVYQ72CicjuMJNRdSAMvkiggsMS+OYex562pUeDUeHlrmbsDlgradk8IFpVx3c2yE5bm42Ma2oagr1nA6kGg22d3WwfzPDAaB+VNEmFYko5g64j35a9loNeeGKFmgTdGhVDgvf3djQAx1dN+o14FoZgLwCN9DTm3ex1ART1IWOkRV2MalQkT3njuf1pqIyG9FomrY6CVDRGvCX0CTKcW1M/RE50pZX6vtKNqAhOAszxX4MDU8grS25LJwTaMbKEqY8ln1TsmClvwhxVb8JrBDBC4NgiDmCYVUSA9HQtKyOM/Ebhhn327WnT/B5CUIfGfouyuGA6JrZHoz/aAmgBI7z4UhEULAxNGiiqyNryNDxoSzVOYEg3T34ABheof3JiPHFtf99AH6bPknNfSR9ltNlkNADPaQEudDbg3kMqK9aVgCG8RJjQas90VayzYimHrMYHdROrw+FFxLVaABuU/sqiPFA74uI87WOsKE4tA3soyq00S2gDkSh2VnvUkYEsnu4IERXgNNXFgF1XICWLrPvdy/NzME0U5uQyHdFMVu/l0gAZ9qPC6EzNZGvgRn5bRwcQLBrFCmUjFRdripSE24VXQRcDWjzlmoETFGS5FkUNshaZIvAI8xDgpWiPeOfHnE4FiJ2fpfMz1qiwKAsAXBbtQZBkf28/naHAu9FG99+yX9Xn51KjAnUJUCj56OOPDJg4Pvh43bPv2fNOART5Rh2M7Z19Fvze3rV/t/xf/I1C3yoGDmQOBcLnfi6MeU7SBQqRWxHyExYg94LkF2eo+M6C5GdHT9Lx4S9exMuPfuvXY/DD/O/5Fl9CNGW4ycpHN0TR8xf27sN2lgit1gb0VQnGreLR4N9FNDEry71rWbkwBbesaXSEuowKTO8WtbSgYMVY7u2Vnd10EIfxhtQARfGP86nnJrL5KRl6C0bZaOm207Rn4IgK05R+oh4dmEtallYZkvKn/HvKx6gcpSb4oZw4qCWlVBhXpaitugP7pTNchTufdFRqrF0mHHnOpjQxjsJT2/MmGt3y/03s4PKyqOVIXFf9Xg4Y4jwMC+RPeYbKCj7DBbwAHJnepd6lvZlJ5cSoVU1/IN62JmUFwp5zxW4iE21AkWcL5QsftHNueCm/EkKlZ118W96vzQ02Is1F65jT9EbOKLMp3Q323cLT1Obse6uit0cSmbGgiuaoryE2usyHNLSQuho3FTn+RPkVB9iTdb0JjJ7jmPhtKOLe8Eo9hJpu1RBXdW1rVArdVY9H9spftPwz/dtAilamVbKjvLMIqAhzL8/HIsBa19KuPJxqg+nStQln3yr6xe/jHFsZP+Lh9S3LC3fDmo/ls3783jDlxcpzoW1zjXXIu02C1IWKbQ8mnSk/Yti5iuDjfbcmxdwRRLKgc45nvYx9RvoVFWbsKb4U66pYcLAWQ2wt8B+fwf+5riJhro+t7SKfqpPH8xdHZxEmBGqO0/a4CpK0L1GDFJ7MLWtBay+dzcTbizKiJ4/ai29N7xnmd1bL/TSjrDnRNLUiZX0JIlARx4zBRyC/OIOv2oykWRFP0XFoSsZW9TAI32to1HTbotHBQQkZbZSDW59PIytGS8d1L8bT6PW8ao5XYofP9FI0+FYNBb0wzn34/Mw50Tsqyp5tX5wWT9YTXzRQEeW1pUb5rEBFVs+uzhcUbeH9uQiekTHdLi6UkPmOYEDF3Lh651HUAUktOZWNkOsxYFrvd7vvITe+eTvDwCuZTtsBZZ0EvvrWGVdSP0H22LSadGhS+3h/7KdOmgUqELXsFwijI1LWmgEUxZ3P0vYOi2nDoIuaCDCIMh0MDL30HmcR6GJYZnomrUFJR9SmJzLTaLVUlMmj1eP5xm/je+VUctp7K+WZeNKV9uMaRrCi5RAzyVpRcN9J/osZRbcohy0iAtcH9wovHt/1bPAqgR1GJMBOIMM1CxzTGx6e+2eWIoqRGvZj4DTGQTqY8Rce/4gO8KLWiF5QnRayiw5dgQh4loZzRWEAfMBaw1DOiAEYp8/Mk18FjmGwPz46MdsFUilZvQuv+8DC0PTqx+8wzusMx9yY6okFkA2YQU0NfHZ6aimn8IM+WUz7KO1sI1XTpQEO4BEUyUbUAoCOw8PjXJDZNCcz6IOWnrrKU1khHRVrZSDlkqc48jkbGGIRGXSCxHysOPY2oi3KPj07R10MgkCYgzjHokG2dxg9YimIHGwwwMqqYbvTAPovQAXobVEqZwA8zoz+oD1hAERrsAg0HRAYhUBwBOmluDc4vo107rU5jk9Y70I1TYzGkDce+WE6A4ACRMtgH3u0hdUL8fVQDQ9GbkgX1Y2Y+rLxh0epEGAjDVUHrshJ8AwjfMjLTLWFFFtFD4p3fYAl50zB5bU6wMM2Jy8ejj0G3gRfIaLE6olwQ/i+KDvW5o5i7E+nRsVlevKQ0RKHBk7cr5TGke7w7PPPhwJgPIEZG1s7ZGCAEAAgTk9njo7PZzxfRKs/+oe/zoAIv//m3yvAIWwIQ8KpINkhHQooVZ7E+ZBR+JVmp8s0Wb+6ZKqbQY4Hy9OfieQX3bxv+4YBOzjyxm4oHBSlnMKqeqRcXqu7dG3DyPSLt+ViZA4NxkLkNv0iduwwcKFcvHb5ri6H+XNN1fLxZUIHyswXD+7xWblMx283mO/P9J1A7yy1Sv0JUwxyESTmS4TAZUEiKCIs6qTcsQIymFNwqohGbokzrNSfYBWpQqirGh9EwEt7pYh3UdgKvTIfzNYJ7vBa4FnxdD78OgdLxPELl8lnJxpdfL8w95hjJrJMOH84J004oTUK1nprhw3ipNu9Vq+C8kAWno+8PJJk4ni1Veg+VtJtB3Qgzv5+H8vQzvNQfGfzyfT2Vtm3bV8EMKbG7HgJiRdL1+ps20cZbDMut4OF7s7z9MiyWazTEDwaGHXv6+27aPjU/IuRp5Xx4bKQUaUZbzZf6mVe0tw1/Wd5obGUIZ2f7ryGmhgAxSipI53D7yMGXnSoh3Zi87HN6vOZtV7X6rwugDH7fG9crTFk9b4dAhUVWBAJ2xJ/dR9jCdUC15Kxmdur/XiVnnrSbBGbfMaH5mXseo2PDVajY2Xqtzbam1m9mfGC75+ZflaGFWqPvMHu9TeWSIYOr2UjWp//l1N2zE09/QxbvVyYe73U7eW/hgbNPod09yP0kVEkIm0Lg5/VglJ6rkSZIiesoKWnuYCRDIYGS3vhBigZYNCDARieMkqayXpyZX6c5cy7eqqouT3UO9fMiLycmezJ0XEyioKYFE0ph/zafY8jLdadxTBoY8xogy76xnwazafuJAFkjGqogwTdbZQFEyWP1++lPjcM1yMPweBpHtEbm2akG+lBI76JHvCFTajHW30A2y/MYS9v6uEu9TzuBP4KHYZ9u3c9yRSM2/Y7vee5j8vdxcbrAtrIZjbgcFeTF7QXoI28GYEKtt85VXXf9u/Kni13Qnmac/jsu80nnz3abEPVyjq8oLkvaXCmo55Sz9CzOwM25rFPx5eWPfG5GYX9C8xJdRjKzAT8kskUDSBwVuAV62lMfxB0ae/AwO13Q9lHWJAYKXLgYU+9+czqC3Bc9EAnD5mpQgWDlbbIDiMvEmzFn2kP0HobkGHpweTRzkgEKxK9DWPseUKxZjxjufi3dwwkMgDB+IK0zDwDCkT1G+DJ9lY6PDhI165dT8cnx7mugc3XIiLQJ3kOAAsM9DgjGOHAYtwwxnP+tFtp3xIw8zRpl+69b/WTtqxWBaIjBFpZaqVT1FFglAbnybmLHjDYMzqQfbMYeKm3USJPMOOSAogABaJOSD9jSYumgJF7JxvnGQEgh2I+J4AQY2IEieZIflWqKTwrMEIG/mKTIt8ZWKWaFxn8wV2JxnjxM94DLVRI/vT8NG1jLUBvLyYtftP4VIfj/NJTp7kA0hgMEEIxc6vb4CmdHJxhDRTfyWGT0Um25LBWrRTyGkAxghrQLyQb9S+XvTCbgd7o1/YReZJ7HNEQDsBB1trannMd8loRpLT9fXaZdnbJ55ITtv8g/8/PrVg51ln1UvC7QDZFdUlgINpiWw4cVymmjQF9+uCDdPDw/fTkwQfp5PjJ6Gx49vkzCvzcKfC7/+jXOydaUCga40Bl9DWh5KF0rohwR0bDS8lx6GI191cUvZACBYpAlXe8eC0WkLx49rdttpOZqC9RkEl4yLtPQ+8plOsnyO7StXzYXkoxUgi/8nk2mmeB61cufyan0al6CrQcGnY6Q2s89c2Q7l4M2e9a/apdebAr1ZNFTTCE0cAJCxdkcSgcCAoh/C//2/96MgApsVCOwFWmJPg7xmWOjktQowEL/zRvCIZF6j95NUDAP3nyxLwgdnb2vRgVvSqee+65kjfS8hzygOoZxTkHzzHoNDCvAMv7yJBcHHL4G/+x6FXx3NAhRqUC4aQM/0Rfyn0Y52Vh6O4khMPu4ox9m+fF6Xn6+OOPEwp0YQ6gwbVr19ILL7yASk6BvUq4Iwt88eJjFyG/7Bd6KQS75NMuSpCpOKbAlXyd2jjwrIESCQ14Mz188DA9uP9hun37hbS3t51u3X7ZlEUVDbO+5e2RmB8zh7G68mMGZng2bXnY7flFOj48yiG3AEhMmXApc3pyku5/+FF677330suvvJxu3b6dbt++nTa3dlyR3Uwb8EwAT52fmUKpdZBCpjWIFymFziKv5jtv3U23bt1ML770Ynrxzh1TiAUynB6fprMTel0wJyfHL16iJw0VuzfffNPW7bvf/a6NsShC3OAsSEZesosqxnxxkTDHv3znHVPMfumXfzk9f/OFLCf0fPYe26ACic//9P/5l+nWrVvpr732rfS1r33NFPijo2Pfk8UrhkpsuCB2jN29S7M+E63aTW17NmBfG64oSsKVPcc3o/EntjVqX+sY36suw95m/h7eKc14FGYbeUJ9Y2/duHHDeRTrWtMoX2SafqaXeT+FAIzZcViMW/HZ9r1YUJ2GjJDLVqnpfLAjA0I7rzjmdt35N/O95nMoWmMW2pcm8zDQ+iB98CH30cnxZbp376P08iu30vsf/Sw9d/1WeuvH76Qb+9fSa69+Nb1/72dpe/da+vZ3/mY6uUzp5HI73b/3YXrzT/4gffXOc+lf/bVfTT+++1Z6/4P303de/0564eatdHF2PV1e7qW0cZbSJjyP4HjihutcH6nm0B7tS6ov7GfS4+QYOYw30p//+M/T/vX99PDRQ9tX8HCCLP7mN7+Z7r75k/Taq7+UPvzwnv2N7/NlgoTNnRtgH9Zya3Mv3b9/P33wwQcs3OnnDc6uR48emocWZKjyHGMf7+3t2MUURQrJ85tpf/9a2t+7bmceeBUXaBXwhEcWvLwwj8PDI78obhl/4xz56KOP6F23tZk2tl0Hu6SX4c7OnhkODg8O0/Ex0mGcpevXr+fzAIYMjBv0YKg/z1PlfLazEWO9tp92tuBptpkOPn1iss3Oh93dtG1FFs/SJx9/YjnBzbtsZyftX7tmZwaoh/2IZ/Hdp59+mvfm48eP7bvnnrtRnVWgI+akSzPeg06CZ6VPgAdQ4BGegpK/pjO416Dmg3Y4VkRlb2dDDzz8Prx3z9YWeYRN9rsuIVkkvQD/YtwHBwfWloon4t2Do0NrY393j2fAyWk6Ojw0WtlF2s7gE6YB2N8v+gqO3gQvTBpGrMDm+bmdM9ZvMI7MyYhWdm8qp7PrC6Il2kdketRTdb5HHQZzB83EE9oL7RikR6F/PIOxY6+I10VDraPaifqedJr/8Hf+06AH8oymcWgGN2knHv8eADo6t6NsXYe2c12u+u6z9LNQfPeHMAeSDIGvUVPrjYTN998Z0aOOgCvjuDJQ0XRv5+jMYjEyWlqqGwwH97HcTijYantpzTnPARU0lMp45kCFFXvtg6MsluxUDEjFaM5KA8SVik+5MVQxdLmgset7Mv5GHSp77bhh3g3VPR0U/dmdM6Pb0XrNBapGY/fcYjrMuElId4W5W1+ZNuOVFigAfsC5YGBTACTwGdPgOC8IiGh4B++bMd3rWhC4oaE/2jAiDSRvo85LPbE/3jMz/GZC2QjwF9Ma8T6Auctof25RSPQUlxNiMfjTm58pjs692Lin6jNgoNQ0UM0PnAXw4scP6w7sMLVWyOtvv9uEWU8Bdx6bk8uYar9XQEWyKIWj42Pz3kcEDM55nj/lXkuvfb5otUdcd6I3PmpPoIYEUyep0LHWTl7/BhQ0oAz6Q7SEQAB4ykOnMCN2AI4oNzBB/itewfQEvOOsww90NuNviywgw+RIBrdHGN9ZCizaI0x38ALlsQ/bBwEEw+8CxlQAnHZu2jMwP6ul4VFEjAqI+jTHpUiHsqZeYDyAF6U2CO0dinrAWlidk2x7iTzvYIhF2Jyb47jZTpDyyZ3QwJ8biLTw9eUxkQuc5B3Gzxs55HOBgZ/3UIK5WmvtPe2lIifYloqES89FF1g37kXsKdqkzi54d5BMpO7AeUovtVoUBnJwgcAT4FvpVXiW0TvUjezHgUKhotqzJmWWAhUIH3ry8IP05MH79u/pCZXQZz/PKPBlo8CPMlAhqd8qLs3fMvTn3IHMoVwOkNaLlUK5/tGhHY9gPsFLResREJ/nVtaPDvKV7j4uaWSKzoKjAlVcGNtw23mvq1x3nndtqiiwhSo2Z8+LWAJAOG/SdqpQMiQftGponqVqXwmd8mBvfZiqhamatDbRK5J5GHnw0qDK6AkAEvDEOLfDE8ADDgB4TOBQwEH1X/0P/91kCFK25Hlgghy5EHGQDIAKXVBhRNGBoXbwPvrChR2o+/b2XjZQ4EBfB6iQcU8HejywybM0/lPZpLEgXsz1eXlWutIUqCA/e4ocO48Y7mgGld3ddHp2kR4/ekSg4saNMVAh4NC9Iyxk2Q3o0UAsXqThjGtdGdjsXGauVobuBp6Cp/kmQjXBC5vp4f2H6eGDj9KtW8+nvf0BUGHhwjAmMtxUipdN2RVSM9BubnheyvN0fHTMIlHoGzzvlgcz31xcGlDxl3/5l+mll15Kt166TSMhwCuEGIN7YHwDXc/OcoEz9StQQCBMnB8UBtD57bfeTDdvvpDu3LljQAU8cUyqbaQEoOL81L2Dzj1kuNp2NVAB49N3v/c9AyqkrEgpiqBX3AdnJyfp7bfeNnp889VX040Xnq/EnQybth8DyPsv/8WfpJsv3EyvvfpqevHFF9Mrr3zF9BqAL/hpgSfNveXv3pnVXo7ivtN8wE7mTxJAN3ly9drUe+2FNO4fvafzhopfkV+jy6ztPRTOa/aWLZW/3r6Lffz8889Tbmzi0jjtR7LBmgmAbZyf8t3ynFwOVOQ6Od5YnCdzapfxRA+rlrYx/7atUzhLaqMCZA9Duls6G/06xho91xopYxsbF7gEPEnv37ubbt++lU6PU/rAgIqb6YOPfpZuvvBiuvvjd9LeJvj7q+nho/tpc2c//Svf/kE6NaBix/b4j//4/0pfffGaARU/efud9NP3fpq+9/p30wu3bqd0CSP1fkobuNSdpMuLeh5xbeM6ZV6twCaetwIqjg5PDOB74+4b6eaLN9OHH36YvvGNb6S33347ffWrX7VLxdHRQbp980b65JOP07e//W0zJleX6hkevTjfTD/72c/So0eP7LwTKAwD/IMH9w34R3u4uIAnARLs7e+lfRj/92jYxjkNwPra/nNmDE8AKkzu4VyCkX+P4egbm+ng4MjOZZ2DOAsxJzN2b22mTQsuphBjccQ9exYAx9HhqQEVeIfedpvZ4ABZCToLqLDzygHubYz1+jUDKvBzdHBoFy8DH/b20u4+gIqL9Oknn1ihR8g8zBdzwiUOZjvRAG32gYrnrG3MQ2dVBCog90Bf0Aw/aAc/GAP+Y4qOCwN6ZEDHfGSkF+iOuUiOYQ4f3fvQzqHd/T2eUXBE8MKd+Jv6ANNaYNygE+ai/jCGJwdPbDf3gIqdHV6kRUuMQ4Z8LBNyMh87SIS+pPfgvID34hJ53sqMdYAK9IkfA+CC5yhoD5rnsQadJMqNrANkXYVpM6SnYPxoJ6aciPSV/vXv//Z/kiMs6Mwgh5AiKVsD9qy5eU2gYnT2VHKgJfSaf3+Wtta7wTQD+0KBivHIR/T4IoGKqli2h1TYOTOI8DRHDLs/FK9r08dH17cuOWj4nPIzKUFnD0Yfmae+jHsD0mZjvXSPFXyaa0q0z9kdsoxKnsyKqJehTYZ5nWU6geyOq6K4A1ClAirwYuVqz5aCTzP/2iiRD/YKrZn5X3srG2b5Xe9HxmwaG+msxDoLnnYHxm83sprH/QCoUH+ljgHXifra9MfuH1Qm7cso44e44Za35OYEa9kfxtmiiAZ458PYD5qxYDaNw2ZM92gfNLHpEWt2R5djwvkZoxXgXODrhvOK9T4YIYHPTXfA+eRnLt7HuY27PH/o6AiDb+Wg05kcaXFhwADy+tuZ7ZEgjGxg8WuLoFCdB4seoWe8jNEwBuM0pXMC79y8C1MH0DkH/pKzifYudJdtFED2YteqqyAHTXMO9D4xO9VUIO85bXFfzU41zEKB6TJtErz9iwMcAQRehQlQyAZDe5vN02xKVOWUcYJRH5fp+JgOewBDbE3c+E6WoiMN1iIXpI5F0J2Hi5MBwTGkrNrb28/RBXIALHqoF2B3QI5ABYuW12P0KBMAIRbtQH4ASAFQgym6YGOCGYHOjlh3RoS43h/4JO9c0TbMRQCY7tB04uQ6WK8WgVSiyrTnAIpp/GYbOTu3dVL4GbPNMDLF1joAj1pzymTcCbnHfSdbRIXthZ3tvG6Y58nxsT2DOhWyFdjel3OQbJxzQAXSBSFi4gkiJx5+kM5wG3v284wCX3IK/Oi3f6NzCsajsT4msyHV36KxnEZr7uz23V4ecUdm83U4gCS2Y5luo/x4PQH1WR3dy1IKVLOIxq38RfAemcyjY6VZsK4TJRoCKStbrfrhoWn+sT0XaFmfzxRrwyLAawMVPAj4owHoE6p4/BS0LsoOzw96O2B8BClg0CYggUMangY4QAAW8N/z9N/8T//jhHrR8IkvTREYAhV8nYh+SQHQXm7RBi64VJzojSnDwTpAhYyhOnijQTUavWKEQDuf2hMQigppboWpGg9bnVq2s4DKIw0dDCG7yJGZ0qOHD83Ycf2558zo0o2ocOUV46BB2pVeP+Q0Ps6teBNgPtFwQGcqrt10nNrbuExspQcfPTCgAhEVu3tb6faLr9AQZQpgAXQyULG1nfNN6zJi3CagwkJhz81wJaDCIiqcv52EZih655130osvvZTuvHLHoks2YBCzZ5nn0Qx2UGbcOKU5mvEHRasqQ6Wz5yW9JN5+64108+ZNAypeevllAz4kIs6O0aa/j0JnrvQVQ3oJIX7jjTfS8dFR+t7rrxtwIN6RIq55mQFNyiVCoU9P01t375pC9+prr6Ubz99gSjYN070zrD1cwFwB+hd/9Mfp1k0AFa+ZYfHOnZfT88+/4HvizEOhg5SNoflhhw6NAf68FC7tk2z8hdEyXPCgYBnfjS7HwaOwBR96RqB2XOLp3ngzbV2CgXq6BGo8vT7AS9evXwtRfuVimJXZ4O1VLhqFgC1QQfC5eNVEYViPvQbs43cl3QHfnjNgDY0IvH6G7gtQ0aXhjKUrXiZb4U6g4iB9cO/tdPs2Iio20r1799Odl2+lD++/l166cyfd/cnXwgJgAAAgAElEQVQ76eL4NL366lfS4dFBShs76Vt//XsWUXGadtODDz9Kf/qH/0f66u399Cs//DUCFe/+NH3v+99NN2+9lFKCkboAFekSF5Z6j0zpXGptxQuiH2sGVEB0bqRt84L/yZs/Sdeeu5Yef/zYIpT+7M/+LP3whz9Mf/In/yJ97WtfTSdHT9Le3m761re+ZXJg4so52FOHB6fppz/9afb+x/6H3EGUBYAPXPR0XuGMQxQE8mbv7e6YbOW5lOwZAhWfGL/ikgfjGHgNF0h6v22mw4PjBG80nEloC+cHgArLzY1ifhY55GDNhb+L9w5heAZQcVoBFRZRcXaWIwAEEmBsdubjAulABS5h+IFMx/mOMxlRCjDyg4c+/eTTdAqgAvmQEVEBwIebNQMVoA3WQzQpERXP2T4QqI5+ekAF2sRPC1QoeuLgyYF7ksqwQT0C78GYwUsqAb/L8wuLqMDYEaqPdVd6Ip150gvQPkAQtVUBFYcHNqa9nd0qogIyCR6eAEkFVNg4LBc1C33i/MI8BRrByHJwcGjPwBD08wAqaOjwiEKX8xiTxtU6P2grFGMH5bGcQXpAhQxieDeCGAIq/uk//I/tjJSXZ9S5inY7NfsNwYohUEGjMtfXdYHsQd9Kv3nZPH16/pM5Ob+qreZG1X18KOK/pEDFcM6Difw8IirWBSpMX3JHJ4EVAhMWL1IGBNqJk99h2LM0N56Lvxgnh8oYuw6uxDPHf4545jtl1Lw/8I4oncvGk9PquCEwGGzlnGfPw76gmhaDxba88dZn6NjrGfCVYp+gWx2u1n7fVsRVsWZOInsFYvS6Z85/T2sUijbjWenBSp9jaWKkKzaNqX6KQH7KQho5s/xuBxAjRQWqzFRUh3OC0d6BMaSKMfAXhvxzRiBYBDdqKFg0JosByyhq80melswLTStq0lKLbREQotF+285Q+x1Fg0PkhGS3RVXsIqrizNYEfcUaCDT6lwhN0ZnRHeHHeQztshQKecruzrARwGDsGRBwZlvUnuv/dKLiuBG9gbPTwH9PvQbDOPqC0yU/pxOhzicBLpy/UjJ5keptgFRnRgdEW+Qi4nCitFoHHtHkeBMjNZT5gLyiSA+mf+K5Q7qU6AfxuN2rPXUXxhyBCnvGU14RVKJDAwz76IcgEY38ihgpkSMdZ9iQ3kk8irOe4AaBDo3RIkJcMDDVEiJ3PBLEv1M0QY4ysUgdgFle1wEpwlznAq15f0daqVMCXttNQfAGqLA9H4GKCD06Xqe+GfHuKdpCphHd2SRlorNzTg0GW4qiotzOCBVBNrKii5EiRqfsjEzWNT3U64Nknnd91faOgxPcjwGklMxpgQqCE0zp9OmD963I8rOfZxT4RaLAj37nN/xC3SrwATyIZ4Ln8pSAp7E8vju9CEyM4GrPTptGq/GwuF4UhvUZ36HGMfY8ydftLCe9v3DMBaAiTxPJHCc/c2pab8V7z/dzpvNthQJGmvTpKsUp1puKIyg+GL21GHBnQSOqB5TDvwhnv5hZaLKnaDJPOhijzqwYlXlPnJ2V/05ZNEjAxX//v/4vfiDWqYbsYukGWsvNB+O4KdjsvQAFTrHgTaLLqi7wMppGoAKGBHwuT1LzkIAx1S+ZeqeipV+6o1FZRrlolDRvJVcqI0ghxVRehSWqgfzRAwB6ERVmCLHiURvp4cOH2VAzAiriGKg4qJAZU1+ZZ1OemwMVvl8qoMIKZtGoDWUvA5LGptiQrsQEoEIRFQAqlOLCHneQxIwRSP3kxpYsDhQW60ET8AaFkneE1E9QLsOY8Y52E7ytM1DxMoEKRlSAn7YMFbK1NaOZh5C6J49FVIQw2nbtwT933/iJpax5+eWXDahgVAcvcWfHp+n0pAAd0dOBMqwAFXfv3rUcqq9///sWUYGfotQVLwko9ZEHkPrp7pt3bc1e+9Zr6QbSfA2ACsgE7EOs4T//wz8ygOVbr75m63D9+g0zsOIHhr42nZnWqLcPRsb/3rOZhthbQTzTN2nqISZebQEPjacnsWK/GRgJSltXymG9CtRK/unXYcyvw5D7/PNMKUNed4AjgN2SAzWQIPlf8sC6xTWnfuqDGrE4aQ1UVGCAj0UDHYX72xSHLna1Vx6FLy4uPI0mKxXkbW/skebq09YWQMXZQXr/3lvpxRdfSkeHl+mjDx8YUHHvwbvp5ZfvpL+8+146+vRJ+qVfumNy5ex8I736re+mY3jfbeykhx89SH/6B/8svXxzL/3wb/+t9Bd3304/ffed9N3vfzfdunUnbWzcSOkSRm1cNJH6iWH4Ubb0eGIKNhUDBu4bR0dn6fq1G+nx44/TOz99xyKWcKFGVAOiuH71V381/f7v/376wQ9eTz979530jW98PX3lK19xT6mgAzRrENfkwf2PLe2TyVj/D/sT4AEM27u72wYm4LyCkVpABVI/wQhAGXYZgAqPqLAczATFCFTQ870FKtAm+qLH+mZCUA3v+vRe291BBAJT+Rwfn9mlFiAB8znjksjUT5CVMvbLw9JAAxSb3N1N+9evmYc/+FjgM8AIAyquwRPvkhEVR8dM/bS7m9MpRaAC/QioQD9LgAqMU6AFaIkfk7OXlyYb8R94FTRA1AM+lzECnxWgYjt78Vm68ouL9OEH93I7TAuoHNCUFRGoQNsYh9I3aX8+CUCF6QXHiNIBPfH+NPVTC1TA2w79WDoNB43sfA1pFVbJgrg/DAJx4FhnGg0R29kJIJ7pOsuifBRQoXO/PVsFbkg3Ev1Fe13q8W9M/RQ/19mBMf6T3/qPmO5qo6SUZPqacgjp3e75UAmwVU80jj3BnWf6Zv/u8FlAh1Wj68m9zw2oGHmbj65MM+fR0nmV56adWPODPkYFpy0yuGqKf+izuWjC/rnCCOUaJBzfx5TvnSmjhsOfJU/rvMCHeYoTPCZomY2fZrjr1zOQfmlXbI9CnTPYZ2cbCoAyTjci06AfVs2NzVF3s/1g91DVAyj6YtYnOjx1kUq+fs2Za8fRSw8oOol7jQd9Jo9MKaDsDsIBz+o63gYBV6Z+wg+MpzA2ogmCEHQYqH78bzMqW40CRlFIbYG3v+5iI1kR9axVOhmLV295itoLu38BaFdkgUVReOooA+LNwM8ix2ad0HjlZBPGZ+l64dluxYPdyx+gxRlTPqMxACKmV3rb5hhh97BQn8VpYM/a+VO87u18MMPu1DrELV9SmVlKJXfO0x1MZxMIDFpgbDLaiw+t1gRX3c9xRfCXKAp8JbDFQAMrmozIAIIajDqB0wdrlljdAY8isHu4gW8E7wSmy57G+yCN+IgAEW1ypI6n5mJdJqb8pN7GqAujs4GRTBctN1Ma6h08s6Lx1MPE3/a8y3GmhPK0VOd+QVKa78DABJmYElp8yGLQRa7onkYnA/Zpe8MjX1iHhOlmjb18zTEWAmoEDWz+0KsSdVKTkxYpc542kCbaI0mZUruW//km5kCFPeFCVueBaIl5KJKFUWdTOaD6LKEZj24i/5nDhqVUI9hkd/Is25yAl9wvikrW3VfOySWVWAEWVadFKci0dqbewNYBumB/AagQOPHJR++mT+6/10ieZ38+o8AvFgX+83/3N7tARTlUa+XKBA8C8U0PKxeyqCBMKDDRz/yoyREDUbEhvBzRyup3Ayv88OiBDEvJb0bW8DDd9vwI7AAK6+IUVZ0N9dN4WU7GymJE0x8fWx6DK9ED1+QSYrwUqKgDY61/e7UY2/iZR6/4gcfQTipiELRmZLGoiVM7uIF287+zdHJGT0z8/j//n79XKYF2lQxGfnRl7SndkA+jGJSnxjcpGjhkcVnX5Zj5pqHw0ejBCIxNM/zI0//Cc2qqX7XVXoh1MBAwoRFaXoT4Tm3r8hwNmNFYgTOF+SDpQTgxlDsbcgmY41JpMhBRAcMM5gVjUQtUtCAJ/o5ARYz64JLWERWaR5zDxSVqOzD1U+UZaR78yJsIy9aWpWdBRMXNm8+na9d3LKJCKS6iByTTLaGIGr1CqwuBaYHkPxi1cDgj9RO8b22sbURFSunRg4dW/+GlOy+lOy+/bMZ5pX7CfsrveHiojEcCiWQcrGjnWwDGojd/8hcGLLzyyivp9ksv5fRTlkro5CydHBUHBbXBOVGhkkHmrbfeSgdPnmSgQp+L3+RhC0OgDMWmnJ+epjffeMMU4G+++s30/M2bOQ861kvjt3a2EH5eAxWvffNVr+eybUZUGDoJ4FHBlDLZ8n2UQ+1FKT7bGn/ys7ikhdupLWsTUYFntW96QMVSca7xtJ677bhjzQyVujP54/uk7Q/7C8AX6spYUW2/wMY5x31e6OkXJ79A8ZLgwHqIqOjRuFw4ZTTnU9VcmvMlftdeiHtrV/cb/xqD6fIe1NOx3REP2OdI/3f2JP3sg7vp5TtfSQdPzhOM87dfeiF9eP/ddOflO+nezz5KH99/mL72tdvp2vX9dHh8nr756rfTMSKKNnbTo/uP0p/94T9Lt57bTL/xd/9O+vM37qZ3fvp2+u7r3043b91J25s3LaKiABVKIdChXbPIEQAi7em9hmJ3H398kLa39qwGDvLNHh4fpv1r+2YoV3TDu+++m1599ZfT+++9k15//XWTy9pTmVahJgW/Yx/Yg++9e89qXegMhayFfAd4cHwMT34a0vGfgApEbgioMHlxmawGDWtUfGryE0UqlfpJQAV4/QnSLvm+I+ixn+7do7Hd+Nu97CwE3mpUwMsfoM2JFW2E0RjvMVUUgQr8bjUuFNbv56zOt529XUv9JKACqZ9w8cQZgAsv6leg/48ff2xRZ0h3KKCCg8L8rtlnkF2gD9KygZZImaV6MqCh1fmA3L24tGclY1T/Y38PkTfFSQDzj0DFJ598Yu+o1hTmIHDBwvEF9EP3OTu3iArIHWsDoEI4o0APGBwk47DOaE/1tWx7XFymJweIIkq5hodqVFgqLtON6PWI+cWICpwxMK5gfAb6oI7VMf8mqEDnD6lyraxv5Y/29I6KnzrQgs9LmzA4lZpg0eNWtAafHR0fGf2li7X6lHSnqANIF5IOp/EJqJDhLp6zav8f/zv/gfEfjDYwxDAdOVNASddv5RRV3ZGePFb6RSfpT9EgOj2z/moDFdEAHedeAesVoy091Zc816Gt3096bz8toGLi1d12RgtX5qz2DK7ohOg2TwsT909M2biIElQwmke5T+mx7A5fIfXTqN1s8DPFg3e8eC+fTDcWwW4Yougz5YpdDN8clyIvjGwqXMwLSr6K2vm0BlAho1++3epdjxLPe7jZ/9l4uQSocODHvOYtj7wXlLZCwYxG4DToJS1HvImOBtctr9Fj4/Jad1Zg2e4QWZNQwIDRrcihYogerSnS4+Ds0xmpuyDH7MWcDVTxuqOeAqjwguwQBLFZv2onRzGaPQiFsd3Zgg5xTLFk/3qKKNBAnuQWReGRl6pHIWMv5lFSlZXaCRNd0+8VBESKvodU04hksGgEROYaiIKUwttmOJbxXgekpU00oImRDCrAbKCA18rgO26M9oLS0AfktGHn0uaG3Vktut6LlzNag6ANdAjdC1lf0+qQuz2BaaFkGyBAgYhVRpjKaK99gb4tMmVnlzUMXPdgloDibMD7A+9f5lCKSFlkaHBbBpxh8I6BY1ZrhZ7+WGMW5qYcqPh2k6mrMQdFaAE4AG8gwkH3a4yNfXI8eJ6pqFkbRfqwgBTaChgFo6Pb5KK7uWEf2V3ZZaxFK1iGkRLpGAfaAhU88ykpBSZYX57BQjY4nl+1DHccleNGfJFnVyjF5mnjEwAMPsPdURFkxh/OQyyCzkgWgZlZRqtmjO997TNzAj5hXRf1DbDR+jHe20wbN/76v3559OTRkjPj2TPPKPALQYHf/Ue/kQ2F+QCwA3pgrO/q9ANF3yzAPZdVnSayyOp9iY9W4fLve0Z8eU2M7hSjO0jUeLIk04VmLvJh4bJ2PVVWtNsFdCRWY7+RTu14VHxLNPPvs3dJZ/xDPKMARn5OUcT7aaWDRV4AOOjgCXkKoALpK/CfGzbMwHF6YmGe/9sf/8EYqMAhnejZCOO0KXduTNVBLwWtp/zLCG0eCZZX+3ACVGAu8lC1eZnXonsbCXUPnnjxgo3nIzgh41K+YATwjsqcK65uuKHBAh4nVEYA7OCQ7Cnzgs5gDEE7MG6cnV8OgQoYmOJYRR+Og4Z+S40Qim7zedBbhaSKtwg1bHieMH2HlIrMQQg3F1BxsRyoMEUWoZym4BS6k8cCUAGQ4YIGEgMq3GNF/Ws3PX74iECFpX4iULGBYlaWo32LQIUX01ZEhXJ5W6EuT2vV0g5/w9Dyxo//3OpewMiPGhW5TgaUqROmpuJlhBup/OueW76+iKgQUNGmfpKxBWtFwyOFkvGIARVvmlL12muvpedeeJ4eFP4TebCNqLh185bVqJCny/XrSAF1J3tBR6+a3hxsTWKIeRAfMhbNSUREVMT16kVU4HsZu3qGpIUS1z21amHWyohzOifbTwQqNM+2LyiIL7zwvKVfMaV5AFS0dGR7XP+8D00X5tka96b6jHTm96F4dnOzvQxehPJ4jO3EecRXp2vpBSs13kEebWtvJq1Ab40k/7Y2cHk5tBoVL734cjp4ktKDjx6nW6j38ODd9JWvvJIe3/80vffOT9M3vn47PffCjXR6dpm+9kt/LR2jztHGbnr84FH60z/4PQMqfvPv/d30F2/eTW+981Z6HREVt++kzc0XQuqn45QuC1Ax4t8+b5cIGBTR/uRj1JfbTHfvvpWev/l8evj4YXrxxdvpZ++/n1599VWrUwEQE/L86OCT9P3vv16lzst71NMNaI9p78DD/t2ffpDrKuDcxH8waCNyDmktYJg2o71FRV03kADej0j9BPnJmgyXdqapmDbSMAC0ZOon1He4ZrIQvP/k4CinNgKogvYR0ZH3s6evMyPJBWs44F/kNRYg0UZU6HPsYxkkMDZ53O2gpsa1a0z1h6iOJwcEKhAF4CAGLnsfP36cgYp9gDNI02T5ljk/0EBABeiAMfciKqiTMGUTfkQnfCZQQqmfRF9e4s8TgAr8KCc1PhNQYeAFoiZcrYW+c+/9D6x9i5LwiAqtM+gR0xhhrBiDQBABFQeIqNjYSLueoxtADaLvaEyiY4OACkUp0mh/aedDBVQINELEqHu6tnLQjH5NVF48czYzYMcaGxhzG1ERwYK4x2ScU40KnW3t+ah3WqBC9Inji0BF7FdnB/r89/6tf5J2t5Fzm/UtlAKqPaeqebu3+NIz5irPlTRR0uh4jkRDvvQwtr+uV9TUcWfVOEcG+1Ekwvyo1htvT2/XfqnO4co4u14fIxI2SWMKmSx1Ev9UREMcZzeiYuIiX16Oeymfy+NBdZcrRzK4F3pFm8Eb04+LPhQ94mm1rIMf4rtT2VC+NX4uuEf2vh7pAEOahyXVM12oxZ/LMkspQuWkc3lmKfnkvc/Iczh3BWQiDE6pMO12697PMCTjZwQO9Zba1sNT3GRiutF0yuNcB3PuM5nTXLoHd/AYyVDTF2P3O4IbtnUfx9qZbPE6jXb+WFHiafRMMdZ767p35HsMPP+9joN9RxkGD3w6MPB+BscJGHgtpZENxKNy/T6MtdH6WS0PS2mLdSPdW7HHiAcA+qhv4UAKIlZgSLcDsaQJ5KYl4G9Fh9G2GfZRIwt3s3KXwnrt7u27k5bkphujbazJ7BRKm6j0VTomMHu0y5SG7qSBOhgWJUADOu5miHCULqTzUw4Kdu5tXJjTB+aiuw/qoEGHIChYQDrbE10G9JRjNkNfc9N1aMRWui2MC09sbyHaEkZu1HpA4XZGp+AHQIKKXIN2RvczRj9QMMqeFBjVAT9Fc+uuA/6DnQc6aiw8Tj2A6ZzJC7yM4Xc6QSqKxvnLgBTYHZg+DIZ48AzatjRlAFCVInnD08vlYTJyDG1b5JA5fDIRMR4xnjJ+2c5RL1oHAqfKFmK7thwMKm7eEXboD6lMsfZK5We0vWTBcKyr7A7cn6qdwzRlOnigv8BxBYXnAbQdmgMQs0KwMDtBGRsveN3vFgbwYH7bX/3ba56W3dPk2YfPKPClocCPfvs3XQbJYEFDSv9HBvL223jKht+xF60Iaat695+n55NSX8StJgPgINqgp91oiF0FYFw3g/GpkwFfYb16g4rjbwfWipYejeIhkdGVcojoxK5IN0QhFsypnoMf9+5Z44Y4D0U05eCcnvc4DFHc8fjk2P49QhqD42OLrsDf//s//6OcDoE6RoiowCFrhUw9OgMG6uwJQIO9zuzpRa9MSQYCFtCE0aFEVOApFaS0td5CHmhGYcQLRlTW42VXF2x9r4PWvBACUCEDssAKU34sioB7DQpF9IbPyohvM11rY0TFLFBhxZfcaz1cd2kwZBiyvGjqixQ9J2wtmrQVAirkjZopbGwFXxUoOwg73Ez3P7xfIiqu7abbL71cRVTQU4IeILhDtGm6jK4YQ46ooJHt+PCIKcDMYBXW2MeriArWkLhjoAJqVOTaFCpsipQjHtor5bENXW3XHEDXG3/x5+nWbQIVd155JedMB0Hh+YqIip4xhBdeGswwDwEV3//BD1hM2y86WgspSlCCDQxxzAbGMERU4DIFoOI6UhF5yj0sQwQqbL1CRMXtW7croALKIOgDUCfmcp/bS6B4/F58kvm/kSRZ4sBrOUgnpX7qieaW7kE9XCmnMs/LAy680Sr4bSoqyh/KIBlvosTEmgCo2N/HRUxh67HWEC8REbzMSm4ori1nRyrnpUZFHJ/kSvmskb/hsoKdF0/Vtp1ItPyd33/inaf1hr3opj1ka/Dc0drb34PbOz7nvqLRfXsTYfCn6f7D99Irr3w1HXx6ke5/9HG6deuF9OGD99LXvv71dPjJSfrxn/55+vrXb6cXbj2fLi630le+9mo6sdRPjKj4f//v30u3b2ymv/Ov/T0DKu6+fTf94G+8TqBi43nAzzmiIhbTFl17jNR+V9bgIh0eIP3OWTp4cpTefvsdq3/z4NEDi9xChMV3vvMdS/v0K7/yK+m9936a7rx4M33zm79cPFijKmQebuUDnRUPHjxIH957YPJX9RxUnwIgBi57iKjA+YQz68aN5xLAxgJUbFqh7whUINqDtRJ4GUTbAirwO+oXgLNwFigqDxEVWfY72MBUFryYY6mVykepnxRRgbHZWX/E9EO6sEPG4h1cpHCBu3bjehVRAWpYBOQe0kJdt/ceP3qU5T0u7XZx9/haARWQyZjjKqBCKZswrxaoAC+AN/HdCKiQ934FVCDdlnvOYvyQ/6AdLpSICrE0GQHMhPyQ0wT6BPiEPqVvFKDi0NgDQAUurfCaOzo8pNHBwIZSbyMCFTaGUwJIiqjQOhnQYmB9nWKzPvt9bwcw2s4yNyZo/BGo2ASYonpDHa9j0S0CFVGvkAyR3FQ+dHyevU49R7r2bAtUFE9lRnXjv9/5N/8xC85v7ZiBhZd7zt/Ol2xvqHXiniH1KlrzyJhZ5HRptQUqolydk60rD8OFDwxl9+j9kaznybAWuDKiU9Snc7P2C1NpTH6G1phOnpI8yjkTDs1YOhNjOsWJJ/+M80Y8U4peMzTXN27KZZY20oie+N/jGXS+6dSMrOg/isr3OwhbrNNiGe8Y0CHv4JkRucF61drVQEXdnl81qGO5h7fpyo4LoZi2OSIZCMCIDBr0tN+a/e7e09XakNhDPhvxXwEhbQeXNFmdyBbrITt7TO//Iw7p7VXeHXRn88h46WTOm5DDGjc9/hFdUH40AummRU5p/5S0P/aW8YSnePK6fEwzxGgQZE0wmsI/1Q2vXDNPM+Ue9TFaPN4risMNmc+c53B+Bgc1u8d6Ee//j703YZLsus4DT+17dVVX79VYGgABYSMJUiFaA4qyrZEtyfLYM6OZkUeOsCX9GPHvTMSEF9keDUGKIkEQBIgdbOwN9FbV3bUvWZk58X3fOffe9/K9rO4WaA0iOhlgdVVmvnffXc72nfMdVZ14ABeVlGymDL9P8QM4krCppqcELCDxAXEITIJ0uGi6RBGWQTvErNRMG1Wp6oXALH6vblF1jJqBh27FuJjVzmCxJ7z63o/eJKCYLgHCmLeYA/xUtUFulK09JTkwuAd1/vR92DiqzpAd2dHceYVngA3M7GecQucnJZ26nOX9CEKh95mf/hKoSNsH/T9E84XvSB9HxYQSVLIflMHfDABoz/B39NnqePURYhSj/n2nsGJSCPaUahjSCGJYpCAP6nRUfxSUVphLrBNpsWBvOpAUa89m8bGHnKINn1Nlp27lmG4SJ+3Aa37+uAbGTeCLVTQ6F1E9UcaySv8X+z7sQ9h13OPsMxTUZk7L6xRi9XjUA6BiQNs8+MNXfQb+6t/9di5uiiB9kTVfOtdZRsmgyxKjKajuh9zpMhpMjyLOUvaZaDN6y1zcmpKvZyccuyg9T2hwRT9g0DS4Kfd6j0bqp7Y5ozhMhkCe2ghV1+Y7T3ztSXX9bNvWDbVhRnqTa1YFdHIjbQhkKQTRPgkRB+UTAsGHR6AeEDgBkGJvf98BCwAXB/azN3+ZnPdQVnQmYZC48cvgK5oKU7Fq3BDgZUBQz1p9pvrvYQSU1E+YaARfJsbRnLpLMC0yHGNC6aA7Ck5VXHPM61sswIry78rsUBPquIYAFDV/oiHpmSOpuRyC/25409hzwwKKHFkECFCD6gJBLFFWTNvc3KwtoecBG0iHQtd3oeJoCHiTsET95Mov9guNQg2SY41AAAjmu90O15KVmM5vmZ1KfE9rtL62ZrfXbzHjGGNdPnWKDUaV4ej0FzQeAW+IhzPWvxAmnrWuQBqUM4zMVCLK1BYHhLxhGu6JRtWgkDlz9ixBgC64QxmkAViqgAXGDwMTc84MKucphZGpzJu8zrGPkB1xuaioWDlzVuvm6WjgU0eATvMS6fru5ek0+h4FUPExOdgBVJxcOcl1ppHhhuaEc1ruo6LC4yoQIzCqSJcqBikAACAASURBVP1kI/boY5dsdnFeXLMopaZhqeykcNzCUH7t56+StujxS4+RJoYNGsdGGeRcXb3I4BrWNTJPBrK8is3cFCqIM9HCcuyyKJwpd2r9mpJsOShQnmU5O26g++cxT/xOAUbk36t9iqhB3JmWMRsBiGby5wBK0zlN4IXGiGAu+lTQFg85UMwNz3Av87SWMoDD8EoKH0VlXkp5Nii7ZFzHq/J+rUdFFagoqAJq9IoSl4XM9ACevk8PM92vDk5Fw/sSiElj82xEnNOdrS278tmntrFxxzqH+3bm9KytXlix7d0dW1pasV53zG7d3jSAaGvrN+zs2XPWPRqz11591S6sLtvCwqTNzy7a0sp5O+yPsZk2qqbefvlHrKj47ve+Z29fvmyffPqRPff803Zi6bSZLVi/P229UQipA3TAyTZK3cmrAD6SXWn+RpCJBgd2xNbX1m1iYspu3FhjY2sAfKBiwhmCAwE58/5779m3vv1te/PN1+0bX3/WTiydkD9fgFSSAVE1RylDHY0ze/PmGjP45VyiR8URgQfQPh0eKlNxkpQ+6k9x4sQSqyoQvMaZjvJxyFSCDpMzpEWCg01d6jQaM1GZ0Ovb3u6+dfvKlJ+bm6ccuLm2JgeWQV810lTDRTlNeJ6omgD4D5Cg7FGB9xhYd65gfAdykkAFqAmmpmxmbpaOGnTu4d4B5wljgK5A/wrc687t27QVlE05aTOghGLjU/XZwBwgE3F7e4dzgUpB6EP8Hc+PPRugOsZM0NdfUanGBt3+PBgjABDqIufDhm4NHQj9hPHjmgAIyooKPAv0A3pUxHVkw2Q9kioq2BRy1G7dus1rB/WT5F7Ptnc32Yx0anyS55NABRtiy06ADItgPb6L/4LzG+MjUDE6xr+jGTj5jFFhye96IMsB1RxcUUP10kmOuRr1/VoCFQCIcH1cs6R+CtldAiL4HsAkOtouM7NNoQxCrBV1mAMNuE4EFOr2GO7Nk1PYYeV1MUd/9q//0oEKJIOEzSEeb7n6ejU9b0XQJhE5zF4e+MawYoTKh3MgfJjmHLz+f4+/UG413agVqGjz19qB7GhA3vY8SRangTTPU72SsLzevQR9kw6LgJhX7mebPHojFnegYm9+Ao0r7B7v6VdLLKiOtWUmCgor7ZkIhDffuHndPAirnV8bcqzd4Ddp7zVckOZCAAI+bK5XPeMh3vPmw41bqjIJHhSNHpjFe6VnCp8Qui2olESbgqQ20dIGfU+uplBwPb+KOSwo+mBjR0Pre9j+qQKjYvG7rVq9jvvmWQqVmyn5CPV7t+1xVYP4AnnPB5m8ouyBjoV+wAuyEU2l6bNXIzeqfIi9OuBPI/NfwVUCQW6zw48grRUpkbS/SdHkSVnq05GD12USnFzabG9V7NZ0EH1MZBzoMrM86H3kq4geST6l+kMItFDCXTwj9RQpemCfi5EAdgUz4SIpzumNeDpQlRFxGI7F+yR4JQD0BmwU2W9OieRRbNgssnlE8YXPRhBcdFIYrxIQlESi/RCJHZg/2A4pQJ4WKidPDuzLYl9jGKyQ8EA/6a5wPzQqd7cHezz5jagGQVIJ4iwJdMlrg/GLzkh+et03xCyz+iglb8n3DdBEzAWiYlKSwhh7ObKChJWgeoXvqSbbSrTE+7CrYL+Oj6u3CwEqBvrRd02vzGanilv6iGjoXiAMGH/YCeET4pkxF7BVmQxYyC4+t8ezZCdIXpT0kG19faL6BrY29mT0DMLYaRcXzezxHAqzqrqqtEngB8C2TwCWV4OUwCOf3ynbYpxxth4AFU0S/MHfvtIz8P1//2Jt/B4cT4ZpDYRoysAYyNqIS4JT3puDVe7i1wxDyAWF0FKKwFqGThhb9cA71Uurwdi+MFDAMtKSAEogTdy6Doa0XK0pvp8ev2bp3TXY4RcNAZouU7tZ61qkiW3IKrk356skBUXYW9pFiD+BClZUwBDoEsU/OFJ2HwKgKFlDUANAhX7Xz9fffTs5yGFcyhlXDwIGM4BoO6cjg7WuPKoBoJzpXSqjUFSlQTQ2NuE9KhTAElCBstIj642IU1GlmtoXpKSYqNKHhGEx7MAHeIN7twEV0SAzgIp6UKsEKjAXMEjRUBmBEijkACoiwxSBKwIV3hw8VDkVuxtVnZ4yHCIokIIGDmxVssdSk22sLZqk7tnG5oYd7sPIGiPAox4fkzY67gHoHrKkBVQggDc5hYqKFc65MiblXNBgofEEfvIMVJQGK0wDGlyenRtVD5F9gfVRYy0FHepABaoFuIohZoLzs6t9BQsHQAXehsGiQNRBpSqCRo838YyKCvSoOHX2nGe9YK+adQ4OVerZ4qiBWzzWFz0qtjY3CVQgKxtwDXlQCRKNGIAKZq6Ci9zb2Qio6NlHly/zHo9eumSzJ+Zt1Bvh8RG5P5TdwkCZA2NvvP66Lcwv2GOXLilDBiWozNAdZdAVz4PglyhQRqyfSuUHd3iT6LpnoKI2R65pstGanHstXBmeiPWoz3NUoZQjLgPpyQlLe3pQ/qXnCEqDoqYQ84+9jqoKyIjmdRZQEa9qgB/nd7ASsO6slb/n67QDFcMrKkqgIu49nHYw3b8AKupjkhxWYLHyjFDBkFMwnK1v+7s79sXnn9unn35s25sb9vRTq3b27Enb2Nq28+dWbf/gyNZv3bGlpWW7dWvNzp47b6M2bT/9yd/Z6uqyzc2N28LcCVs5fcH2uqN2ZFO2eeeOvfXyj+zE7Ij9zu/+rr35/vt25crH9tzzzySgomfTlOV9AhXVflClfGmKKCYZbHAWJbtvXEe/nRP23nu/SqAyHCcEYAEAqv9Rl9VJn135xH7rN19gv4VKlmACLJz7mPzGck729vYJSCAIG/1ioDsh35F5ryD+uLL1vT8FxhPNoCOYKyBXzbQnJ6YzUFHQ/uA7oZN2AVT0FNQB4ICfGIecb8gHBMsdKEYzbYCcTn8UTbNL6idWVLiux7XEmTzB60L/wzFE1cTM7IwCGrjW3j5leAAVM15RgUA+AJqgSUC/EtIL2ohNT4H6aZpJEDs7uwNABfQgnqEEKoL6Cc+DucULcxm/43kDqFAgosv5wyt0ZQAB0RsCAEAEb0D7t+bVKHgGBiDKPkoePBO90ZihggavAHIo53oAKjZsbDxTP0GvCKgY96zOBqDCEx3g5MM+QP8P8E7vbKkZOMfpVFQhE1Nz1AK0qDjyLnwAVFCf+BpFdQoz/WirZYCD1/aGqSGn60BFCYgkeeuVhrQFPHgR56AJqIjvxbjChomEh//zX/2F7zuBZKS59CSFYUBFo0yPprrDjL2B9+7Ntm6S+fd0u1/Thyuy0u/R/mRNFfDHDWyY01QAHH8PoKJtBK2UV141wMzdLwmoICDjEWw1+r0HgCEeILKrXS9HsK3p+YYBFfp8CVpE/UAz0DSQpBA++j8gUAGZi+piBhg961mV0fI9AU5S/yBppwRPGozXCJDy7Ceal2rD73KOW3A62u+xmzmTRdC/ukb3C1TgKg0rW/QNwfgjUxv7jL0y3AeA78DKutEROzys2pMcX4FHjfjYKcOjjilA9wSSKXAruztnm9OPcSqtAJsl0xU4jh4G4YNGM+sI+qYn9H+QnmhcwW0sEdgYWAnheiLGgHEgKIx7kh7IfXZWODhN1ASuE/S+sGvQ5Drpv+wvYWwAdESVpWQS2RJqRI+fkXAXAW1cBzYfElioy93eQ3IJ1gCfw9hDj2L/kmKJ1GRdUZaRLSDr05RoGpUC7HPRIDP7uDZoqmBrBeWVelMQyBkbTXSN8qW1V2Ev4H7hX6uSA0mTSqYJPRuAMn3mCigSCaxqWC59rL2vZxZAETRP8WwEE/0545wEkBA2eVTpcnwTAFIAsMFHhs+OyIZsNPU+CZGWgQrG9byKgjIC695HxYbkBhNEfE24duyv1qH9gnXE30B5pUqdLDOzOI7EwmYNQ1sECTr7SGgSiHp0dJhkjOhE5fkS6EnFaS4fvEoIz4C5hM2J52W1EGleQd2lpF6yjjhlVtgwXL8H1E/HGSAP3v+qzUAVqCiC/kkwNhmVpeKsARlpAnJKsGRcGTwvZymMpwik1IGKfP2MatZCXPfmHwgMKYEK3qII5PB6f0+govLM8bzFNY8DLUrF1AZUcJjFww+MuwB2AlZvSwNqCbRq3Qoji5kIkenv1RQwFL2igpRPHQAUAiYAUuC/3T2AFAIq3v7gVxXlFqAAkXbPTCeKftRRuZtnfeQeFdkgjIzkauA9B4dDIQ4DKroGRZ0pEkJZBzVRee1wqJvOeXyO4I0rkaioCOUfDns0047AH08ILRTtfxY5ugEKJYpANAIsyFoJoAKBGSgyBFrYlwEVF/iOU2XROfdsYTSCZda/Zy+Wznk0B4u/lUqv1+/Ywc6Ord9at62tHRkiNsZGpidOLNvE7IR8sV7Pbq2v8z9kSoPqY3nlJIEKZmE6UJGbysmQUgCnmjXSBFSkUlLMjVfdgLMSrzpQgQA8giloHseXO3lHDUAFe4TAEHCgQkZXpspAAO5X779ry96j4jSCquTSFKgGA+jQedCb9kQqSu33bQCoQKYw1od8lWgeLqP5eKBigQEoARwkwXSwQc8a1wNQsbiwYJcedaCi2APY2xcuXOCeQqCU2VmFTKoHbwYodctstCFKrw1gCAlbStnyszgJZVAh3ov1Cecsn5s8iHL/JscxKjFqHmcZ/CoDR0FTRU7byUk7cWJRPLwNGbnMxApuXnegi9EMABUxpjIglALlxfiQLV6+Kp8fSv10b0BFOZ5ynQcCVi5L6udVaVAynCnfPLPu1vpNViOdOTVnF86dspvr63bhwkPUBWvrtxlovnNnnUDF1MSi/e2PfmRnz87bwqIqKk6fuWg7HbPuyDR7FxComDF78Xvfszffe8+uXv2MQMXi0mnrs6Jikpy1BCpqFFaVZ2nLDoZzQCBBNDu31u8w+P/662+Q9g39BRYX5wkirK6u2ltvvWXPPPOMXbt+zebnZ+1rTzxK2RFBgsq8pv3hurQ3YrdvC5CIvhS4J4Lkd+5s2O7ujlMSjRsytELOAyDBmaWT5RzAcO5QUUHgenKGQMoYSs0RdPMqLbzHDPZuT820DRl1AioggwFU4KWgb97nuA/uhzHqPkeUF9A9pPUCddO4qJ8ACtwvUDE7N8drI5AfVRh45tnZaes6gdzM9JzLq30D2IK5wBnBuuizGaiICjzKNgdgcF38O4Ae/I71in5VJVCh4IoC3SVQAWcXARRmq8IBPuywmTa+izFEM23JN1W0ZIrDMa43XlWgousVFWZTE5p7VOrdK1AxMYa+Je1ARVnBEEGUUp6VZ6QEKljZ6P0+mLwxKh7u+G4JXIacxt+wl0NvHwdUxPslUFHqoGjKHfcMOoQAOfD9P/3jf0dubezH6H8VQIXMAPc1arbugJwLoXsffkWzKqxoOX5kUATpZqWeG6JWB95qfYZ7uYh/tula/7BARXMwfdij3WtFhdZDvk5sj+OonxrvX1AdyU51rvO/B1DhB61Sqdd071agokw6rOz9mNfBb1YTEQof/B8QqEA2tnrp5aAoDhJoVWDHK0tdtD/EKaKPW9149Wx67vOGXj2Nc9tyAARAlX0bc0Z/9Tr3B1RoV7bdXO9FXISeoyeS0H9kEL+j4C4BFWVxp1f9sonpSW8E+JAOBPeRV1Yg2Os9FqYmpxiMV0BfN4iG0NI5AiqUZe70SF59XknqKORujkFLz8i2lD4WLz+qKEDhpOpP6A31MEQvAq1J2Ejw0WjHeF8D6RinE2LfC1FAsblzD7TEGLP+FoFl+fMCffBd0Tard0ZUR/CeQTvk68KAMumqFFzWS8H9oKpSD4mo9AtfOKpYvHKmBaiAD82kzp4qEfAx9mqBvekAQuhWVYPoPtHYGr/LztEcpkQkVl+gf0PB9FEAcYhRBOAScxnXlW0h21OglfYEbCakFwJUDHAEH4y+C9DdWFeuJ4Ap+hVOb0XqLTEjsP8FAMoUUiyACqRyur0XFSopxhIggCeH0HYYHbX9vX1+B8mVrFLASYlkrFocrqyWq8sJJoGEXehUU6rwwOJ4DxXSqYqfIHSDrpOBirABwkYjGOtVFeXf6COz2br3PIz+qg+AivrSPPj9qz4D3//3300GWgVdPxaoqAMY9cC+/44Mx0oyZxms99mjog8nggVkLcBGc6C/PpLqmjS9C3FTKgeqqcLgaPhOW5U2P9rw+eOAitaNU4ILPg0VgyLe9z8moCKPAUHULF9lvOk1zOBvm8UcwAxb3l0qp31CUF6Befam6KA3xaFACnBJ7+0JqNjf4++osvjwyqcpy7w0CJjJgPJJb6pknhURwfY6UBFBobpzh98DwAinqwmoGB+btG5fhkkJVIQyCCe4DCqUoEV9CQMEwD2DLiIAixIg8CQeKmTxeTtfZCwRqpAcqAjqKyhuNokrKioQmGEDVVCCLC3ZKLjE2XJDpYQBVBA46YOz042Sgab01R4VPA2kqsCW6VrnYM9u37ptmxtbDABMTc2QJx2c3EcjMMLkeaOi4hYqKpaWGIhZPrXCBqrKjnQqhkT9pCyOMoAR8wlTWFUn4juPwBXX0tlp+HzuIKBHxeXLl0n9dPbcOVYKIKDUcZ7t6OeAvuzItqJzA6MO5bIJUKo2xNa9RO3x/nvv8JnOnTtndaACpej4TBjcZXBFoqFaUYEmuc869RMQJQEE+skmcf0+zwjFIf5z6qePLn+QKipmTizIOIGRQstU+43B7uK0g0oHzbQvPfqoGqLSeM3coAhAXrz4EA1pAGGeRJuM2fQsHMugfIgg/90SWJRBXBquBdihLZQbvDYBFdyXBVVJUEfR33RnDn8bc7+x7uDRYWtw+pquk2Bzd04AVKBXQAlspP1KTD43zQ7Hw4+FWb8oda5QAmVQrAxqx3UlG7PwLwNI0F+V34vIl/7uO6EfjbtzYLGUW9wzZSl+qWLr0TQHKiL4nQAhvxvGy4w3d/S6Rx376MPL1u1s2aMPr9rNtXW7sHqRQMXNtVu2tHTC7mzcsrNnztvszLL95Mc/tsUT47Zyat4QlD59OgMVWxub9ubLP7RFABW/8zv25nvv27Vrn9lzX3/GFhcdqLApJiD0Rw+NSfiFXq7shQawKoMLo6wQBB3T3u4BZ/GXr79hTzzxhF2/fo2VSJubG2xID6DixRdftJdfftmef/5ZO7Wy5Jl4OegYa6FsNfwn2dw57Nr16zdSMDcqKQBCA+THHM/OztjEOH5mOR9ABfZYABWiBAKgME2gAnoWQAV0RR2ogJxAz43+COgHJwhU4DNra2tFxZ2aZMb6Qu8EmNIIVNQqKjA2yJtUUYGxoiJkboY6Ce8jEF+vqGgEKuZmqKMxltmZOQai0WMDc7SwIKACwX/owTr1E76DyotwmqO6AvoSr6Alwu/BCYyxDaN+QmCEYAVsFKfcWwPIg4blMzOa7wIgwhhywsN4qqgQeB9NG1VRQeonABWgrKoAFTq7FeonUCo6NSXGTPtgfII0YZWKCmRK1qifAlio2zKlPEGPipC3oYcxX8rOVfVrjD+uF3IkbJ0SqKC+ToGaCJbkoEK81wZUBIVX3LP8GXbE//ZH/9amJrGWaKgdFRWyMfgsDUCFgpXNxnhr7k6L7d6WdR3XycFwz0ROvkPIi3zhL+vebTQVbe7HvQIekqvtMEbTfdrmKT6bxpAue+/3aH2+lrFq7+pbEXeunIeBoG578DjdOxq98tr3XlHh5l8lmF7q6vozNo6IHKLeaNabxKaHHEJHlQLITiskbeppN79W6qfWsHzqU0d2Hs94Zu+6VOhf7aVR0rUkW8CrQkN+lWAFd5kHmgfm9i62OCsKosygcQOWCVlVe/p+zhHty8Lupd/r9wfIgEQE2vtOadhHICZtqlLWlKwU+UGZ9R9BIWdXjcoC0kkhII6qhXH5aQxce/JUuYqQ1fnMp+iyqJaKfgL5/OMMIiCtagHZ0bJH4CeRuYlOh3pU4D1UbbJfBgPNqJoYtaMO7BDpaXyG+msCOnKSiRX4IOktvak0nwm9KbjBNJqQAdJfSFBTlYWoedT7ET8np0ErpR6aqm6Q/mRAHt/zJszQ2Uigw1hZeYpq1SPIBlSLqBo1gtgChYLiq6C3DSfPVZd0oeYh0fjCLUSVwDieSeukvhMCVkA9hMC6wFSBUiXtIv5NvY8qCK/cjOz/6BlEkMSfX6osXyv0swBEVaBqawpIithKxHSUtAiqUVQOjBOMgL/Kv2POUJXCPhxaT8TrtDZBEywqKiSK9LwfHHuD+PkgCIW1deAlaN4SWODngvvIKdNEpaVYWrhU2bdq1jDYP7A3cA3sN+yL/b3d1KOCMR8HclRtFFkL2nB6pEwtpnUAlWUAY/L1BaBpPhkLcEo0AmcPgIo29f/g71/VGfj+n/+OD70tUD349ypnW/H+kFh3YzC/bdJopZcht/uZ3SGUUOzOrPAanTgHSfhvpGTm3JqBf1dHIiGZ6yfzuIcbHs0Tpb/W3xvNvOHU8SUg0RwiLIOlAzPX5gGVVrp/iULdjcAwUhOYBeMAAIVnaaJkEgIU1RRwKgFUICAVYAUAC4IV+3v20ZXPKsMqA17IFEeGBh1+p34CUBFVCgnxrzVMkp4MYS+DsQQrmoCKsVHw9h8xuAXlHYHUMIpkYIEWajxlQNYd7vJBotoirgM6hihLxfWZUUDe8FhSZKUoQA5lE0FY0AXRiPJGU8zc7BwxmxTzjAxS9DpAFmo0HEUAzVDSCjDCG57RMfe5Y4mmByzyfeKZq9yUCVThQRBQAQBif/+QlRSTkzMKSKKcGEEkn/v1mzdt7eaanST10xQbWyN4E7QXyohBOW+HBjWDPlHKW/FeFYAn32y3yz2kEkc3tIuKE9wb/PXvv/++rZw6ZecvnLfTZ06LnskrKbCnmBF6oIA85hMZGQxce9lwZK+XewiPj/V57523bXl5yc6fP2+nzpzzzB3xjHY7RxWgonreqg72hx9+yMzw555/3pZXlt3gzqWkoO5IFRWO3aYeFZc/4JyA+ml6Yc7GYSh7lgnWGPsjMjUiSwxAxYnFEwQqWA7uQEWMEeM/d/Yc1xRZJTSYQxvUA1Gk48pcmuUZQRO58nvlHNRlUfpeeEwt362HJkqHIRxQAX6RsShRzDEOiYSA3Yqfk8CoBvtD8JfUT/4wCwvoU4Gs/RzA5bn1JnKp3wg9qFKGi/qpDgjEHJXBkHoQog9wMWSx8w+n34dUVFR0Zz9omsomdM3gBx+/TYfjzZTClGVtTJnykPRSRQV4o49sZ2vD+t09m52Zsk8/+8wuPXbJdvcO7PqN66SIu31n3S6uPmxzM8v28k9/aqNjB7Z6cYUB9zNnHratg551RyZta3PL3vjJS7Y8N2Yv/s537Y333rNrV6/Ys88/bYsn1KOi159iv6EmoKLck/XgXbk2cuZHWWEwPTXLptnoUYGKCmT7o2cC9g90HeQwKipeffVVe/HFf2RTU3Ae6iCFZigcV2Z8EgjZtrWb66JGcrqha9euJUAAwVY0zh4bRcb/NAEFVg3MzVI/4jsAznAtVQoYG2YDfGdlA+SDOzEYAavxnOZuf+/QeiNjdNgR3McLQEVQEY6NqWIjzjuC6pCD+C8y6wEMhDMLWY9S97KiogQq8DmA2tFsmhUK+wfUITg/7LUEXt9Oh9WCuA/+LRB+ynojysoDUAEwBj0Y9g86PI/on4R1AZhTVlTEuWK/Dne0o4IielTgd9w/qJ8iIA+QCq/QTRgL5i56VAAEohOM6rf9A7vlIE8AFawKLYLyDJqPARia5FgxttRMmxQAXdvZQ4+KUZtCxUJfFRW7OzuJ9xr2ZIwD64GxxPoE9dMkKMImp2xne0cZqEWPiqpeOv63kSIrMjIjMV+ifspNWemU+/zGOYogBACfoHKIoEKS0UWPClFDSnpEsIRJKz6H+G5UVJT2Vzx/zO+f/OG/1RqNTwoccnuDtmQhlYfaxyHDeGybo5PHBdqHzW4TeH78amSpf6/3Fke4qDjymdbvba/QqVWZ2TIX9wFU3M3zlnrRtcrA19RbKGcJlwlZg98PRTp4NQYRK0ST+VYRpIJNUWaua6/HvSMAXPQ6KkbLeS8qNTL+4rqiZULoTRZ+WeX30DS8RL6Omgg7lVraLN6XIX/UA3wK7jH4W9h74TuFn1Am4eBvAfAySObnnxQ5ngAU+yzo4EYKuyHv5LZd0GfiWNgwAS6SK5+Z8wquIpEp5iYDgBFULJsR1++jZrZcvzjrHmDFr6nqLCq9SW0MGpt2wyhMvgRI4nmLZ66cnPSLe/sepsA6RHIYM9ujN0BRmUf7Hv6cN2VmpRvPtYNr9PX6DNJXX5grJQggiA67jFUo7PnoWeANy8H1YwW+AAIG8f258BgMgtNngD81aXsHu55s5XGVlCUu8CD6FYyNyk4iNdP4RPKf1HvE+3cddZgMB7ACVI8IXuO50D8M/rEoIA+oe6JXVsXuLWIB7NdlfSY4oDpV1EG58hVBjrzPRMcbCR4M5nt1SmrczYodgSRqlI3qCFFTseKQz6AgN8aOeZyadpuK4IPugfdRiQJfVHEG0UDh3gjU43oAWg4dNNBR98RR93UQY8D9pO9UtZISOqPZPW0Zva/M/OiXhnM/Kl8eNm0tMSr0H2hF8TzQp/TJ++oDhu/hObgPsZfCZnIwh3OBf6NKgsEHjAPVEg6QjJrt7GhNWJXi84i1wL4QkKXebaH3OWeHHUP1KOwefAh7Af3RAPrwb24rhc2rShiBTNWkXf2O/R39T7WflJChqlzV1suGd7aLYm8FGIIxkg6UFSBZ3kaFhZhPBLhgPzAm4vfVuoExA3saFGLoIzmRQKroj8ZYG9kXcBaVFEYQCXJBaJPyrR8AFXdjYjz4zFdpBv7qz793zHDbFXQlY2FYgKOkVfo1Tc6gGT1sQDjQpaHun6U2rQaZYriDzk0dCMkAh77TbNgPWWKwxQAAIABJREFUffw6iOBp1am0sAZiDOSeJMur+S7VDJPqZ8rMjBxDzJkFVL4IRrEhl1D+ACmIxpM+p8NqClZU7KuaYndv139GdcWeffLF55Wbl0AFHoFOPZohxlJEsN0FdQ5OVrOBS8c2DM5wnqtAhRQBKyq6R9YbVQa/7ABvylRbixKsCAO+7gyVQEWAFeQfR9YBm3qNpFLVUYJlAirCOKFzzqZaWsiUcY4eBMjimJgcACpI9zEzRbolNdNWJQWBESjZAHm8oiLGHj/D9ikbnuFv+X3QhRzaxp0NGhjIjB0fU9ULAno9pC67Q9QGVCgQUfSoOIQhrkwcgRjDqZ/KZtqyd+RYhTkeQAWynM9dOM+KCvRwoOEP44FGSt/29o/I5c3sEhhCXvmiAJ4MvrKxFuYBe/m9t98aACqMzbAAVKiiIjtN9XOf5cxHH33E4OZzzz3HZtq4BA0PbzhI6icEZZAhnZnw+BlWVJgJqFicFxe+c34KqFB5Mz7En31jc2JQgqGZNg0vgHI1uYT9g0oR7LvDA10j1iOc18gSLmVgCVqUQMWAW9hUieFyrC4xS/k0AFREKXUhnusyOX5vcow5rhDZxZgqZzhw5jBnXfzhuggWq6F2lZtd95QBW6/i0lzkHhVlQDzmqbx/vJ/fq/Zqqnx2SEVFZQ0agIr6GpXXLZumD+i8hoBDzKsS3LT3AVQw2836trO1ab2jfZuZmrQrn1+xiw89RN1wLYCK2+t28aKAitdff932dtfsoUfOsEfF8slztg3qJ5u0rY0te/0nP7BlNNNGRcX779vVq1fs+W88YwuLp8z6AirQTLs/cqiEgzYVzCDFIFijAA2aIPbYPHtxYclee+11m5lB82oBPnCcENwHqHD69OkUwP/GN563UdoUTUCFHK7YD5A3oJUC9VMEn69fv243btxIS4N7oqJifGyEAXgAFdBZ+DebQhKoUGUAqJ6wz1DphoABgrqkfnIAHJ/FOU9Axf6h9UfGqWPxLHhuBNCzbsgVFdgDcPiilw2ugevH9SC/MS78LYAKVXugim6UsoyNsR2ogE5idQaDD5L/ACmCXgpARdxLlSRB/WQEKgDgIOAAvm1Ul4CyDxUVdaAigmslUBEBtqDOKoGKGC+CRGVFBZ4/AwRopj2u3g9F76i1GzfVa2NKCRYlUBFBe2X954qKQaBiq9KjAs3G24AKgBEIfKTgflFRAXoL9EFicAWNTvFf4VgPtT+LN0e9Waj6SmkOMH/RoyJgSTwvq/XCifakBfwd8xhBpJAxpd7ItpkncKDnEwI0TrlR2nOwo0p9VF4ngIr/9Q//zKa9ooKBLc6504XcI1AhOfbrBSqG2ePt63RvY4qAWdi2fC4HLprukWzx2rO3Bv7lDdzttrrrz1Xv1+zLKWhac3pch7cCMf7x8opy+1qSvggkwu+pARU5vXggQartIev3TJ8bgj6l4GQEHYvPZozC9S59tPyCHBaYoIzrpldpc2Q/TMFMBc4jEUTJXPT7XL6HH8h7eDZ7BHjhH5DGRRHq5nu3/LUE1eofEfWTgovwWVK2c2jXqKalHdu8EqiYrOyaEqhwACp49TU/qnBvnL/IeC8qT1QlXXy6XLNaQmBcFT5iyFr6Yh6IjgQ9ndsRJVh5VrYohdTQGuNTXwZUmDSPtdcDqKyqA7wi8YuUQA1rFHsj7Fr6R35tggxF42hQ/SLIWuaYpgoc0j1pPzCb3pMCmSjm7A+RxR6BZq6txwJQwYhEiKiiCb5+jA8Vlriv9nm5xzUHqSrEN8rszCyvFVUUMa+xvqxEQd8CBx4IwmMLe1VGio14pYr8JfmX4TtFUDv0mKpcNOcIaCNYr4oe/x0VKd4MXnI6+9+4JimmhFJWEqu0Hl5RErRNTHiUPmWPCMRmOurzoIC7+7gJVYt9yprwLJKKfwdQI3BJtGpBOcU1ROXGxATtA4xXQX4AG95HwpG0o86hkidYcaqfsF1hN+F2UWETuj35S4lOS5Rbva5kEUAy3stpljB6LbPOrPaDgK/s2kWsT8+KWWHViydbRFJG9FQJYEO+gaqidXYA0h151YroQGHrBHBR7gckEZb2SgAjIW/DfgK1MJOOuEZOczcqFoioNqE9gznwag/MG6i0JJ4ccH4AVNy1nfHgg1+RGbhfoOLuQQoe61/vbDRaJApUyCSpK25IWjVoTC+vpNDvg4q+DajIor3hHkPBm/qUNJlCUc4QF7qXCzYZh3fxfX7Ee1CEskrzKzSfcwraHBpGyhZFNjZon9DciRUV+/u2EyDFroMV+/i5b59d+6Ly8CVQAU2jckkh/Qz+14CKCBqVgb9QBBFkjayC7AyXzbRHGewBeMHSzZFQarkUNQyYTAMFh1xBmQiu11ewDlTQyOh1DQ03mSnoxqdoprQvg/c7Ahp0/CfUCBZABZWtAxVwvpHNUFZUMMN2epoUP2UzbZZ3wnx1eqOoqMD16sFWKPLgrCyBDB0F0Hod2ubmFtcaRuP4qIJQfNvpi/CsbUAFgksy/L2ZNoAK9gVRhgZfZWa9J6ghWwAB+GimHUczMuJZcdLvp4oKUD+dv3AhARWpJweCdr2+7R+i+kFARVA/0dhwoKIeRMHv2MvvlkDF2XPioWSjRGSHqKLCazYbMhWHABVkelKWFLNnKkBFPqsAJD76oAAqFuZtfHLcKyp0PkqgQj503179+c9t6cQJ+9rjTzDzAtnHZVBBjt6InTx5kkAXsoNj38dPGby5qquco8gSHNKDuyJNq85hg1aoyfGqr9dQ0aFB5mPoQFMrUIFtBgeXjkNDgzp3WGXOe7m593tBgBJARQowFhmIdEy8B0GiTEgB61xRoW1edTbqAaD8fXw600nVZQ3kVl7LqmPMPRVfSLyL7YGK8toVZ6XmvJYNacvv4F7xPQb3UoPJvu3v7Zh1D5l99/kXn9vq6kXb29+xq06jhB4VFy8+YnOzJ+29d9+1G9c/skcunbOV5VM2t3DK9o7QTHvStje37LUf/40tz4/Zd7/3PXsLQMW1z+zr33jOFhZOWa8/bz30qGCDnkPzZhXNdgdAW05QgEw5wxKZh3t7BwaKtrnZBfvbv/1be+KJJw1AAgLje3s7BP/QbwaA4+u/fN2efeYZO3/+rI0SYG4CKqoVFZAp16/dtO3tHVUhHhzaF198bmtr6zyPcFhQLaDs8FFWViC7EPISAEEAFaruGCVNFU4Tmz1HRQV7CYgiA/cA8AE5R6Bh74AVFdAnUYWAYH/oIDNl+FEXAACZnnJApmNH3Q7lBCsqnOIJwRMEkgOowB4OaqOoGAmggjQUnQ57O0RFBZ4T90CQGuMIqj8CFbMz1jPR2s1Mz6qiYnePc4Y5gpN2LFBB+gdVnuCZME9RGYLfCfZ7hQJ0DQLsSe4heI4KwG6PHMYK1IuiD3ODZ7lx/Qb5r/leAVSErIxAOhYk5pnZhp4tC9mxu79dASoOdvdbgQpWoPh4MY6o2pye0BhQtQcgnhXCDlTU5c6A9VmTvQjPROAswJoAKsybpOIamD9RSmhv8W8ACEZG3GYQFUIEccLWCzstggRhTwT1U2SIRtUbAhrlfJbXESAxan/yB3/GoAcSOphMUQcq/BkrtvyQIHGrtXxPgddipl0oV5KCmiXUkL/eD1ChxqA58/zublrXTc1gRTzNlwtW3BVQ4QkZXh5Znej6GhVz3+CpJd74wZnxfmWFG5nHlgGCum5vmivuOx9XZbbuAqio+EiNYEX0yYqGwwpcKyCaufMHnq9IEirPJGWT9wtMzwbd1pPfV55pvI+zFtVQ5e/Jc435J4NBUQNSuudpjbLdE8+tRCrp6fBRAqjQ+PRkMcWSN837HECFPusfCHADYGskWzhtVxk0rV9NGIzb7zWgomIrFdUbBL0ahsVkn6j0JbVV1U5FMBb3U/a7+nBgbLJlqyGLtucegV73hB8kEEQmfRvOmHxpr67T/pWPHLcM/xgVGmxiHs2V5ex60pSqDxho5xpyxag/O0cCxBiYJTuD6H5YLeULC7omVW+qHwMmCva4QA2Ym1rrbDuXPoGxwbZiFJozJk5MTqb9Sns/emYEqOK0SNhHuHeAQXEW5FuKTqh7pH5WGks0YlbPh9BNqqiVvYmxQmdzPkH5hIoK35Pq6STwH++rmkD5s5y3mvwQMKCKBpxLBLRTVZBTGOFrSsBTVY1YKQRm4MWzhX0JAMXTrvwf6fey+Xz6nu89rBTGqx4XueKc/ShJba0m2AQuHaSKTQv7jQmY0U/SK8+iegh0mBHHY9UCE4by+cXzAqiKKmOFrlT9IRomNXTX3uOp1+krBAZiVqq+EAga+yiqtnKvonzQVMkkWjXNofpypKQQp8nVeROwEToB9hKqNmKuArjAPB0eHtgIabJHuV+xz8N2gn1M2QfZ4IAf7o096A+lzz4AKpoF/4O/fnVn4Pt/0VRRUQj6YVwQdxH3DhT31zpD9wNUMKO9MBeHAhVlz4d4EhegFHiOkJcPybfvxXjPtCrpMjH36flaJjz9uSaE65M+bL1iqMGrGnyb4dyFAqsAFWqUBSHNgAvoIUD9dHjAwMWO96jYIVCxS+Bib2/fPr9+vTYyzaEEvQS6ZL6aGoVhE0h5VrA5izkCC6WxHdkoygCYYIAiUHYoJpRaMsuj4O1XwD64CaXYS6c4MggjA7N0elOQH8EBzp/Gp6ZbMtACmQdQUQYAMCHh4OM9BjdYWioACwF2Zp2MjtnGnTukfpqbm7eZOVRUzNgJUgmhogLhEJUf6qcUGYIhMUcBVsQiCKjI1ADV9wG2gNd8h4ZhplPwTAU9Kg00cHUH9RPm+mTqUTGpEmJUVbDMUeWZMDJgZCnrocho87mJ8lzQYDBbwXlpcW71fBo3+OvfffddO3X6tJ1fvcBMZxi3dDLY60IGeqfbZRNWrAFLK70JNXo9IIivNZHhEUYFgjPvvl2lfmK5JWYX1FeoIEIJcnCEVpxIOVdx7D768ENDP41vfOMbtrJykr17UqaOB33wO3pUMCvKnTo84wfv/4rP89jjj9v0HLjaUcKtclMY+GVWCZ4VT/Gzn71CoOLJr31N5cRoYub9MLgfme0vxw/rMDs9YYsnTvD5WdnDKhgHKpx3nXsjeVS+gyrZeg4CxGcqThQ7MfpZz5yrTc6gbPLC+ywkhnZ3pnoqgWXOdXI23fAu1gRnvYwL6N6FAcvzo9+5J6Mx/ehIot+RU6Jry3eLTJtMOZeHW6V+ymcu64Z4zrafYYSWzT1LWqi6mI+MRP09hQqyWomAQL2RZDF3/KcD0sfpbum5eB4003aXoH9kW1t3rNtBBv603bh53c6cv8Bg/9UvrtrJpSW7s7Fmqw89YjMzK/b5lS/s8juv2ZNfW7Wl08sEKvY7E3bUn6C8e/Xv/saWZvr2T/7pP7E33n7Hrt+8Yl//5gs2v3jGur0p6/UBelLi+d5pUniSy2lvcejKRMXeQDPtDYKyoIk7sp+/8nP75te/YZc/uGxnzp613d1tOrlrN2/YU089aa+88jP7vd/7PZudmXEecl+tAMN88lBRIUcTAdxNu379JgEROGroo/DZZ58yuwz7cW5uxhYWFxj8npwcI0BCmqMjVFGg549XVMzM8PNbm9s8ywQqWFFxkPoZseqr17OZaVRU9Bh0B90AHeSxcQcwehyTzjqacAvghkzDSUOAXkkIHQdW9knph2sBuIYsAiCBTMWgL8Ac4RWgAwAHVONBp7F/06HkOQAsBJcBQEA+3bl9u6B+8ooKVqOMsG8JgYq9XTs42EvVICVQAVnJ8nrfgwAdAgzHGHHPqKgIOqGoUlFg4IhzAbkKOY9XgNlB/URn2bNsIf9v3rjptFBwML2qkUEIZaCKxkh2DZIM8BPXkvxQQDFRP02KLgFUfPs7u/ouAwjg2D7gukRPjQgWwoHH2gLgwpqiogL3ppzyqsISqKgHUUP+xjnnPqBQlCMOnR16TgkeCpbF+FWth4BdpuHhvtzSOSrtp/LfEVApqZ9i7cK+YuWKGcGjsEvCzopx43eM6X/55/+G+yOACqyf7BWnfmoCKmoyr5R1reby/QIVEqq/plfzhWOtNe+5sXNbhn11cLpmXS/VP+Of+lKf626AirYb8rv3ClSUvmDtwgyEhpvncyjtmANmye+o3Le9/0k5vmFborp+US3bstY+bu53JK8w09bttzYwpJ4c4pnDPNsNQAXOU5xRceCPp8+VQIWCcZ20f+IshTmYnqC0D/nHnH2eDRaAMLIx8AMBa7wCqJAMVQA41qEJKIrrJYvcA+8KnnuVtoOqCJiTYsmD2G2yIKizIkOeTwD6pZofEfdOSTL1PeY3kB+mjHXRPMHGL32STG8FmRfBfVwusq1z4LJ6k15XOol0QgeqjsNLfREG91Ta06iu8UriqNKJwHwAO1m/+Jx5TCSqAEinRJ+i7HMC3wMgggCiWDMAKNE/IfYQxonqCVyPVRLeNFygjSisSl+8nG/1oARbAWyhLhO8CA6Enep6OJ7BzTTPmpfNA+A/mhYHVZrmH2wJom3CS70U5BhEol3oLfYsYDWsgI+yRwTtT0/61GcUW5FNNkKbLL8CxJGvg2x+gES4HhNEvHk6Yw2eRYYxoFI4aIdgh0ZgnZ9jBUL4S7pTgqDZvFy+pp4TskW9YQC4TE5M2d7eLu1SfIafZUKkepewV0r0O3HQJIAJ+uLjE7T94gzqPGd6KlFBCbgJG41JE+PonSYAKxIdMAcYnyo84NNHX5NI1KrGyLBGAO1gOwUQQI8uKM5c7ig+5VTZrHIRaBB9RWJtyxMXciUo8dh3o9ulPZ3orCDLeM61jrShoo8dADICFgC11JQ9bFLMlWwzgdDoQSqWiwfUT1+qIfLgYv//mIH7BirqwXEXbYNPJQP5nl5tKQHDjK2BWwyhfggj866AihyQqj5DIL3x1wJo4PjvtsVsedWmrNfywaoPWRrKuoobMUMoOprXQU6p0iRKns+yuW3U5uUAFpQbkhoQNEPwGUGJACpQORG0T3Wg4osaUFEqqHqeddX4yAGxUGb1AHsYV3jOoLqA0hkdE69zlPjB2WeTUGQBOFBBpeAZB6oAqFZYxNxFJUDwKAcvIR1m59lUNrSyDEX1qcAvnlXZh1LMwcddGsrSNyrzDbAChgiUFAJpyJjcAVAxO2czc7M2OTttJ1ZW2LSKBquXd1KRpUALlJ030/aqingeGio1oCIHL6SUEUSLJk5htHLMwcnY69nNGzcSUIEsVQIVDJ5N4MYM4gRQgXGV1E9lJjkCv3KStN8P9/YZ2AqjLbz9ACqQbf3OO+/YyunTduHiKoGKMMIjiAHMD8YA9iTECIwqlI7iugSSjg6So1OeEazPO28FUHHBzpw770EaVBmo4VsEwOQg183JMNzNPrz8gd1Zv2UvvPCCrZxaUeNfn/sABJjp60AFLhXPePm99/n8jwOoKOhf4hzQgXDjEvt5fGSUTX5RafOUAxUINJKj1J0hGWbKhLl9a83OnF6yRx552OU15EBudo77BHhWT1ULp4zGbSGjy7MY57h0vKPJa/09XIeOi09lBOSypDVjjk6tGXe8n6ugBvUOHLvyOmXgLP3d913d2QVNDoKa9YoqZZEpoybWM92EIGA0fiv2RtnAuqHKon7vMtCY57l0LvOzKhDfpn9yU7vjdPJQZ78ekAF1BoH1cQIVBHv7HdvcvGVHnX3S063fWrdT587ZPqifvrhqp04s2ebWup2/+JBNTq/Y7fUte/3lH9nTT67a0tkTNr1w0rpHc9axCdve3rKf//i/2eJUz37/93/PXn/zTVu79bk9941v29ziWet2J4z9JbAzUEVW9PeoPycakSvoEamU4nDGuel0+3YDtE9z80aqtjsbduHsOfvi6lVbOrnE4A+5+tHkembG1m5et+985x/Z5CSCtYPgU5KxnlEHBwW9KW7dQkBeTjAC7Z9++qky90ZHbXFxzhZPoKJCQMXy0gmbn19kFQGqCgIMmJ6ZJiS5vbVNmYaqCQAVqDiYmJxi1ZpK9HvstwEZcXAAeYfMNoHhoEKAHETFXJz36Ns17jSCE1OTtnd4QK5kJSQcUK4HrQ/0KObkYG+fcpeOvQPFkI34HZV/AI8j8zaAZ+g4ARWoqKj2qMBZQ48KZVGi8mFOzcL3dwhUzM/PULcSqJjx6gsHKmgNebA8zmsJVJQVFbhPBMYxhgBtAuAg/7pXiURFZZwNXJP9TLwhN3VcIZcisQFjwDVwbfycnnJeZm+yubO7SQ5ugD6s/oD9tLNLIIfOaL9HoAJ9jABg4b9oJIr1wxwp+WKcAAHuQR1YAyrqcqQuQ+P3kN1lkAX3j0bVpV0W1AVx7bhGCVSU1y3lNMYZQAU+E/QR9cpVXKsEKmjnFNWhuMb//M/+tBWoiP0wIOMlTBtFoQDxwffuF2tI8vR+LzBUYLdfNOP9svM1jrvxyaryrFUftAT5h+mPe9M9dzPWqu3RCggVwckkm7k52oL/btOV1E8RNC+AirSni4z5yhULSs1sG9wFxFNL1pCNWVy58JV5Jv092E9MXqk1sR8270HVE75AeVbibIctFlm9DNZ6YLIEJePvdZvwuHXnShf9P7KsiAqJ3J8iBasLuzPk1vC9570lnXGBz8Yb6VxU51h/awqCa6gKKIffTM//OKAibby8jlGRGn5QgMFITsArgpha/jKZTsHK2O/YAjk7vTrbR4eosPHgJitToJNAH8UDMLA0pW8R9j90DgOmDg7FlxBoFqAiAE/V1mFrCugIUKdSUUbwwAPyXlUhgFwJFhgXgAvQhQKA5trwGbvUhXjW8OnzM1TPMqpVohcHMtTxOVRCli9KxugD58F2PAN6fTH4DtDP56hco5xZL73PSmcATQQqRqnD8XckduA8giILNMOYA8YlPOaQn0H9JFSdoMqHyLinXSZFls45fLoA7rAHGMgOMMeT0hBMR3Ac0xlVj3wGn6bovcAxZOGU/h0MBLh5AFVcF/YoQb8T2OfbbtMoEYV7FgAF7uP5aQDdsF6wXWQrQ0Z1ubcpc9goPcCSoPISOMn9g7ntiY4Z64iqSdhf7N0ZfUeYZBqfl67TPZy5oaGiglRi3pMi1gGjqPiKyaYTFVfIA/qarCoFPVmmgE4+rTLdlD7lCYXYAyEXCSBhvlwlS4Znain8jn2jpu86q0FLJ4kVvZKKSpYHFRXHqZkH73/VZuD7f/G7xwy5rsDuA3i410lpASrajA8e7vsBKhpt05bna7p+tm1y0534XKKduvuHb+bBHAJUuNKW7orG3u2OVz3AWBlZYRA7bFEJOtL4KDJQIExpDHujJQQ9Dw73mXWJUrwSqNje3WHwhBUV+3t29Xrm4g6BnR3mKlhTNRCl3AI9j4y8CExGQCIMWGZuMsiAoMwkKZLiuwFUMFuyUlGhbI0YTxlAL5VLzDk+R4cZjTBB1eEBGlAmQUmTWgq6mopOnMnKSBAdVARywgDgMpJaWgYHAznjyjpBX4LOUb8KVMzPkv97EKgYJchBBUlqI2Sw+liPASrimcLoB6iCAAvGGxmVCaxwoxTP2gRUALAgUEFuRSAwMC5VzhqUGGEQJ/vdG3+rmqZvRweHzADinBMY0cGlWdzvkxZGQMUpu7C6aqfPnFHFhDek475AuSSyUmM/kGOyx+AfwaSOgIp0lnwwCJy8/eabbPy7urpqZ85dKIAKNfbCfpchlSnEJBo8YOwG40cffJiBipUV62OJg/s0KioAXqEs1PNZwCaD615+/1c0fglUgP4FxpmXD9MYY2MxnUkCbzZir/zsZ6yoeOprT4p3FU1hnUscxx1jR2AT1/ns049s9cJpe/rpp5ntoWyeDFTI8BQVW6x9rFfp45dARKxrnKV6IIsNmIss11K+B1BRfjfdT+HoY4GK+lrWJXF9rPg9y6Hqp7EGON/IbC8zgPUpHPDgS/a1SJsZzlpuph0ypP4zxlL/mS5zDGVUOdrjgIqcWTs8Ynb/QAXuAPl3aNeuXbHtrTt26syK3Vxft0cee4ygw7UvviBQsb1z286tPmQT0yu2v92xv/2b/2RPPnbOTl9csYnZJRsZWbTOyKSh18ArP/ovtjDZTUDFrTtX7dnnv2VzC2dZdcESJex8NI7sRzl0bdW9NFxAjgNIpGiWfNjbP7Qb67ds5eRJ+7sf/9gefeRR27h1W3pjTJQD6Ofw0MUL9vmVK3Zx9bw9/PDD4swuQcpa8JN5hH1jReH1azdsa2tHVRudjl29epVNu3ENOJ0AKU6cWGSQfmpyjP8GUIFKiQAq8D1UKWDcoJDCtUEPhUA5qhnHJyYdqEAgCYFxVVQEUAH1EkDF4WFXVQSj4NodV7UAwFyvqICzDqACPNrS88hAk/yBnMV/uCcq39qBijnqL5wvfC9kFz4PnRLAR/SoADAPcAN/J7AyAmBowSYnQf20bQeHewR00FwTQAVARPbN6HVFQeEUIQhw3y9QEd+LHhWpmbb3VcLOwr5Eb5Gg5AqgImRPCVRgvRNQUdgieL6d3S0bHx/hXKDCj1Rau3uSNWSC7JFicHJsnHMMZz8CC9BjoZvxeQQNZC9MMhMzUxjkLMXSfinlZCn/Yg7xDOw/5s2060BtCVSU1x1WUUGp6bqoBCoigzaSQCIwWq+ooP6vARX/+vf/DSkgkHnLHmdsICp9VdcFKZCQMibr2mFYKP/+kYaKTL3/ywwOtuUvSraR3axnLsGKpi/VHR0P4db50YuvtueVtQX/jx/+vYIcdw0CfRlABZO6nMYm0ap4ANl/L8cfs5Bcw1I3FAkZ9VlR8NS/XfSoqMxN2E/+ZQbXikpJ8voHvcvAtOcs9kjMwrVhe4mKx/vPxQLH3HmlBe4VDXx5TmH/eg8EBti8X0Jjtv4QoIzUUMW5FHAgGsOI6NGvIk1PtQI6fJbhtgutr4z3FOGDAGnCxi1/H7AfvT8F7caiyphy05PS2mzOdDIKYCmHDryyu+x74MGrb9GwAAAgAElEQVRp2tRBR1SAUJpjJXcpq7zhhaZ4SFxDI2Q2OlZT3mGvqJITEOMUOuxJkqm+cE8Ee+GrRnA3zYcH/ymB/Fkpj0mLDD/bqxMjW92TqOi7eRBflQwaJQARZrE77ST8s6iQjLGm/RZ4LCmHFRDGdYM6U76Xrhuxf9qFvt8RoEcQnb6T9zZk36fipWdyerjUMyJXjfO+YAMYgz8+xn6dPCNeYRKVRwykM54zwuQ5+MwYRgTFSZuUguWljPZ1d0olgQ75oQQAKJguxCCALuhP9a4JPZyerZBJvFKc+0jgSgCdmrPDX2VShLNG4JqkvfIqUjWj17wh2QHzr2qloKcL+i7FJ/KZQ++OTBeFvxP8oD+tKhzIKdKpBWWTh8Ewb7DVxfihGirNis+dP1OSzU6Ph32tag2/T7E/8G2ePQKz3gPE/XcBHQKXSj+Soou9SOSPRGwlwN2gzEq+se8lyl8mLqkRfNhYEXcDYpPH7oBF9LZ5AFQcb2A8+MRXawa+/5d1oKIQgjwJTUBF8Yw1I+a+n764Tpv9Xg1aH3enwQyByjcGMmgcyfVE1Gx8R/SyUfMXfywUmMPz2UCtjqWSURBXaBxuO0hB/VEuQ2jboVZHy8y2eRqlQg5kODXThqKQImVlBSoqHKjYP9jP1E+7u4aKCoIVTv10tWgaKj1YBgiHAxXCY6TQovohDKAoRw0HG8oBShT9M8bHpxjgDce3DlSUIEcbUFEaWjHmOB4YE5S1AvPIrlCQWsaRstEB6uD+vBfLRA+dxgIUIDKiZIgeqdEp6DVQSurLBh7vbq9WUdECVOA6Qd0hBSpDJwLNYTjE/JdZVGUAAM+AcSKAhDGqQkIcinQKhgAVAA4qQIVTV4mfU9yc5bzHdmOGOpuBywAsgQr5A1WgYmdr295++207deYMqZ/QTDuAiggUAahAZo36qsjgIVCxr7kHUBHOPA1CP08Izrz1xht2EkDFxYsCKpj1QQJ4GqHY7+GYpZ4bfBiVbgOpgtH70Ycf2e21dVZUoJ8GLiEqJue7dGAmqFlg4CSgwisqnnjiidaKCtG8dBlwxdr/7OWX7cTiCXv6qacqQAWdUfqzAMyUjfvxxx/Y+bMn7VsvfIslwuJKLamfRMMW+7fcP5UIrS9iHeirBoY848Wd/SYwQqGVAPgyb2hoJJ0gbwhYk3kBLsZ1h+mNqlHppmxDpUZkKC8tLVXKxnXrKlBRATchLwugIgzSSiBjSHVF+Wj177S/N7yiImUN1ipg6qqj7uyX8xjPoe9g3qJZHyoqHKjod+zmjS9sb3fLlk8ts8/DI48/bltbm6miYnv7lp27+JBNzZ62g90je+mv/2975OKyXXj0nE3ML9vY6AnrjCA4vWMvv/TXtjB5VAAV1+zZr3/L5ubPWBdAhcERj4qKFqDCM/4E5rjjRro/ARVbO3u2tbPD7LCXfvADe/F/eNHe+uUbduHCBdvc2WKDa2TQP/HYJXvjjV/ad1/8bVKCMbOyUK8DgRLPvASocO3qdQIG2CcAqq9cucJrQnZMTIyxF8rS8gkCFZMTY7a0tGhzcwtqYj09J+fw8NCmZ2ecSqroUeHNtBHQ74AyyZPvUFFBfXgIkABZeCMGXmlUYRzsC4hGzyY4zOQgt1GbIAXQKBtz76IyAt0iHFyHHiiD4wisg/oJZfzxd+yMaIw9h2bgDlREzyHIkCagIsB7gQ+4D2QR+mksMKsS+wdAxdISelT0Kj0qAvwJ2RCZ+Ni7qaJieko9i9Cgk1RbaNItEAVjw3dCV+I6TGYoKhZCh+I9BNABVERVBuZQqkOBnRKowHVKoCLoJ/B82zsbXJMpzxoFSIHxTU6IWoXUhQgIOJ3RtFeHYoFRzRpzjvsBPImADBhNy+BdXc+XYy3/Hec7bIGymXbYWSEv6kBF2AYBVNTvEd9rAypoSyFQ44kVGEv0DSnnPu4Tc/yv/sc/vWegoi7z8u8N9EHpzZYAfB2cjMBO7e/t9zzmnSL5KSU1pbhL85j0uQFPoZKEdHfjqTVyrXypzWNrvnLQxcS7hE+Cb7/4Sng/QQtT1+MRwE5fGebyRUPVFqCirZl2qLegforfq3SHxa6pBfWoHRvWvxxqfT7yNiuBBPdPcT0PSKVzFSvsAUYFzis7uaVqSNSo8A9wzZKuCfZxPZivbZTXWoFC75OgB00Nt+OTqbJzYEAtRT00JcL6q+4fBTEjg1jvhWxr99nic/y0lo+6P0aov5UucM6Yhx/n1EgOlkQwl/SqHuRt2uXw9WJft52vJnsuza6vZfgh9Yh6UGGp9j4lZPNBqtSffncmFiobW8C/fMGgouKeYXIcdDz6CniSmAdLc28BUBT1aDsgoB7zgEB6te9DXnCGzgli4fpqcB3ngvRApE9SFb16C2TwhEAYA/1qvszG38xOD0ohzRjH4cl9oihWHKED/v6RUZsYkx6NKtAOg9EToiwMKmD4hsoqpG1GXROAnSdqQSdHtX7EGUJXpl4P7icFSIBxkNYZZw0VMkWPCthE6i/hTeIJ+nQ5Xh6FaFTtzb3TmS/i7QxoAwjx6iYCLBNuxzklcQBNBA+Z4heN0eVjc897JQKrJAo6x7gunhufiyD74dFh6o8R9g72DoAj9CidmpymncoKB9iRaDjtFE+x9/ET1yew4Qkgqibp09bW94OyMIPtoFBSBocAL7y45vCpnY5ce1iHI5+1LEeTRAiUyo9KVGfwfaffxvfJvOB7TcBI7nOLf6s/iGhnpasgG0V5RlpZB3ZLkE/XyRUalKeg6yrOicYpWY2/x/kNucL+k7D1A1R5AFS0idwHf/+qzkCqqEh6xdMLQmMO9KioWYMJYAjFf58zcRdG/ZcLVDSNM5fUJeslwJrG0uByLmpIe2HQVZyKIc5Gcw5XxQzJ1p2DIekpCkurzV4f5k40fScChWEIyCLIHJOqqIiAfFeNtA8PGLhNPSoqQMUe/37l6lVeqgx2hqJLDPHRBK5i5EtN5M9GdkA1wJiUoCkYocA0gIrpVCYKzu6gm0BFRSjJ4BVs2h3kDC2pY7xMMT6LcSGAoyanokxSVpGaeTJDHdkdoGNwgxlzBoc+MkxZ/dDrMHMSxgIyJ2FhQmEjw7TXH1WPis1NBshmQFsxO23LKys26jyZ0aMCWjr6PIjDs436ScY7jaViXeK8ofoDWavM4nUgJgcJxA+LOV8D9dONm6w+QOAGQEWifkLzLvxHY0qVJiVQEXNI484pSxjIQc8GNJ31RlKauGzU4RnRo4JABXpUXFy1s2fPpqz3BAzByUElC9cEwBUoNpThjMqCXme/ClT4/sO8v/nLXxoC1AhWnj53wXkiYTjAiEbwTyWfpeOhPapMWKACWP8PP/jQbt1cs29961sEU/poRF5wAgeIhtJWBhgdqMCeeP/d97iWX/va12x2ft5LqRVMSdlC9PFA+KKKip/99KcCKn7jN+hEkGPeqc3gSMngRDOyA/vk4w9tcWHKvv3tbzNrG2MIgC3Oqjhmw+jOvKBD6J0HjlEl2D0ksFB3VStziz3qvSPCiM0GvJfuFxUq5XsliEFx1hBYKEGWEkTBfsSZw56uvjDj4sjFf1UAlQXk6eP1fRKl2PGB8jnLbL4ywBjjru+3qMpSjx1dsZSV+R554iugSlTm+QebAizlOPP7kG3UFhXqJ7TBXl+7br3eASnqrt24bqsPP0zQ4eqVz+3U8rJtbKzZxUcetYmpk2a9cfub//h/2YVzC3bxiYs2Njlvk5MnCVSgCuOVH/4Xmxndtz/4w39O6qc7m9ftGVZUnLGjLjKgMvVTU+BJzwqHPPSG5gHNECnbrW/rtzfsCGeyc0SZ8vxzz9sbr73OSqYb6zdtbm6WOmVpccGuXv3CfvPbL9j8/ILt7u3QUSn3S7lH+u7UXL923dbXRfsEubm2tkbaJ6wdziiAClRUnDy5TOqnqUk0cZ9jRQX0BKiPkDEOWTw3P0fAcWtrmyA4ZG5J/XTUj0bGxu9BlgmYhPOuhtfQgwBNAKBAFlAG5ZVk4ADgxe7Bvh32pM/w/AByIjiBc8GKCmT8k1JPji72h+6J6ohcUcHsRM+yY3UAGiBDPh0esodDAjfYiweUBXBiJ2xudpHPvrEJ0PyQ1E8BVKSKClYP5uy1BFSMjrDvA/R82aMCv+M8RwA8mmnH7wQIDjtJ9+HvqU+DGQH89fX1BFSwR0Vx7vD50HOYD3wWP+OeIf93tu+ASZDXhr7f290l8EOKp3GvBkQvJO9FQlpI75Vz2FHlqPbPhDdXN2bNjrIHlF4BDLASw/VGk51TnvEAKkjr6RzbAVTEXi8DCfHs+AzmPhqYl6BCXD/kVehojCkqKsoeYLh+gEcxnjKZAu9jjr9coEJ2xr28Srq9ip77MoEKZt26bC+yuCtYxF0Nug1safvylw9UhBaKuSoD9uV7EUys2/3K4A1pVbhGRYPoeJqwUZK+Lx6TtgaoC4e8Bm2cdrAqB6ryBUPvx7Nmd7uahFEZQmQ2FxUSvA4+5NnXQY+a/p4PL/+Vt97geGPqoiE05AV0Q2RCN01HaROUlRLRDLj+nfIz4cmqGsVZAAa+IF3cfO+8RuE7Ej8gBXGV8qWYeaeOCSqi4J9vuodGWNpdEUhM+4iBX9nz7FXXIiOgj/GK9TnuSJa9K0qwgt8rAqmtQEax7gM+rH+JmeWge/IeXXjaoIINpR/JSJDNDExrgtOc4DakyiGQJUoq+AWRrNX0nLCAy3tin2GOoeOmp2dZ+SndpMbQCOaLTmiLOk0VFEeJTgo9J3jGmLImgEK6RH4d9jBsAIyLemQMAXIFwgnOIEFkT1RS0VuJ1YcEKtA/Sr4S1j58KzwXvgf9FLopbPes25TYhcQDxRxGCUJwH/h9ef49QQvPEXYSPkcwhgmMwVwguwo6FH53yMdI1pQIkCQJO159JgQ+ko4L9htAEgcBMLdZZoYUUnURA+8uO/GMeL5UTeLUl2kMHjPZO9izMfQ1c0FD6kqvHIZtSQDCm30ziO/0uBhzJPXhPtxv3quCz+NgWN0/if2l+VLjcDwFq7tIXZX7gXKeuPdaGq2HDCpAQeoCj2ewstj7dZU6KPZ92cdCzB2qMAk/XnYJ9puYHCImgGeNeFPqMeOVFxhsSe1U6vWwswL8kHx30K9QUA+aaR8nbR+8/5WbgWqPiiJylACIejQJyiH/7e7Ag/YQeSVQ5JYMzZjGIFZzZIt/HbjFkChYthKHrFf5far0Bl+gaMRaA3TScHwes0rIRiZtkHIEbc8cFmX9WsMMvi9rJ6Zyv3iijG6LB1VABQwB0gOwuTCon/ZsZ3dPTbR3d1hVET0rrl6/ngyPUPL3A1SE8R9Odyg+BbvlxCg7ExyFU5XgAII6oAkgwh+NJ70nRZtylBJrd2jCYYZxBc5y7BkpYQWTRQuBn5GxL8ccGZAwRkLxUNkiw6noUYHNh4DR2MSkbd6+w+A8gj+zrKhQM+2xcXEfEqjwhqg8Uqn5UzP1Uxg62dhRtYTOtpryIYAUxmtZURFctbBO0Ewb9E/LSwIqTp05Ld5sZKs6FQMMJ2TsS1krC0SZUjIKuKYjmC9xk+Jzh7sAE5RZgSAjTTHyp+vZQP301ltvEahAjwo0vS2pIzj34Gpn2aaACjZXw1g6Crx19ncTUCHfQHOF+/7y9ddt2YGKM+dXvYxWXK8lUKH1K4E0MpGSygP7BkDF+o2b9pu/+Zt26tSpClCB+4URTaDCcU/YHzDK3n8vAxXoUZEdNd0vgnPc+d6EmxUVC4v2zNNPc+/DWGJPFjoFogQDeIbnB1AxOzNmzz77rJ05c5ZZHQiAxSsFhgyNzWT8pmoY59FtdFKGVWvV2ghVgjvuRDU7PhmoiPdTAMD3UD1gHO9X10ffLt8rf6/fG3MQAdHqe8hGqvKWZmABD5mDhXWgopQ19fciiBmGbyVIUAPGsJbIOsZ/KHlGVn44VNWxijc4XsPAiNjPbaqkBCrw/LlHBQ4CMreO7Nb6Dese7dvU7DSBiocvXbLdnR374soVO7W0bJuba3bx0UvsUWG9Mfvx//Of7cTiqD302KqNzSza9NQpAhU7O9v2s5f+s02PFEDFxnV75uvfsnlQP/XgpKB8HtRPjmT5wPO8itZCoIqCOJFxhfMAEO/62rpNzczaxx9+yIANnGT0lYFs2dzasNHxUQbpNzduUyY8/dSTlBtrt9btxAlQVeWASGVu2WOgY9ev32Dza8gNUDmB8gkZ+fie+hygefaCnVwJoGKM4EgAFaiMQJ+AEqhAfwnoGOxNBPQBvoL6CX061N9ghNRPAVQo6wvBgHE25z50oIIyEc4fssBwzgGxOVCxd7hvHVA/HR3ReYbjHNRPGag4ZGA9suMwx9FMe35hnnR1eAV4gflFRiH0JfREABXIxkOlGkBB0TTA4QZQAeqnKa4D/gagYoD6yZ3e2LMl9RPGHcAE1iZ+x7OUFRWqLpF8wwtzXQfp+V7f7M7GHVKBYe6lczJYFToEf4+qAwAVeGGt41xDBgRQgYoKbEoCFXv75JYG5Rg0CQBx9B7CXGGeA1TCHGB80YMLz4xXHagIeRJAxd3Y7mGf1YGKMmg8KD+hb9HkfYtrWgcVYm0CqIi5xvhCz5dABT5/d0CFqJ9wPtT8FM20sSYK3pTPe/yztwfmm7872AS4Pi9tcrTp721yOQerSl+tyf/R39q9oC8TqLiXJ6tWGJRz2VRpgStHBnaTrq74j8Uw6vMXPmIbUNHWoyIuWQcq1Jdq8NW2bqVur+zDIXYOrxXKus44EAkWQe1UfjbpvXJ8zUCFbOlst+KekMvlnFeuUhgPVf3WaiXQnpcfosz3hIQX1QBcW9/GbUBFmXkcvkkEXWXLKvlNNp4AhQgmRqNg7ienxxoYsdO/8Jrk1XewwfsrpPPslEHBrT9wHVBPAsi4C6aC+C6Do2WEwZerQmMU61pPgqwEFyIom9c7hQ+cOku2aQZRqMe9NxLWnZnhrkcV4GfXQ694kK+G+YFfgvFxv3g/iTbfOcAE9XpQ/wJlgot3H6NVZYCS+qA/4Lfzs+4fqjrUqXyceofV6FHV71UuBBeQjMG9PWZHzGT3yg2vbp90EIaRHSau+TMgo90rQLiPwIDgyRuYEwIhTolWVveEThWI4zTHnsjJgLk3uBdFqNYmKhMiez4AQr0fCVd96nElhOam77EX2b/A+ysIWAC9shLKsG6qjNcGgZ1AOmjXh+ELiR0gkne0yTBOJpjMzjGeo7OnM4X5ZdzE+yOQrtLpjTF02DpIWA0Ag3SizrwxPq6qKAApYRPJXhynPYpkElVuIOEkN49OZyxAN1bgkBOT/igBGFIf52qcfF7L8GBVI0Z8pHL0fJ5LQIDngomWorVSNRVkjmIlZK1wurKgMwv5mAAP2IZMltQYywohVYOMMFZQgpb8oO+XAHcTQMeeMGZHqKYoY7IPKiralNGDv39VZ+Cv/vx3qpuc5zgOc5OZi4y7XwNQEdnpRBbbgI0hQMWg1VH8ZQho0bhwcmySNKGwUMleftXnqH6P3IYvvZPQdL90XMwDws17qJjrmtvROkstBtKwoFST8xW8l3z8JMmj2ZgcCARIILCrQMVBAVQIpMhAxa6t3brlvSM828BphDSGzCccges8L4QK1KfAS+ZCeZM2A1nyTu+D7zBzIlVU5B4V+C4C6VGq2ic3uIISkXXYdp7rwcLKjoh+FaNoiomMxxinPhVBDBqwHnCH0kMQgM2q2exYWb8MEHhGDqswlEZBoGJnc8u2NjdpRMwtzNvU7IwtLi/xPd7HnXJVVuiZEJiKwEkEH8qxRxBD46wBFd0Om8oGvUQZpK4DFTeu3yBNEisqzpw2UFQQqEDAABnHXlHBzK0y2F3wWNKxATWUl4R29g/Yo0LBkVymHdRQbUBFGJkwkkX91KsAFbBsEDAkXcjBHo2IMuANgwPBoddefTX1qDh7IYAKGIQy5gYqKjyTQ6dGQAWMjQ8uf2A3r16z3/rOd2xlZUVMNV7GjJUiUNFX34wAKmjEdnv2q3ff5dhQUTHjQTGeSzdiYJDqdOQeFS//FNRPi/bcM88koIINvbzBu5yKUQbsPvn4A5uZGbfHLl2yc+fOK4B5KDoyOW7iv017CJnCbpD3jwEqStlSkUE1oCLAF55D50rOIrKQr8gGduEX4ynnogyilfcL5zaCVtW1zpUYbePFtbCvEUCtvtRMmwmuFbkkD0yZ/nqVAYtyzPHv0tErM/tKJz3kVOHx87pYR2R44+/IyBcFXYNeas8bGKCpGKYzSrnMwA2vK+qnBFTcumGdwz32U7i+doNABajaPr/yma0sLdnW1ro9fOlxm5g+adYdt1/85Ic2Ztt28fELNjW3bNNTp+1obMZ2trfspwAqbC9XVGzcsGe/8S1bWDwnoIKAkHpUlBmyMef8yTOeM3EVDFIwHwHytdt3bG5+wV55+Wf29DPPsJLp1PJJOmZwJHDWUTH2+Wef2tNP/4adO3Pabty8Tjlw9tx5yahoBl9FhGxza8tu3rhpB/uHBC0AMHz22WcMwmKtAqhYWjphyyeXEvXT3NyMzc7O83NB/ZSAij6oANE/qEswQzLrUICD60oMY2JcQACOPIEKk3M+NTXNigo0faxSP43YGCgL4ajDgewc2hFl04EqKtg7QplhcCzxN8joJqACn0P1B4AKzDfGUX6XQIVXfAEQxz7G86EfjHphINgNWsV5m5qYsq3tTev28P4c57HSo8IDLOGEl0AF+mThmTH2OC8YfwlU4PniO3F+AmwpaQ8DVMZnAVTkhtx3B1TguRIA2euxjwvorzEXaEYPoAJOOysqvaKC1E+jquhAoEXBETSXRAanKBeikgHCCIDlSK2igoHIMruzxdAJuTEMqMBXQ9aWciK+A8AHax2AdimXQ4bFeGJMUVGBZwx9gO+VFF5ldUbI/1xRAbBvEKgos09j3C2PHpJ6+Nv1d2GzlOe9eP/uZGj1gm3fqeRDlXK8xcU5plCg4RmHARhDFEfTlVrmo21iK7Z1bf7qauye5zQCvzVaJOpd3uveKiraqJ9Cj9d9l3sebz2gXgAVecy1JIu2/Vd+oZhXgRQ5w1tfj2BolSGg1PXx76ot19RhsQBayp6NisPyFUHq8t8tBRU+tsgiztF5yI4APWPeoQejOqJ+3oclm0WSGxtNI0ufmePjiSu/XF/x+zf3eOiDc+8eXrJDSj/bbUdfj/JSddq3egalbMgaUIELpEpSXY32PALSHafdQeLVoaquoTsY8Edw23WI6HZGUi8SzDXsDgavGcSOmOrgvWOvBLe/ekmJ0in8i6gOVwKkqgrYH8opc2i/OYCEcSOJJD6rBBT5SvgH9DwAD1A/TUxMJYpd6AmMGUmABGHcXo9kOQbhPeCvbHf1XcGewe8zSPhCIhn9NTjxI6wkhY+bKj9I36MqAekn0T5pw6s5ctDZhY5TT0Cn5jpSggn7EyQ66LBZc8Y93otxl/sj1p/0XJhjp6Ji4J/XFE1rAHEM+HvjczwTbKoIvotCOfS8wJWgOEIfuKgYYKIEK33VtwxjC5quOH+sROJA9f9xRhl78H4TAJii14lAqNo5KuQ4xoVn5T7AWrkHnL/iiY+sJFI8pQm6575yoSN56B9z4YT3A/hiJREABQdbGJNh31GvSPGnC7kW+x7XxdxAKrGxuVM+q6cQKm4kb3voD+nAm0vjtLTsNVJU0GhdIfuOmGwbrwcVFfcgeB989KsxA3/159/LGzxH1IvB1xXuEKCiVTe3G7iixCmij9W8gruaxGYBdG+GQvVGTUCFeMjz63igonLNmqE5OOnDwZmKGRhVDjXDdDAoVX2qYcZy03fLEd0NUAGDB07zPgLve7mCYntnu1JRcXsLgRWVRyYDMwXII7zeVBpclL0X5d3h7OZSQjXfDKBCFRUCKgLkmJsVLzUUEJ4zMvAVxM0KoTaDboyFa5MzHPAXAgpukCDoHVUBbCbN51NpqIwXXRkBLvJ+Oyc1KaDGFBSmEePWH5W6GzI72zu2t7tn86yomGfPgsXlZRtFYMLHQU7DcASYhSIjk+BA3DwF1CNTxbkeHbTRuVTjbwAV3UPQS0yovBEGJp9BhmuqqABQcfIkA5MrZ86qwTj5pr38FIqVylilmhEMKuccQTTxlaoPCZq0dlIz7Ww0MbMA2ahbRUXF6qqdPXeu0kh0bETBo05Pja+1X8ZZybK/f8h5mp6apNGqpmNhbchw/8WrP7eVk8ukfjp34aKyYzzDKICm+tmiw8QyVPSoEEcrKiquX71q3/mt79jKqRWzcWV/RYZXZNTQEI7MMAIVXXvv3XdF/fTkkwz6RSkvy7ILyowwBfHZn/4E1E8AKp5lOTMM8AAqsK1ULj9GkOyzTz8mUPHQxYs2NzdP+iyWrJKGSh3eKXZ8/7IyaGxUGdcFaNA0D9wlhcyqAAGlRC2o1CK4rE2vEt78EuFuPkvZqY7sQIERNalOG9SNZEeCygBWCZSU4+V2YPC9z8yzhcV5ZddQBmVHf2Q0B8HFV5ubAMa85OfybVbLUKx/LhyV+rxiX+lvWQ/hrGAtwVc6PzfrAcmQ4uVktOvGtoy44YoYcjD4WgFUiEca1E9r69etc7hj8/NzdmPthj30yKOkKrryqQMVO7ft0cceI/VTvztu773xmt25/Zk99tSqzS8u2+TUaeuMztrezo799KW/tsnujv3Rv/gD+8Ubv7StrVv2zPMv2PziWev2wenrFRWqZWsEXZhl6Q5NVHfB+8V6QR5sM2A/br949Rf2W9/5LfvhSz+05599joDC8spJ297ZssWFObtz65Y998xztrSwaD95+SU7d/aUPfzoE9bjflCSAtfa9xsc85tra7Zx+44ddQCgH9jazTX27YBMghyMSjyATAAqcGYnxscoS+fnFljVBsACgAKC1uj7gHFvbIA6sEcKKpwTVE6RaoBAhfbgxPgkHWpUs+EPlK9+Tz7a3uMAACAASURBVAAnCuIDXFdDTOoROOMOVKDKC39HphwC99FMmwkCBVAB/QB9y8y+vtEWwL7E+sOZx5wE9VNUGkS/qKiowB7Gv0+cOJGy6yBvZmbmyHuMoDUy53BNzMPt23cIFLCZdlFRgfNfBrjZZNwBIcxb/A6qxtDRAKIEHKGiQsEaVtx1Oqk/E95TduEIe05sbNwh3SPmYWx0IgGWZRA9Eg/W1te4RpAjkXHLigoCFWimjaaUxqojzDPoKVhRASpJNNl06ipWgHiQB4AydAR6WOE+aowOTmgkB3gvKQecQ57Uz3MdRAi5EuA01hG83gCbgrqS33EO53C8CWizYnSE+5XZktAdnlxSCuUAYgcqKjg/k0nGYqzoSxI9K0JOB2ARdsT/9Hv/B/fHlwNUhBFwVy4I7SS5B1U7/n4C1NI3Lf6A9wVLo2oS76VOvTf2qpbSjMEA5KC/NDhPbbQ49SB+0wyXz591djbN7nleY558XmvWhCg6h7wGNeYwKqzCUikqH5PdU2TIyoJufpVnip+JatFYpYISaiAL142fBAS07afUAFe9DeDDwCci33/jqwxC5383+57eGKFoXN2SQ1fZzm1ARdhOorYMX0v2IYK/8Yqgb1mJWrHnWuZCmeb5CDD46feKNSorTVLsomGeovC+vG+b7E3nPYKwFZDBfcxyl9Q2bz4feqMNqCAlbLAHOIUTPstqa6/ojyz3qJiALcHqNgclWKEZPQEQ9GdynTeoJmhRyq7csBx6izYE+2OMUg/jPySARGUBg8kOhOAn9B+mhP4j1tjpfdRn0KlW3T/AWoQegY0iX3zUDtH7EVRI7IuoPpJBVUz9TFAh0zRBt8FPUrBd8YkAZwDgRPUA5pmNy7s92mlILmMvLVR/+OdEm4R+YLnhO+ZHPTfKZMBw81U1ActLTAMCgvD5sJ2YqOmZ9BgDPgc7BuuYExCM9gXsFAFJ8jEx1gBNIj4SPoR8fSRYTtLewdgjNsNnZVDcg+3+b9rY3nuE6+ERh7CVRLEMYCgS3np25MAeAv50J2EXYJ2w/zzJB/cKQGSg2bufEX1G6yPASvJbFcThkGpeo5m2jmmDJHeqp/h+yIDwhTA3YavI5snVmbw+K7fEmgDbA2vEytBRVb92SQ+tylKAfoiTRfVFXXSwwsh97XiM8nxjDeS7Z3pT+hplldWDioqhuvzBm1/BGQBQUTUe6gf5vyNQQauqUgB5VzP6pQIV5E2J2xb8K/W0BRd62RAZAowMpgPl56q8V3dOyifz6xefL43140CKZAw1zGjbdweBCo2B96WAFmoeZXpAjGGMJKCCdE97tr1bAyp2thIXcWQeCFnu2/joeOJIHXCeBwKP1T9E5l5pEDLo0emw2gDNtONZg6ohlFHJO5mMoDTXngfgRpgCUCIDQ5Y+DWKWq7rxQSsPmfTZOApnOgwQIuiYP/QNAFiBuUNWaqqqaO7hgfEjkIJA1/zsvM3OzbMh6tLySbNJZPlXKyp4nrzhFL6r+2cjKe1f0gENAhXITD7qdmzrzh3rHnRoNDLbBuWcHvhlNoJTP6GiYiWAirPnmLHLoAoqKmg8Aqg4st4IDEsZrJEVEg5sABUwBDF2gDgJqECVilNnUVwgwLi1ZW+++aadAfXT6kU7t3rexienOD6ULCNQgv91DTRb28lgRSCFFFsIinBuULmiLFUZeGq+9vqrr9ipUyft/Pnzdn71IS/pUKlmABUBtFSD8J5tRN7bvn3wq8sCKlBRcfqU9bxhHTNHwM/qzeBg1PRhrHhwHO+9+847NIyffPJJm12YTUBFyABWVMAg9f4UMJJe/ru/Y1aygIopGolsKO4VFTonMnQ/+/QTm54as4ceusj1OH36tC0uLhpAMWZrOHhFY86BZRqvMP4Z0qxl99XkTP0sHyev4rnS50o56Xu63McxLhmV2Wmt3lf1JhJiHHHxX3Nj7ngMZMgpUGa2sDgjsG4E3KzI3MJl4DwjAKxsNgSj0QBYvfly2fYg4KDzWT5vdsjbgl54jqJZdF/l1HgeAcAdm5j0fgO9MNzbMiSrC1UJEN11RizG0y2on0SDMmJdW1u/Zp3DbZtfmLO1tRt28aFHbWd72z75+FNWfWzvbtilS4/Z5NSSdXsT9tnHH9uvfvULe/bZh9hEemL6rB3YjB3sHtjLP/xvNtbZtD/+l39oP3/9F2zS/RvPftPmFk5Ztw8HAYCwZyZhPEU2YjnHylkSZYEC93Bke6TxwdkAZc3Vq1ft0qVL9tprr9nzzz9vly9fJni3f7Bn1j+02clpe/zRr9nM1JS99NJ/ssceX7WHH/2adbuj1u0hiK1eD9ASuNte54ANxEHL1DsCP/O+ffH5F96zQFzAbJ49NWHLy0v8T6CwKi1QLYFqmblZ9KdRphzmVEDFjh0difpJjvChN1PsM1iNZw8HVBRx2MsKFMCxgmPK/g3gm/Zy+tgVpOdDKf/BAfVDUADRAXMOY1wbepaBdad+IgBtqFLZc6BCVGS4RjSnjmAFAIboUYHqiOBlFlCB8StxACANmoSjEgXBBQAV6PGEeQFQgXkqKyLxKAFUYA5w3eiJgXOZgQqcZ3FuQ/aCGxtOfmQi4nMYsyovojcE9Peo3bm9YZvbAJBAOYTvTKaqs5BJoeMA4K2t3awA9Nwhva7tbm84UCEaBYBmGIt0p0Di7qGyDaGvxqcmKJNJo+BVgVgTzBP0mkAnJAe0UJG5HRfykUGbAOnDoS/6AEWVC+/h14zvREBQQR0PPvRHuC6w70AhRlnt9AaxtyIpJGi3cD3YNfgsgDX1fME56tvWFnp4VLNTY334+YkJ+5f/9H9vBSqiii7ufZz+KWXHXTkhKfczbMUWoOHuLtYMVChaLfUV/siXDlS0DTAHHeufaAs+Hwcm1N+vBJOLm+hzRYB8CJAzYDf4dcJTSJmz5fWVez90Zf6+QAVNprR2fqtj9CufOke8UxDXuZp0kUgAYfZxfgWwoc3SDqoggzfOJvn32URXQeDjXsetr9Sf/Lry3LWts/Z1e21L4mN3aiclpWgKwmdj4pT3MGgCKmQnNZ/NAGVpRzuNC30nrxwM3aLsZ1QiKODc9KpXVIT90TqvAV7VwYoy8B8hgEIGhC8eIptzWHvGFLd1n5Ny3nspYCowJgSEcS0AClFlwQpIJC3QvwV1pYKvtLFJXwOKKwEPDNZDdsN/Sts77zvYJKBtVPBegAX7IHgz63KtYk+z7xKTCTMFFD8fVE/u12LMtEAZiJe9y7NGKiDJzPAVCJyTyiuyj3TGSDPsCYrwk2LOSHvlz4/n5j28wkLbG3vFkz+8VxLGr/mJI5r70DA55siBBwJhMdZoat1Nc4j9hnEL0EGw34PxBVARQXT6nxH49z55WBvZNdo4qjzKLBYBXuA9+OYAKvBsrFLAPQ+1v+UPq3pCdFxKEuv1sfaipBY4KNAHsQzEWtC3ZHoSvcwcLGGsJGJI2nc6F/KPxCggMC2ang+AlmlzSfYlgIaVNM4o4IsXFUO071kdpb1QviKGEFUmCax0ai5cHzIxEhgxTqxF9BplDMf3cJpHZ0nQPmR5Ne9NewwVOJ70w3hMgHPFXlF8KcecJBdj9E7rzcbsSrLlviwqux5UVBynuR68/5WbgdRMu3Xk1YONTOLysN+FPaOYUE1EJFPBLY1kWCV6hjZDqeXvlDhx2iMQFRqzAB8Uz2l/1a/BB4Q2rxs3fpFKLXZ54RA2nok8IB6TGkvDaYNoxMZfPFs8lqSUP3hxbw7VLbjKfduMtPqE5N9lwJfvO8e5I8nRDAiKLHpU7B8cpoqKHfSqqFdU7GyplK6Ya2TZk17jSOWMEVCvL1SboaegazZIwulmk08YWOMTCajA5xDUgQIKvsi4X1lRUb9XUiBuPAZQEdkJMHaUcY7tovLVyPTB9YOLe5wBDZUY9ryiAvRAuDdBi1439awIAyst/8gIgxgIeCFohSxagAHLJ1cqQAUUaVAjKTNI81MHKuJcRsYAla0HLGhIjKLssWNbt29bdx/lnZPkkkSTTjSd5dZwow89KtAsNoCKU6QQUrYqgrZ6Fi9VRKBwvBmoQGgPc6igWQ2oYL/cER5H7sq+sbH4m2+8YafPnLGHLj5kZy+ctzGUVzKrftTG0cQcDsxoN9E04doIruHFQEkq/ZR8A5+nKgo69otXXrYzZ1bs/IULdoFABW4b1E8dBvpi/+U942cNAWzGbXv2/vvv27XPv7Df/u3ftpOnTplNeEUFjCwAFU7lgeySACrC0Hnn7be5fk899ZTNzM94Q+98OgKooKHlzsdPfvxjAhVff+55ARXeMJ1nllUeOGvjHP+HH1y2melxu3TpUd4Hhuq5c+d4A4KII8qQ5n7xjJJwvtUCrqkCqhBbBXd/2xku/14GHI5zmuP97ABXy/Era5K6anKne3bS8U45ex8wCNe3+QVx2o+OTLBRNgAtgmvg2RgRVzKACgTOZQBrL5TB8piZYaBEO2iABS6esa/sogjG9foArQJAvXugoglEGaIpi7eqQIW8wC6hQVRUHHV2bG5+xm7fvmUXLz7MioqPP/qEFErbu3fs0mOP2dTUMoEKyJCfv/L/2vPPP2wnl5dsYuaMHdqc7e8d2s9++F9t7HDT/sUf/4H9/PVX7WB/137jmW/a3OIpO+oBpMhABaiBmN1WALDJMcKZ9Mwk7AGchc5Bx9Zv3aJ8/OSTT0jvhcx0zAn+jeAvdAb8uZ3tW3bx3KpdPPcwNfNLL/1He+KpR+zhh5+wXg9OMBwu9fLCvoDsvb15265dQ3VJx/rdvu1so4rpM9IGgbcXumF6ZpqUgSsrJxNQATmFADmqCTQGVE2IJxd9H+Ak37mzw4bgqITCi0AFAk7O34s5CKBCAR2MepzABM550DlF4Lc8b+EoQ0bgOtCl+E9NrpFBBuAafTH2KEdKoAJjEfUiqh+GAxWQT/hsCVQsLS15ZqPGjOdjM+2NACrm7eBwXwDO3NxQoAJjgbwP4AeqK6pIRLmlqkfMRR2oUJ8rARUCADB/0E1jHC+y/Wfn0BAcgXXouhz0D1lKXdbrsnl60GWFnkXQpg5UJOBnAs20VWWKBu+wWUgzgcoL8GqDzpAVFcjszEBFZJci0BCAv7Kui2NLikXJvkE7Q/zP8X5UlfAe0DHQz7y2MlcjoEeTNCoqakCFlHqWtZGxWQUq9pnMAKBCFajI7O7bFpuN5x5b5ZgjCeSPW4AKVKrI7M+OSLnH26T/XQViKwLynssXPOimZSldjDY3Re5GbR1bhLSCMEPebHhLMZ7mQG6Ye3enE9qvw3cagvRN9rbuVQVJPIRTGWYecfPY05hbwIGgBKw8W3Ep2nA1jdc6D7WKiRT1dDe0PoQU0IoLBvhQJO0xCMngoPPr1PoTKmDd1JREBnqlYrlszu1c7/hU6hGQBlg8cdh+BA498/uYqdbSOd0ifykzkT3w5v5r3g/eeLk2ufmMlr5prmivr5vWU9n/4ftITikpaNj+U/BY8g2fJSe9yzhcl3LJg5FteyCdu+Qf+f4pGveW3033dN+LoG+x5k0ySv5oBrMiyBpgXOmTEHxyf4or4msXDZ+jjw/fYBA0ssTznopmz9GbIsAAzbPTLHmT7VSVExXjepiisjpcR9+b6N2AILgnP8WcY96he1i9PTZOKifMFfQgng9BcFY4EjSRz6aKRwXN8ZjKo1MAPPWHYC8JNAv35DyCF76fnE6Hetx7ZsT54nWQze+Z7wFaRDUDg/yoxkACAZJCvEqA33caKDTtjrMc+zB6gwD8iuecwFy6LMD9ggoKiQ2kJmMfBwE+eLHywule6Xcwlw5jjWfMvUSCAioqIVBFgs9yLVGbHI2qoa97xnkXE4PHN9hrQ8AD1gC0n+iZiTEhEQd0obCl8Ay4P8eLhJMAfTzpIJg1ZGcCCFECVq6KUrUzgB+uBXuW6HOhz+Oa+B77kTi4EpVX1CsEGJQQRN8X8iEp2SwfubZehQL7mPRg3pAcIA3PPYGppJlSYm2cWdpGxTkmCISxdZS4ir0imaxkzagMwWci2TZVc7jcEXOCziRsYbJNOMVb7CWMjXP8oKLi7k2UB5/8aszA9//yHzcPNFIVkvHk/yDfS4ParPMrlldNcfbcoLc0TGr2WQ1x8HcrGbW1+zdq8bAQZCBVwZX2wFSrcxKk6DS+CuCgYqxVjSjxluveTdRN9b+3Jdi0BeqggJveK59B06a5iDoAzWh1DipgSHLolIFMih0+p9ZeCU4SnGga1uuKvqhzdGj7bKYt6ic100ZTba+o8AqL27ugqpDQ5lWdQxGC/mBHNAukUUB2R7Hu+HdTMDP2TxhmpcAndzYaSo2NJ6AC9ysrKkJ54GeiogqKm2KeZOD5fz6jYQREFkIYl7COoFzxnAIBVJpJsGIazUMnZTg5wENHyK8NoCIaeEbQI97DtRAUAlAxOzNnCwuLzUAFFD/pKZQRRJ1cAypirFRwRUCvDlQgQ3vz1m072j8kRyeACtBOIPCtUmAZ9mikXQUqLjBLmNnnbGqpwAONkZFeCpRR0ZbNtAvqJ4y/rKjgFkTyRwFUoKLijV/+kkDFIw8/bGfOn7dRNPjiGo4aYApUVQCokGEkbvVYaxqfqfEZvoP3lKGDoNyrL//UTp9ZsdXVVbtw8WHZKJ6BgnXa399rBiq81wapcHo9e/edd+3a55/bi9/9ri2jRwWBCnc0vKICYxHdkhrY0U486trbACrMCFTMLSJgWqX0CG7vCBLhOiVQgWBcAiqY4SJjEDQyOCPvv/+eLcxN2uOPP54kN7KUESxkafSIMo55XiPgVAAXad+3qL3YUyGbMqiQHdamQEWc+TYZWJV1MqLbeIOZCUQ5Hs0xgppJcqjtHhT5Ks8hGDE3P61muCMCKwhUsIcRDHJl9gioGE/VFmU2YDlFSZ4Uwj+eqXy2ql4arKjQ1z1zi8Tknn1l8Yy5/LxliQb+HMby8Z+vUj/JM4TjUwUqQJGzuvoQM+IBVGBv7extOFCxZEfdCdva3LCXfvAf7IVvXrJTp1ZsDM20bc4O9jv28kv/1UYJVPwze+W1X9jR4Z499ewLNr+wYkd9rIMDFX2znb0d6qdyLuWTogquw/M4wz5F6lcACrjNjQ06Q2+8+SZ7wbzyyiv2zRdesE8+/pigCvQaQOaD/U178tITdnLptB0dduwHP/gP9vQzj9tDDz8mkIKNvUWRiUoTnLMr17+gbISshCMHKr3PPr3iwfMxm52dUY+KyTE+N/pUoKICe1L9D6ZYHYDKCjQpxHmfnZuhs7JxBxUVRlASzwI9TIeMlRMqo4e+QbY615Q6VcBxZDgyGOAyRY6UWwmuM6KiogmoQNYj9HwbUEFQxYEKBhccnA/aKAAAJVAR1E/YHwJEREUSQAWqGDCnuCYqXAJEir4ZsW/hKwYNEp6mrKjAWYEOxTMHUIG5hsONHhisrnO7JMAWfU7zFkAFgCYAFZAJU6hyQI+WFqCid9RhBQ2eG8+FedZ8dAaAiqgqwecQvKGOBvVTqqhA7wpvTAkqAQcq8JxlM/BY0yY5E4mZTTIWmbHlHiBQcdghvZToGop+RQUgyAAAxztiGwVQwXvA6S7MzkiOiIoT3A/7DI499ntUVOiZbomuzCtCQw+xD5X3Sfmjf/wnPM/NzbQ9c9Vze7Ksb/cFykzw42VgDWmoCvnGrx8X5x1s1UfDu9n9ojOQz2zcsBWoaHkgNiSNs19/htD39e+2Pkgb4NH897vR8XXd2fQYck/uBTSKB6t9pwQqohAzMl1bst3oYzU+Xssz/3/svfeTJNeRJuhZKStLtqyq1gIt0ECjARAAyRnOzcxyZjgz5Owsd21P/L77t8z9MXdndmtnayNIaEWCIMGWUN1otO6qLi2yUp99n7tHvIiMKIEBzQizTkOjKisjI9578eI9d//8+9xsb3XTzA6xTmk/woC+ywkaAGDFfundRVm4GdcxqRDKOdE+Ul8EL2r6+/0Ov5oGKwJbL0xqYmAzz3H1fhgwEtp8advG/RPK6TiLZEcPnY5FQhbC/Ciurx7It+xlJqLlzA0GtpHZbTUZQmmnvDblzbO86ZdZHyNgKFAy0WSZsIY6Q2DgkbNEQR3/OEmFPrAlSAwAYgUE6xWscfYBAXBj49C7t3iF+o06T3Ae95mUvWLZ67BlLOtffTiVli1BPgkBdAaFNYDuwXROI4sVaaIUAt0adKYf5lr9VnxZiz+jKDSy2AtSqgCsUBYQGoYgOcfA+2DPkM5RZ39rpCX23+PRxNCRSQqpaID+CCYXYberb6vxDm0n7CfW5fNEPmcHBGymMM7jfdWlIlWQz5BPlypC/2Cj0dcqFVUqyNrEvY6BfmMmdG2cTMLYfT+0EZJPOAeSVYaQ4GAgkoaAdH0hqwQgiD8nvB5knbWGGMcO95Y3yovC257v9RnsGeVYwN8h40LlorxeiCY6IKkGdkvZ0rX0WE9O0FiARcIIJKn8nAbfNekL7SGAA0au9V3tGc/H1X7RpzX2rd4znTsAHjCP0UfYb1QBsX5RimxIwQ9fGzWRR2NmzhRBeyDvpQmUarfh8ojxuNxXZPdZPMPuesS1RF9Rx4M1JQBk9VDcXM/ljF76GMbu9WfLsizYx5A5kUw60TEkgPYUqNjpzvH0uO/KCHxrQEWe4cun1S2g3QIV/qiHP9O/OxaQcjgShZ2+LaBC9afjV97vtoLyQPceUu228yQD79mDmGfA7wyoCNvIpTUFUuT1Iel4eSAMDjqNzDSjotumQbJpGtbbARVO1aVhaHrKDJa3u6SQ+oaJvruRExnUKcAiPWpuPHvwHUg4sktr9eEoGIPgj8tXhNfw77jzrhugzl93+t1Qx8/QgA0DPBgfbJAxUKEbJ/8VRWrDFRaaprEFIMWMQbY9cDgptQGjw6IKXngbuuJgUwCogGM+Nj4h5XpNiuUiz0UNfbvTbKdtqC4J4X1wgw/987+F4w12Q6fbkpXFRek0WmwzjKECKKKul6weFYGK2UePKRuEglEHZg5Tu5tgQRHAEyiUKv2ExoFREQZS+IRYbQd+btkEjbV1GpA0aCyb0/uGzXllaUkuX75MaZZjR4/JgZkpKcLoQtYGYYpCBFTQmLbsDJyfxdqQvWQOG5810JeNsY5g1m9+9b5MTR3g+Y8cO5EAKmCEhYyKMHNN5YCUXYP2fvbpZ3L/7l350Y9+JPsPHpReSc1aZkABNDBgSSnWymAgKNDry/Vr1zgHAVTUR+scf5+baLNncyggpqDCu2+/zQArNPYRlGXGEEKnVkRbHdYy65189tkNGR2pytmzZ8ww10wmFP1Gdk2JMkbqyLlMmj8jSpVOAg7p96GTGj5bfs+9Dz4f0g7wboIYAA3iYGWcVc+sOFGquq5hKkU2ANpm0QQp5YNnGFJhQwySloqQaYHBzzBiBFQwQE7JJb2HmoGoAYG0U+/rXN5nvrZ5oFHfZwEVGH8tIBnVRmHPrFhhVJMjmU2YHteswEjYhnCtjb+bD1TMzj006ac6M9UBVCAj/vZXtwlUbBCoOK3ST92SrK6syBuv/w958cWTcuDAfilWD0ivNCaN9aZ89M4vpddYkJ//53+Q93/9ofQ6Lbnw3MtSH9sr7Z4CFbi3AAE+ufwJZQgxVxEIx3xYW1uj7BTkubBWv/baa7J37346I3jOtb5HT258+ikl1n7961+T/fTRRx/x/cLCotRquE5Lzp0+I2PDE9JuNuX1N/4/eeHSOTl0+IR0uqR8SY/zBfYOQJBN+eLrW5RXQvY7Ar4b6w15+OAhg+y1WoXBcsoXDZdZ42diYlzrPIgQxKhWMX5rUqvVA0bFCLPEVlc2pN1W6Seu430tgMl6GTaXse6jHT7PUM8DzwPGB+sNPnO5ppD+jnvs38UYkjWJTDnINpj0E/ZRSDyhf+6s4m84HufGHuiJAQ5U+HddigkBeZwXgX/cB3wH80OdNs0iw35HRsXSKs+NZ3Cjsc4xxO9poAJbJuaTBxa8jyoRpcAF5oEDFZ69CeBBa1To+OM4HwcEEzSBAnvEkMzOzkqjsUFGBYAKMCrCNc3BIPwEUDE3NxexUPz5QQ2ojbUV1iMhMCFC1qTXAgF4xgBAu0MpDBxTqlakz4KhyqhQMCrJqFBpLZWSCvd3X0MwNxV8jRNA/HdPXPE2Uv4K10f/kbEaMCOiAIXJcjBzVFT6iRrWLiEVSD/5eh/uJ2iXA2bVCmw1jL+uaRFQYUElHOt7hds0P/3L/5XzYyugwpf2UOc7XNMSv28TgB343iCyYEOdE7DPvbB+sGuggl+KT6pBqm0ukvqYQIWWJoteEQkxoxC1Lii7vEZOo3azx291RQ9IZh2THVTfOVCh3SUclz9t8gYkNZ/8DBpctlfK9sjbjz1Q5nVu9H3+zYYv4uAi9fxt7QiBinD6ODkjOV46Tm6LqK1sgeddgBVZ9yC0D/MSJPKmWSSJY6MY3X/YzxZU1vFB8pjKCIbrlw+9JlwVKG2ngUQ9FgHgsDBweON3DVTkjZMFVhnPDvRuknZfcsqpjRzblAy0d9pMXEMwFGAzkwltn2bg1zLameXOTHNfonQO+n3QrHMPACv7mr56VFhbGbvqqxToFyJZAaeEX6VMB03UQfAUAX7U0dL6RiqZyzW8qDJJyhAwFrCNBfYC7LXY11qtJv0Xyk0bK0ZlERWkcGkeJv+lZNCcARI9YrrpWWBXr0l/nbKUbdazJKAUsCEwLpFvF9XpM7/LmALJ5dfGbmB9NDBSt7VoHjqYQ2YKal0EezKuC7lHSEOrL23+i0k2oSYHaz7Y330JCX0ObbsBAMZw8OcQ46iKGFpLAjaG241IloFt7IF/2jGwA8kysoLf9IuUGeBM7pAtCYAAyY0EfQCUkJ3hBagdDPMEUJVkxfVUVswAA9a7UKlWB1p9G0n4lvasYt5TsqmgIBcBNkuo9HmA63TpKypbAw8Ta7KUVHKVc9vmCueqAWYEHQ/SQgAAIABJREFUOZDkQ+lNXSPof3uh+YBh6jXiFChp0RdBMowDlpqI41JjMdPJn3sf93DdVYgk3nf9vYKQ/adAxe7MkadHfxdG4I8RqIiNs3hrSQaTkkaiJgH8oYEKXxiSgX3bdlK3WiUfEk5DFDZWQ9ej0aFx/m0xKnxRGzT8dw5U+AbhxqEzKpxdQaOPgfquQLYIm6syKrTY5lZAxfLmeqQpyoXVsjZ53zuG6FtmORZ3p/bTEPCsoxywwjf4cKGH0dTu9qNikzgGgRMvCIr3HiAIGRV+PZ+P7hh7UNhBDe+DG8W6iejm5XrcvtFpBgIMNtGggxUqg/kW0R5tI2Jg1cbBAQ8YNFoEuskCqwjeIDA9uWePSKXEQIKagkp3RHABRqtvrmp4x9mizEY0BN+vnwAqCjB0nVHRlFoVjIoyszUAVDhlGdeaffw4E6jQAl7KkGGNCmT0F5SiG4I/0b2zZ8edsM31DW7uvPcpRsUAUEFGxbQUYQAwYFKMalRIUY0Szw5Sw0NrhACoUMcLT7RlVPQ16/ajD9+TAwf2UQoJjAoaJBhfGOSoLdJUWZQoyGPGFQ1Fk35yoOLB3bvyv/z5n7NGRb9kDCUYxQANLIs1ZlRosTcAFdeuXuW0Onf+PLXpHajA3zxQhN+VQqxU6LfffFMmJybkhYsvsJA8l6BI1quoWTeFEvsIoGKkXpFzZ8/yOnAAPGi0f/9+GeqrU4IXskLc4UCfvUBa6ICGhrY/R6Gxn/UcJ8cvGdRPO7fZAQd3uhSoYCaOZfpgrjFLyfTV9RnNln4K15BoYQ+AilIZWe4o7DtM+RcwKqL6FKxHEQAVUXZnvK6Fm4X3Az/TDnrYx6TDSrgpsFTdcfGaSlobheOOoLkBU1n2SNa4ptdQ/1762Hh/sfYQsEExbTQN2VBdmZ19IK3mqoxPQEppmUDF6sqafAWgYg+AihU5gRoVlQlKP62trsjrv/h/5dKlEwQHy8NT0itNyOZGU3711r9Jd2Ne/tPPfybv/+pD6bY35cIL35PR8QOsUeFAxfVr1+XqteuyaJJA6D+C3wBKkBU1OVmXM2eeIWCI4sdYB9bXGwQ25uafyNLyMuuz3Lt3j8yKK1euyDPPPEOZH4CroyNlOXXspNQro9LcbMibb/5PefHlCzI1dUQ6XQWouj1kN6lk5Mrqitx7dF/aBlJAZqrb7sr8/IIFrot0YAie10oEF8fHx6L1UWsjVAlUDNfqXJ9U+ikGKlqtngEVynRkMW3MS9NsxpqO55nPILPRdO11gAB7dpit7vfcA+3OKsB1w1oUOG9YoyIEKjBfXDaJwB4zLJM1KrAH4/s4D86LMcb+hutgHBjs4FxSoAJBmKXFWJILQAUC4ji/F9OO12LU71iO9pjBYtoaCHFJpzRQ4ZltmDsYN7wHUKEMAPSlQJbM5uaGDNdjoCJc+3z8KOfQ2oyACrc3MM7o6+bGCjNRMR4YN5d+0poQRQZzHKjQGhXGqIAmdAZQoSCFAhXcFwxkTjzDDqSnWKsauDEtZMuY9jodaI9navocSQMVZFT0JQIquBv53orghv2OfqM9DnzjfLrnFFlrIgFUrC5qYMTkpkJ7yoGKv/+L/8rxQ58RbMAzAPaRFvcOXYQkMzdrXdT9YZcR+D8GoCLsDGM8+QH1zP3Ac7F2AFTEgfbsEczC+30uuk2QO/Y7/CDPDsgLILv0y+DpsVZvwagIc89s593l7BgAEjh+jpFk9Her82f1WwNWg99ipi0TlXTeM1hvmdEDe3rUpmxmCILdUZvtBuezSCyR3DTaw5no65E/x24berA6c27mzAnY9KGsm2fsa5HkOCCaadcF53TwghIvBlAwszxiIWbMmhzQLRcgDJmzwenYbwbDcT0rEIxIgbEO0lfW3DDV99cx1H6yaLT5jQk7Dv5JUf0bjr2d11kjnAdGTPHMdGVudhRogI8YgCJYu13+EYFnABWoTcnkCtTJ6sBvR50qDY4jPoBxpVLCEHwPKyjtcjXGKmG2eshKgvsDPxoFrrHvwh4oCIP2zhCi5JExPzgmolJDmG8ONmkdCZ2PsXqEAT1WNB3fwXmQ/MEXgRwNoHvNEvRFr6GBax03WzuCxBBlcNgr9UjqFAgSu6zWoTMskciCsaXcU8QuMLaPj4/VUPBtCvsiwUgDUskcQBDeJMSiQtpW84mAgzGIorhFlMBloW9jKgEYwTzwZ5PftbgNgYeOMmaUqaEJHi5F7LXHtFaajqn7OZTqMgaJP7N87iwp0xkkPlZMXOT1TMbM6vL5PeEtwxy32IeuMXoPWEeD8touDaVsCdgGSMb0caLdbLEAgnM2wOgvZK8B0OCyXpTeAUz6fPb8ud2IOYux67S7jJkgIZWF61ut6BoYK/ydsCBkNM2fZqKpq1WgjWi7zQedPSmwwpBlRn6eMip2aD08Pew7MwLfKlCRYxNHD1WkURlmdcZfipHgeGXXvyXBgQFbLMjuigY+MtBtdwrOEQdYdnab8g3G0OFJdj40GmM6oKPsaaBid86EtzqPUZHVK02e2Ma0NufUdulwOdRgnIEtatzqhqO6kKgvAUS+KZutzW2BipXmRgRU+ObnmzSACjW8NIjskhP+t3QQIN3XdIAUbWUBYaDpQe0LL77pElRpoELtFDPsrVAVUXdz+v2nG9wOAITzDxkkIaPCpayGilp0l5kkCPwiWANqpBlEEUJugAIzGNptZnbidy+mPTY6TjkMGITjExNSqGrRp2q5opqMrTYNOgR+YLA54OMbKZwXGBhjlo3qG37IDEExbWQ2qPRT02pOqPQTGAuumYsZDKDi8cNHAaPiEDP50T4NGMRABYwDz1pNB7A180cDGgRqGpuahYB5tw1Qcfz4cTk4rUAF2odArRbTRqqPFn7PAyoimTYYSjTaiwyc/PqD92Tv3kk5dOiQTB86oo4AzjiEWhaDQIVm7nuWuQrAIIbhjIq/+Iu/sBoVyMzVDCqAfWgnXkqH1TYwS6LbJVCBcTr/7LNStxoVYbA/YlRQ51K/C6Biz+QeufTCC9S/pyKPyZeBsQHjZwiMikZDPr1xXerDJTl39lxkIIHJAyfkwP6DpO56ZhLBNZNlo2Fs2VZh0B1twzwKARx/ZsJnNAuwiOz73QaK3C8wRgXmPYK7aJezp9qdTTl4cIrrlzpRg1KGWwEVkH4CYaVWG5b68Ggk/aTZyQgAGHsCwAZBDJ0HDjRkAQPhuKXBiXAs4s92AlRolg6AqD8EUJHcQ3OAClGgotlclvGJMVlaWpSjR4/L2uq6AhWTk9LYXJUTp05KuTxO6SfIuP3Lv/w/8uKl4zI9PSXV+pT0y5OUZvrVm/8mnbUn8o8//6m896sPRHptuXBRgYqeVMlmwD19/OiRrK43IrYUgr5YP7nOVhEUF5mcGOfz3G5pUGJjQyUCP/v8cxmfGJdHjx+TQYXAOT7H/qDsq44cPXpQDk8dlqF+UTYbDXn37X+WV157QfbumxYQvyD9BEYFa8H0u/J49rEsri4RqGAtJtTDeLIgc7NzPDeKMAM4p8RTZYgBehSKZiHrKJBe4boPuT8sgnje6yN1BgBWVxrSbvWoEaxrKejfWtDbiyPiPNhLucZzD1Ow2hkVuwUqnFHhIIMXf8be4kEMnJ8slW6XwE+Ujdduc05q4B8Z8Ap2OFCBZxbnALMEn1FWTRQcxHMH6Sc8txivLEYFnhN9htNAxQb3ImV7AERRmj3O4+A91nuvUeH7NfqWBirAREP9wsePZzOBCrcfQqACNVVQowLXdHtDMxHbsrm+xlol2l8FKuDQKlCBoAKACgRrypzDLKYN1gyAn6YyKhAswr2F9BOuofKZAPB0FQmDg7rBqbSCtzVsswMV+Bvagz3CWRuU5whM1iRQodruaaCC5zZGha+vWwEVlXI1AVR4jQq/J34OjJ/bNSr9lMOoiNRhtOFe1DOMiQ3YkjtzD2KTLy+jPWcf2y7QvRtGhQd6gsbYr7vzLbbENbJK9fEqeT3JvrZLM+oeYqlejAluNyKDN2S3QEX2FbzWweCnfn7VM489uYEir5HtsSW8MNCB3LtjQcKwf2FAzp9L34c1eJrN88AxXiCbv5tcDm2zFDMknnMBUBF0qYcEiSjga/7sVvfN7mtUxNxs+hA08XXH+5crs5QjCaVAglp0zvDQWanZ2coqUCDAgfvtpqwHORXgjGsbpG/gbhkV+rjogHoQNFx3fY3mGmss+8zhtYlDIMWSk3Qv0eC01wQAQI61DkkYBJjhtxtdnKCAs+DQGG+XqSU4q9zBYfrK9Ms0aQnMegSPNQFIwXSurQjOsuCwJmvQxrZEHJXz0zmoAW8NVuO8SPpi8WrUVQAjo6x1KDxw7HMYa5QCHZqQ5bLK3OMMOIC/grkAHxg/oyQgY5G4z8LkCfTXngm1X1Qq2b9DBiHaZHLVZHaYP81AN8ewKwWXBA/WtXB5TAN67udzjrrUFJkdCgz5/ui/+z6LwDaSFXyuuD+PvmLP1/mOQstWz4BJKz3kDhnjQesrkokSJBti9WCgHGwc1mVQ8MPtNpdL4ndN+pt+pAFrrDsaADhu43EuWCFvZ774moR76+3X9Uvvpy63qPOBuiUKGOGF+cyC3van9PoFG8qBJmVJ6H3k9fE9q9tG5grs0H5PKpTsVL9bwTf9DH10dQKumQZ84W+MpyBR0ZhBGBMyNDh2seS2XjcGR/BdZVAoCOnMNpWe0iLiIVgb/h76ib6++XrkbIqnNSp2abQ9Pfy7MQL/9N/+MruhZij5h4kFIc+a/daAiqRKajIoMpgllNmcSFqJZkAC7FBnPbuxeYZjCLYkBixCV9Lf5M7vED6/4mOoa64b6LtzJMJr7xSo0PFTQzb75QV4g9obdqB+wzeKoEYFN3JIKmnAPWJUNBuZQAUKV643Nsi0WG5sJOhuuilqUA96/AjacvMCXQ+BnTZkpZDNrRkh2Ew9Ez90Htzg80wI76sqtsfjjWuRUVFBcEsNqhioQHBJDfioOBkDH6q36EF1DzxGBlBQhFqvi4JkCuA4vdrbDJ18aNlrEVfVvawPqywVN6AgeOAOOa6DAA42yPXVNcr1kFExNs5sgdGxMSnWKjTUELDg+PX6vBcIXOAnN1NmGao2uRfowvURGANbAvc7Air42CgFc3lhgUAFa1SgODZopoGR40DFIwAV+/er9NP0IQbPNONRZVnQRxgacHg869PH1I2cLKDC5cBYn8Jps/ZMrSwtU/ppGtJPx5VRUapUpRdKP1EfWzPNaThFBbI00wdggM4fr/2gIAEysAFUQDMeNSoOzhzW8WGNCmXBqPSTMTICMNZSyzW3pi/y6Y0bcv/rO/Iffvxj1qgolGODsQ8dTdbwMGZNBFQU2DZkdaM9zz77rFTrVd7zKBMmzJgtQLpcnyUyKiYn5aVLLxJg4v1ilhaeCKXwAoxpbDbls0+vy0i9TGkppxbDwKKOJp6XsTE1gqlBizmkmp7MfqFMVlC/JShsH+0ftk6mgQt/ZkPwImuNCp+z6DnPXMygrYtMXTXK8czMzs7J/fv3OJdnZvbI5MQ+2bfvgAwNIYjnLARf8DzImdRexrxQvVIYnUItdBQ2xrxWUAuTBw6XOaEcE6UTe2ZQ2tDksx6Mm7/3bqWDMMkxgCPi67kzKpzKj7usGVhp6af0NdJDGAd5LXMszAAMfk8DFeD4myuh257VqJh7/EAajSUZnxxlhvXRoydkfa0ht29/xWeqsbkmJ06fklJpXDqdEhkV//LP/5dcfO6oHDo0LbXRaekRqOjIh2/+m3TXZuUf/9PfyTvvvyu1alnOX3hJ6qP7pFfA2qX3gg5+Hw5BRwr9rqysLPHP4+MTlFQD00N1cyFNoEEIyBYhcH356hU5fOSIXLt+TX74gx/Ku+++K88995w8fPhQRkZHBDI9p08dlcnxSSn0irKxtiYfvP+v8tr3X5Q9e2ek3YajqUAm1moU9b53/55soCAzshM7XdlY35Cvv74jS4tLlHUaHq7K+NiEDNdRrHmITBOsxxo8L8jwMGpUVCLpJzCBMMextmJ/WVlZl3a7KwCu8QoZFXCEqGvLLMQmmQB4XgGkFIso/Ig1ri2tlhaX5H4amCS4zwQ5mAWGvRg1qLSYNpw3BSoqsrGxzoAFxhT7Nf6uTJV1rhkAKnAefAfHYZ5hPXGQAgFmyDsszC/IqgEV+/bvM51rXZtRUBzsB0g/4dz4HfWvsL95MW0HbN3mAYvH1xaXegqBClwfQIXvTQCe1tbXCB75Pri+nmRUKABQpgP6+PFj1skYGUEhdNSsUYkDXt+ycrn/DRWl1WxQKop9hmyFJULg/jQb62RU+BqLtmI8MC5DACS6Xem2OgxQuPQTAQwkMbCYtko/YVwxHjgP9ulSSf8W/ovswb4W+9Q8n9g+cm1uD9I5cMJr1GqWtWhWjtliaAcDJ6bhjO+iRkUs/aTAvhfT9mAV1mi0k/Zfz2pUEEADUGFZCdKXtbWlwRoVVlPF7Yi/+/P/sg1QEQfFo/Vri7rUu7XMc6V3vjWggqt3tgkf/DXaN8z92PYL4XfzHaAMKartzpzdVt/HHKjwZLTcoO83AjCyZZDyRy8HwnAJmKAMAoO9lvCx3QjEnw/6X5kEnIyMe9+Tfe/2QFheUkO6TSE4wTXYEq808Js8OmpTYjiCh8QBJQMGdF3xukeDo6GZ5W5zBqPhSVkMRMeFo/WZz56EmfUdPKBsEnZhC7wOgwelfb3dChDzQDyyoT0wrYlH2a9dz1k7UWgLOmDhckO8z5YNTjaYFxMKm0DpXKyZKlHl7fCgP9kGUXFo91s1AO/zyetVeGZ9vAto/Tq0AX6GB1e1foPWS8I5PLNeg/xa+4KST+bL43yQ6nFf2useUYXBC7pbwJa1KoK6lbhuq6k1tch4LINtuyrlaiXyywnSW/BZaw2of6nBYvOlYAPC16F/hiLEyqLQuYEMdmUHYAwYQHY/3hI+0AcNpMdzUgECPV8Mutp+6Mf5PaMz75I+9tPlxLz4twEJWs9B5Y4oHuCADX11tee1OLzK++IYrbugUkWwGRjLqGpSDa7rCRjqV2oftdaDyfiWyhoDsaQy9Vdipo4+3xoT8MTBiD1A2W4dZ4w52QEEynq0hQg4GlBAIIqJcVozT9kRCvgg+QIvl6dGHxNSxpjnENuwOhUOOvpSqQCnAZMlkyMzBqw+SwC2tI6qy2NyrqMmWVvlYZl0CKkn2m0KSpF7w+RKTdIlKGHzlPar3RfGo3z87NmIAEf2U8EsZU8oGIcX4ga0RU0iHONBW9EKxXONcDaPJQb6WhmuR5qQps/40xoVO9+Rnx75HRqB3QMVqaJA3tctrPoko0K/EBsLFr4Pvh9v/rFjEW8UGddXjyo56gnLIglUeOZ01m3aNVCRAkFCwzQNVGjAPzlgAyDMLubO7oAKjnoGWGE9TrAp3GTRO6coN7dwvgsz9GJGhYIJyqjYDKSfNhisYFFtAyrWTLfaNyOl6GuwTTMsjOZpdNAYrPBCTRo8ccMzAi1yxg4uC0xhLOYuJzQ6rDUqfMNyoMKzGCKjNiii7vcqMjINjPDr+9/9uzgXGRVWGEyPwz+lp2Jw25sqleWsBp0iTufVzUc3YpPR6HYJVKyvrMn46DhrUxRKRRmdmBQpqjSCBlKKJpsBZkVLC4oHsk/eFz8/64QYY0SNvLgeBDI+F+fnyc4Yrg1LxYPk2BhNXxfHzz1GMe1HsnfPXmbw7586zCAQDCMaOkHRdABcLtngQIW3xYEKakCiwLoxKjQi3Jf+kDIUMB/xc215TX7/yScyPT0jx04cIVBRhk4rTYQiA/dgK/QKaqgpUKH9xe/MQurAsItZND6VkKXy6w8+YMD/8NGjMj1zSPqU7xqi0dIFa6WpxbSj73v2KA1Ug8jAqLjxqdy5fVt+/OMfU/qJEW93SgAAmHGL4KMXUKWZ2+vJ1StX2P1nLzwrNRvTcN57lpzqwWqNijdffz0CKpB9TQM0Agy8GJlmW12/fpXFtM+dO6ta9SyQpg4FDMNavSZ7JiYj3U4E1chJgFHHwGw2UJFe39JOot/z7Y7Lcy492yd89NOgBjLRf/e738ny8qJcemFGhofHZLg6ySLMUqgoOwaUYUshy3Jok8+LAloIjmr9A2QdJXcON/DRLjp95jR6O8NgTfqz9HvfL+MxMLZOEOkIg1MKUtiVHIixGhXJvXd3WazpexC2ZwiANRMArOh6vyso5/xk9oE0NhdldLQuG82WTE0fkbXVNbkDoGJiXBrNdTkGoKI4Lr1eRdaWl+Vf//n/ltMn98qJE0dkdBJAxT5Z3+zL+2/8q7RXHspPf/qX8vpbv5Qjh2fk5DPPS70ORgWACjxPWoOp262J9KH9Pyu3bl2XffsPyMzhkzJUBLMI89rvl2aNIVi/tLQst27dZF2WO3fuyKVLl+T999+XF198Ub766iuyqvr9tpw9f0bKpYoU+kVZX1qS33z0C3nltYsyueeYaLkbBSrgUK6urcrs7GNptbrM7kOQHoDN119/TUdlZKQuw7UKr4k9CP9QFBtziwGSAmpU6O+Qp1JGhWYk1kdGpdXtyOrqGoEGABV4VnX+Klg5VC5KF+teX6S12cJqyMw61sMprEm/sCmCOisyzJoLnB8A0l3v1oAKr2+BvQr/vB6E15hwBkAIVOD6Lhk0MTERrbfU/jVHkmBFtSLVqmr3LjyZZ12JdrcjewFUVMrwYDmfAdjUh+uysrLG569Wq8r6xiqZJg5UeMCcu8NQgXJj/jzDDnFgBMdp8e8an2EADDgn2otzhjUq0DffT7UItgIPcM4fPX5IQGFsDAyYopSLKrXkL2dUqARAUx49ehhJXfm+jra0mpt0fJ1R4TUqCEogsCB97r8ALiBBUAIoYnrRraZm4bk9g/mF39FOlX4y9ivHUYMX+jOWd4qsUm78mqBACQ3bkzZW17gP8RrGqMhaJykJYfIfy4uLKjFiwA0Lw1LiIGaqenvQVsw/gIWQrWAyRASCdAWMilAq0j/DPcPxGLef/NnPv0Ex7WyFp92CFGpd59QI2AVQoWEtfWUrSWWHTH0u+X3cKhibmKCpN0EOVfyJ1+m2S0euVhS/3h48CS+TbFsMjOa1efd90WBb1mt7/y75rciuS9drzoKMtgNU0jfUQPUB8CnIuA/tynR/wnFJHxd+poFElzOKk9Fog2RNMo1m6+WiYbSbPeBmGxslB1zQHLdkXSw9rw6o69HDhtK6CG7bD0Jynv0fJfxZ43B+Z1OEn8F+JYsi+od9GYl1lrGdMfcZrMaaRQkbZTVoxry2mf6wSQJpZnkOIJb3zDPZJZkEQs/az8m1UiWLuAYY0MNcp1iUP46fOJPE2CSRDJYl1qmsjDB5DXa+3lItkMzsdgM6/H6H13OfzbPG0W4EWqn/D1qqCM8J/0rlprRmo7M2dJzg5mjyAlkOIvRFPfhLm9sKnRN0sBZ6oDf0uZUd2pdmWwF81hiMmBtq98BndPlmz/xnTQvb79Su0f2Q+6BJeznIgXHhOU1i0GsPaOBa7z39LmOWaLxAaxEmATaTEXZlqMRzoH46fLVQioiB8SB5gewBshT0oXMlAPTbgQtKZlrtMfrXBgTo3q3PPfsesgus1gLOiWvQf7HgOPoTSRd1NOEEQX6PzzjrweXFMLe0NkpHbULzp52Z4OwdX0qYLEeZM12HmFRjEsp47/OKc40JZ2A1mHwYa12UtbC63Tu9J16vkfBxxCJWUAfBfyQwKdMYSTX0961mB5IwHWjlOmHxPGVjATgyUMoKVTurxZM+w3nBui9k2DhDT+eKAmOamEnmMvzrIAZKNQWr/ULWhxcV93iJzz2rpeLjxvvKY3WN9bX0qfRTeqd8+v47PwI7ASoiNgWfrt2b8FtnsQzqxUb62tGlUkBD2ijKalICyQ6zBP3g4EsByJFryA58EAf4cyfBgGGacW0zR3yDzjtXOpCnC3+yUeGm7ptq8nxZdyKnTZa2rgbvFowKbAbdjjIqKP0U1KhoNBSwSAEV61YXIMp+RNA4ACqwwWBRx/ZDgwU1MEjT06CfB5dd29hBi7yxI1BhTAwvWFwplrixkmFQ1CKW6GsyI1ODNv4adMxV+icdbPX7gHOF0k9u5HjaL66HIDyLZIlQZ7taq9J5CAOjnjnP4mLlsqwuLcnywpKMjYwZUFGSsck9MlSGoRIDAg4ERICQbXzOXgkNL4xzZNQw08QKjhmjAkAFrg+gohoAFbFD2Gd9CgAV+/buk9rwsOyfUuknb4ePNccEhoCBKZzLnmFjDj8MQRpkGMNNZPGCEaJZ61FAADUGQqBiZkaOg1FxaEpKBlR4jQrUf4CMFYKUIVDh96jb1uBZ+Jzhd4A8v37/A5mYnJQjx47JzKHDClQYWNFtt5kpGwbH4/MkgYpPb3wqt2/elL/+67+WA1NTBJbYd2Yv9aUEA1ig79qJASAHKi5f4bHPXrggI2Oj0X32uen3GEZ5OQAqECB8+cWXmH3tMCWNS+BkBNCE2rI3AFSMViNGBe6NZgtpJgwexgN797F9bmjid6V3a8ZZOqDgQEq4LmUFHdLj7vNhJ5vrToAKjA2K2P72t7+RSmlDXnzxEsevWqvLyMgekUJNCgywa+QgvY76c5JuJwKcWsA4ijjoam77iTro6pN7v8Of6UDDVu9pnCakDwDDxdfN/e42QMVuxjp978L3RSq9YiSUCQcHtChdefL4gWxuLkl9tCbNVk8OTh+SlZVVuRsAFcdPnyajotctC4Kbb/zif8ihmbqcPXOcQEW/ekAarSF5/41/k9XZW/LDH16Sjz/5jVw4f06Onzovleo+BSpY40V3xV6vJv3epnx184p89dVn8sKlS3Jw+rj0RVln8Uv1dxHsvXfvPrPRMe99rcJ7SBDhJ5gPyJw/efoYA9v97pCsLS3Ixx/9Ul79wQsyOXGUz0KvD6q9SKfXkfn5J7KwMC/wNxFZIFASAAAgAElEQVSEBYgPhs+DBw84J8CiGAGou39fVNQZ4G4EVKCYtkk6gYmCOQdHG04R/t7qdMm0AFABVoY6+JqFSacNBQix2kIGYbMtRTzIYEp1W7K4fE+6vU3Zu3dKKuU90kV9DXAPmUWm2foOLjNbz2QevMgznitnRYRABdZXD7i7XKEzKvAZpSIMKAZDgCyBak3aBCqeyOrKKuveAKiAY8rBY1HxUbL+liJGRY2MChS/9ppTHuDA8ViiUaMiZkbEQAXGHm1DwANyUpAmJLsMQMX6KmUnPJDvQIX3lUKCHB/Iej1igoYDFaUhDcb4KwQqup1WLlCBWicopg1HGn0IpZ9wD3G/MW4OZrntg6AbsirRnyygAtJP/ownsvwieazYhozWN/4JwKPJEfaFzKEkUOE2tX9fnykkLmBthQ2/uLDI/TkGKgDwx+tr2B5lpilQ4bJVaaDCpdC8nb6/+PF/86Ofs4ZJVjFtmg4Jk38bPyZYs9P7UJYtrsdkezp5wcyB5Cq/kCc9ZGyAeUH7NFDB1jCTKWcXzXHKsty7UA7I4ssWPNP9LZ0jtt2+nR/P/+aAR2ib6xjF59oJ0JHFNg+DSelhVEAn+KsFseMMgdQo8NBk/7YrUh7aVFk2SXqcs/q5Xd+xa2dOEdO20jEIr5QzxxlJ1yC4B/w8eSVrTDzwPzAqmhodvfIAFwbzwtoU9o3EfcyZTg48RJ6vgbORhKknLLllZ2tlCGJ4AefdAhUIxiOYzhXWpHd86cC4ads06IiBYIFiAgsI1rq0kT5+Dsp7YBnnUZkdA6PCcUwzgGzuYg46w4ZhWg9rGECDfYbZ+Q4mQLLJpX8syz+SRLaCwt4PDZTbGqQITyQb5XtykiUz+Mz6vUJAnYAA6iUYOIAxUTmqIWVeGuMgSq80ZgKy/PXMGsuIgtEW26Cd7sCQsfQoTWW1Fsi8NQaF/wQARBvGamjp5E89SXY/4UY5S5333K7BcTL1Bvfx06Be9AzlLOReuJzMRQvoJ4uH+5hyB1Tv2tg6lL3ye2jzDWOFOQBwCYwWxCM8eE6JrSFlTRCDMnBNwYSSSn6RyZGROGzrSMhEc3AR9xFzjMF62M0APYa1loP6lyqdhGcBoEMInGlumSYnsW9IkCqjELYyTbh+GINGGR8q2UQgxAqCO9iCZjvDxmWxaL24P2dslhCk8Boo+l2r2RklA6r9jJhV3otxD0vkQD/IiDKmrLMwor3dQnHedpwzAnqDRfopULGdBfL08+/cCPzTf/txZpvdQIhtMV2EtzHvs8+V/5jaIhCeNc6+SF47PCa9IWRcIAAqYsci/J5mK2qfQg8md0nJkIvKb1OBFnx687IxZMcyTd/ce/HNgIr0HQs3Lb9UTh/YRqcAOhNEg9fuBzC4zYJIJv20C6AChoAHxlk7woAKZgNnABXcnExPHt/zIsgeUNoKrGAAzTYnrwMA59lZBAj+OCUwysbwgKPalNErdAgREEI7/N648RUCFa45yI3M2qC3XguabW40CFQgIA7DARm2lZoW7PTz+PeYAVqtyvLikizPL8pofVRGxycIXozt2SPFMoLxMSsgZFVwUwtADO+QnzsEKtzwVecP1OI2JTnIqKjWyKhgXyklZJlG/V4CqABAcWDmSKJQ6XZABWcrM3308XANyHZDwS8HKgTgkdVM6Xf7MaNiZkZOnDDpp2pVuqy9PcQi1TgXi2alGBUOVPQtGJYFVHz43vvUjQdQcejwETIhYKS5bim0x7cEKuyxu3blKhkVBCoOHqTGOIePxe2SjIqIqWKfX7l8hd2/8NxzEVDhbcX6pcwm9LCfACoQIHzl5e8RMCLEw+wiJQ/w+L6wmPb1awAqlFHh2S5O0SYw2O+x9gmCQMO1qlTKFZWAIrMErIRBRsV2AGK8x2QXNw3vRZ7DnQVUhM9rmJmFbOZPPv5QRkZL8uzF0yyMXK2Oyejwfijg67oWBNLSi3H4POK8nv2ubIrYGE0DFcpCS2YV+vu8v6evnTwurn/iGYvpPrtTppsc/nnWUdJo3iqQkW5b/v3oS5pRgZVhqN+RuUf3CVQMj0BmryAHpmZkeXklBipa63L89DNSNqBiYf6JvPvm/5S9e4py4cIpGRk/KIXhKWm0S/LBG7+QpYdfyvTUuMwuPJZLLzwnJ05dkOrwPun1USxenXt18AE8b8rl330g7fa6vPy9V6VcGZd+AUBFmAUJqnhbGhubcvPmLWZn379/X86ePSs3btwgcHf37l0+/wAZjh6dlulDB1mfoN8tyMrigvzu49fl+z+4JKNjh1ifAmANAcBWU+7fv0tZJCwvuA5Ae5x/YWGBew5YASN1ABX7I6ACALrKEalUDhgVeK2tbkRABeZfrT4i7a4CFZB+AlCh+5dpccNigZ6ubditzU0pIVuz3ZKlhVm5/+hLGRkdlgMHjkq1tk+GimAYwimsRFmfaAOeYwTw8Tv2M2UixNJP+F3BEqXRu/QT2uI1prKACg8wO1ABxxiMipXllQGgQhlMowQWUKMCrD/IZjlQ4TWnCNjC9CJbIK5RgfFD8N8ZFZjb6AccXwAVkL1SoAKJFWtSKitYgz6jb2RLUKqqkihwOTcHoKLNwua6HhqjyB7IEKjoddsEKrwNbkvQnrFCpF6gFCwRnBdzAY4rggNeZyUCTKwgJoA29AfHYl4AnFFGBZIwlDWKz0NgIG3TpPc9yiQW+sq8Qc2MtXWi27A/oloTls0YBVNcFgZZnd2e1ndJARWuiIHrhYkRClRoHRWVcgJjRDMSsWeDUYFghQNnHpiOAK9yWZ4CFaF9vzWIkLfuRz5RsE3EwWpNqIDdx/kSZZjn+UzZf/9DARW6z/rabqHJgJ1AGzwHVckdjxzQKA58ah/DwHvuaKQS10KgIu87oY3kz3H+sbEZkgW8DNgUKr6S+HPkDSpKEvUtamsOGKdj4AWZ9SxbARXRmJn/4O/VNcoO7FE+xgoGc13IY2pYj/LGIH2vY0lmY+IEIK5fg2t1FNQ12VRjEWTdj1wAI8i21q4qCKEJFjpu7ks484G1rlCYlwWBlRkDAJ81p4YKlM5x0MOBjgTYE4XpB6M3DFEE7BlnBpj7r0WSKb2sTAoGpU1PP2bFaC0KZKczmmIJZjoJ1H5wsAN9xHv6FmCX2JyJx1DvPYECk0LGe98r6d9abQCtsRfX8vCsdJe/4h4TJfeEqE3MsqGcK6SQwSzoIyESe6lKWfFF2R+9Jwx0G0PFi0BjfMCsTNqU2m+Otkn4RtJTJhHU6iirxGWh1Z+2moQ+GFYHgtcKxiKcbwyUI6kvYChErFqTuYqfY/NDrGYD7wNkmAGW8PwqPYR5pfLamqyGkcNxTCopl2g3KciiSUEErszGIDPSi5sEDVWr3P75mmrf4zSxZ0v9f5fwYlGNKIGQ0qJIXCGYgSQZLdCNe4YXbDYkzDoAA3tM7SaVpdJnWJNReQzBOE1KcltEmcI9SkLpcxn7pmRoEIjV4vVkZhjQpMuYslXDF9ePrDWTdVEgvepFvtEmlbjC/cR8Qx8hVRYCgVwvvIi7XUhL9MTP9lOgImtFfvq37/QI5AEVedlBiaD+Tnueg24ks3PUVNE1TDeVbwOo0CZ6AxyZwIJtFPcdAhWO0sddTncq+f6PAajwDT5tBAxQFKMDQsAmBCrsALUSDKhQxzcJVED6yRgVmxuyvgFGBaQU1iSsUdEwpkHSUdWCUr2+6nhTvsid2a7VFWBhMC9QqwUn3fn2QEK6z9ycsKmac4UNnaG7wG5xnWpnVRDlNopnl6JRMeUzDN4xs9UMR9o0tkllARW+iTltlBmL3Z40AVQ0mwQqPNO/OlwhuwKbpm9KOCdpg2RULMvS/AKBivGJPVIolWRi714plNRgCNsRUikdKPC++W2n0WEa0/gZficNVNQqCFKXVYfUhFY8bRxsCmdUQGrowPQRZv16sMaDDKTL0rAwwMOz9KMaHWoMUAMSwS6COU1tLooVI5jM+6cBkY3VDfnkd7+TqelpMiqmDk9LCXrdlPrSYDrnkgEVbgTT8OwAMOsweOf3OQIAoGHZbAqACkg/HTtxUg4dPkzpC5yboB1kYzYbqgMfZNNrY9U087l249p1+erLL+VvfvITOUhGhRYlJf0YxpPpyoJOTSDEGQudjly5fJmng15+fWyUBpvTtKmfCWPZigp6kTzUqICMzPdeepmZ22gvgpY0uFiET31RBypGR0py/vz5yClwiizuFwKiSwsL7NWz58/LyDAC+2CBFKVQRBHXJBPBA0nhHNtuuwjHPT2W7ryFx0TOS37kIwIIfI7PPnwkn1z+QMb2lOTc+ZNSKJRkpLpPRob3M8AcPj9Z7Q1BCBi7eE5hMPteFX7u3yd7xZ3+HMDCjw0BDM6gLGecf8d80yKSflx4jqjtLOrNXg0cl/5eur9bgRjp7w5Bsi+SftKVodjvyvzsQ2k0FqVWr5BtAEYFAql3b9+W8bFRSj+dOHNGikOjZFQsLS7I+2//swzXmnLp0jkZmTgohdqUbHYqBCoWH9yUZ04dkvmlOTl2/JA8c+6i1GpgVAyr9FOBgy3dHrKqVuRX770uM4f2y7lzzxHM6Bc0GE9MyjL+IMm0trYht259xTUX9UwuXLggH3/8sfzpn/6JfPTRb+T06dOyvLQoF54/J/WRKrO/waiYf/xQrl97T1597ZKMjExJr485BEdcZHl1WR48uM8APop2A6hA8BbAB+azBterUh+uyoEDB6IANtZfX/sRpIbkEY7fWN+MgAo87/XRMRYORFAbFHVIP+FWq/Ot2XpDJQAz6pC1mxtSLfRkaemJ3Ln9uUixJcdPnJRKba/0+yMyVKpy/y2XquqIGqPCnVd1njrGRKio5m+lynXcC5brmupFCXsRUIF1COfkWkIZCK2xg4A61jIwKrDWzs/Ny9LiIoHR/QcPRIwKHIuaMAAKQqBibX2VwALGEudyjWdff1EYWzP+imwjrutgAMAXnI9Z+CXU1EA/1iOggtlqoswLBoes+Df2FAb++z0BUIFrjo+PqjMcMZhim0EZhSr9BBkwb4OvFRhXgEjQdfYaFQ5UeDFtBCRCoMLHD+1gjQrT8saaDfYPJaNY+0GZov7PA1pZ9kq4tgKogFvOAEi/T7lJ/ESGZQF1TixgpAEdy6aG9AeCFEXUVTKgAgkSlpVIQFejNwzSuMymJlQoUIG9SIEKnR8hUOFyXN5OBynwHuP2RwtUbBHczdwTt2RUZO+iihskE5HUjs0+Pndtt5yk0D52oILfMaftDwNU5FkI2YHr9B4U2gPheITf/vaAiqRHGF1jC1skLbO0E6DC+5hlVwzu12G+xPZQhYbQBqWLssAKN2dzz2q5Gi4No9ZvhuRT2GhnoWgno0/yxkWLNGvw0pPC3P+LbJ/U+fNnVMacsqC9+39um/t71+6Pih8bsyDrGsjsznuxQDH8UEjHWra4Bu0twcDsc3xfM/FR60HBaLxRWSoLlNoerYFw3bN9rgyCFQ4gxS0LgQoySjz2YqFPXBPyNrgm9if6DTBuwOhgnQPNZuc+ALKmyeoiQMyVntJ8Zcpe8lxd9S9xHO+h+U3Jx0ZVEzxRIATr4Ico214Dz57F7xn0+A6C1S5dycA1g9vBzCXjVNsK21z3H6uDAIZG0dn8GkiOkiph/5gsdYJ6gkFML7SQGrLYAOtZkf2jwAXvkckuRnON9Ty0LgrGGv41WZuIldA3HKwfqgPsSQgWMzP/X59qAxp5X6NtWueQ1Rh0oETrUunc8n0Z94ngAKS7TBrZbSeAYwjmu43IWJCBB1nznp5wIHnm/iHtKJ/D9tOvi7kCtQ4AdLAP1G5EnEj75RJQKilmtQmZpaJsq3j+a8KD1lADY9UlMPUZ0mLpYeJEzHhyB0vlz1VKinaRMSV8DnJ4jS1DBopJj+pzEMcao7EhwKJ2sANhXh9TC6HHiaUem9H5EwAnEYMIV4gzap8CFblL79MPvqsjkA9UJHb82Ij4JpyKHGNZTxp/GBvPfwigQq9DY5Z20W6BivQdtvOlQZBwJRowWk1OJ9VvTYN3vHlwJoWbWfKupMCRQHJkoLXmIA6ePTxH+DuCqDBEQoOLodMUUOHST5B/alFGBgH1DQMqGpsoTrnOIIHXqNg0p9sXYA+g05Dptbnh0XiwzAw4vUppVaDCX1pkW/WZWWQoKIodBuvTQAU3kTDBwgxfBAW0OKjqP7M9Emu7hoEFBqktK92PDX/iGs788CABvq/IvloNaLczKjRrpW2FT/sMSLnutgMH1PYuFmV9ZVUWn8zLWH1MJvbEQAWmkWfEOTCitFU17HEeDwCE88AdPA9M47go0FzA2LdlcWGeBWehdVpDNj0yEiwjiCZOr0eQIguo8PvrgQcCVKSXqsEdGtj8HRktzBRKAhUaDE/WqEAUbn1lXYGKqWk5duKoTB+ekTKACkpYQUJMM068RkUSqNAaFZ1WM+5zADgAQPrg3fdlYmJcTp4+LTNgVDDgUuRPFMKCvrgXVUsGAOyZNvYzgIqbn38uP/nbv5WpmWkFKjh2ClSUbW7jGeI1WCQLurBtufz73/P9xRdekPooCpSrxAiDkaDOdtQR4LiaMfzOW2/J6MiovPzSSwzksb1mGMLX0LYWCCLeuHZV6vWSPPusAhVsl0mhYZ7CQXh4/z7n7J/88IeUAENgURkVXoR3cKHPAhby9so0UBEe5w7Ybs7nfQjvSbdTkMezt+WTyx/Kvv2jcvbMM9LvFGV8bJ/U6nu0ALYb+wmppWSr3YnCMwoHjuoBQT2ZZNtjwCENPKQDRmFQMav9el6lOGs9BvtLYq/R+6qHqmPkQIWfM/t7eXcm++/hfj0ERo8BFXp1SD91ZGHuEYtpV2oawD84fTgCKlAwerO5ZkDFGIGKhfl5+c2Hv5QhWZGLl87IxN4ZKQxPS6tbkfd++QtZm7sjf/kXP5Qvb30u4+NVOXP+klRrexNABXb4Tg8MhHn56MM35fmLz8rMzFHp9Yal168S7PQXAvxweBD8vnv3nrEHNgSSafPz83Lo0CHWk5iZmZFupy3PXjgjiNNiXBFYfXT3jnzx+Ufy2vcvyfDwQWNTKMX88dxjefJkTms3NVDLpsXiyyiojH1GweiqDNdqcvDgfu45ni3PTHpzxGvDda5Rm40WQQuMLvYKABUtFtNeocQCGBVcE0zyhUGQMpgsVpSvvSGdxrLc/vJT2WyuyOGj03Lo6HHZaMARrRHU6PRbUi1rFn4IVGDvcfaZSiZVLMtOg+shUOFMgJBRgb66s+jSUOgf9jk4ohFQMQuprAUGTPZPHYyAiohRAaBiaSViVKysLhNY0OewotR5ZhLqXgEGi18vrFGBtilQAVZLjYwKABWUqdxQRgX2JpzHMwgJVKC4tSVL4BkEQwJrv0s/QWowfGkQRIEKSARiPvg9xnG+92EPQQKAM1UUfNLij75uO1MFf/MgPTMKW22tWVKv8zv4Lvd6JHuA7ZYqpu3XTWf/+fqFJZ11XApaXwIvr1EBSQZ9AIwhaqwTDzh0uXfrHFxcWOD3+S9ik8YZki7hoHaAAxWNSPopthc6UY0Ktxf4bBiQgZ8Yt7/6k3/845R++gMDFZ4FHQf0PO6bH+BP7wNbrfy+q+s8cqypoIRxCwzl7BC72lC+KdMi9o80mKTv40v7uBCu3zWjQs+TDhNqbm08FrrXekAwY9zN5g8HZKdAhX/HE1PSNkN0TldNCn2bLeYenu905v+ABafOcnCJ7DkVti1kKGwLl6QYLzpMdo3UpXytdN8mBBIieyb6xYK0283A1KTjHA/YDVzXrL4B91XzpVT+xiWRBy+SB1SQ/WxBfAVhbb+yc4d6+7SiaN8XuEdqcW+diSxejILT8Amt2K8yGToRI3pg7A105hAH46xBWGVLhfYps/htfDz5AfeHrBZmvutsYbIengUDT8gyIEu8zyA7a0OybSovzCSKbpfsSASiE/PL7rn7U/HtVOYDXg6C0N+2ehsKlqid7Rn0TA6wuACfTWeABTEbPkupeea5BmSxWPH5brsjwyN17rWe8U65JbZB5bkSCaB0xrXNZN4HBeMjVrsl42qdP7BPVdrRweCojkf4TKSmGsEuKwTu44xDIrZR4MuFa7f32xPMWNuCyWtx/Qg9j9YcwX8u2en7Lp9Hl/syVr9KEQ2CnwpUxLc69DHRFthIChwpUx22jtsnGvtR9geOw/1FcpjKbqPWpI4vr8u8CQVcYsBAk2DhV8NvJZhlIAFt6a4CW2iTFiHXpBQFQWO2QgS8cuFWFQPuDVE9N7yLn2+0S+9DcmroXmE3sg9hBY2BaB1RfZ7wIsCG+W5yWpTUDJgn0VTgc+11ZEWeAhXbLfpPP//OjcD/+d+zpZ+SWfe26W8hebplx/PSelKLuxpg8a7x72dUeKtikMLXiH8fUBGbc3DDki9LLWGWWbgD2neigj3JtiVWrtQZY0M8+UF+jQrX7Eu1LPM+eF/SgAU2J2zASqvT2xIU044CngoSYLGnLEQAVIBNgX9rG+uysR4DFU0aEwYwGKXSgwLOqMB71qhA1oZlcmYBFW60euABCz7ZGKYDyiB8ilHBngS3xgMyONazJjWjFSrrWoMizO7w+4H4HxF5C2g4UOEOPwO81k9e0xxrGnhA5w2o2Gw0jF6LMdEAAbe8QoFBFATNEIhBEKVUqShQMTfPIPTE5F4ZKpdlct8+aqJb2bcoaKoGotJoEeBgBmspKU/hsyQNVGgbYGy2GHQgUAFNb2ZrOlBhc63Xk0cPHyaAioOHjjF4gmuHGZLbARWqk24UYWias45HUwPrCDKymLaCZgAqUEwbQAVYCidOHpfpQzNShgwGNVGZz2kBdQBhWqPCQRLKGgVAhY+7/8T9++Cd92RyckJOPfMMgYo+gQotqA1DG9mw1MsdyLDS9YwJNyIsiP3lZw5UzLDoqDtmNMJgsIjWjDDlOs30aLfl958AqOjLpRdfNKAChpQaljzGiqYplVyNlnfffpvFZ1/53vcEDBcyKow5kwYqrl+7IiP1MoEKNxDdacE8bXbacu/rO5T/+qu/+isGV1H8VinpkN1JrrHR6hYUMwzHNmu/8OdqcByTer67BSsS1yrAwG3KnTs35fInH8nJE4fl5Klj7NfE5FGpDSMrPX7+8vY1HyOV6RnOBSo8CTUrWMhlNQwCBOyJvL/7YrwVUJEIZKQYFVnXzOtjbkBk4At9yQIqIP20+MSAiiqAvbLsPzgjyysrcu/2bQFQ0dhckxPPmPRTryJzs4/l6icfSKc9J8+ePy77po9IoX5I2t2avPvLX0hz4aH8w89+Ir/53YcEKsCoKFf3SL8wDNOeexaACjCHHjy4LTc/vyzff+1VGRmZkG4f0jioAaSOpTomXeriP3r4WBYWFrlej42NMlh+/Phx+fLLL8l2wNp74jhq1BwQyuL0sLaU5e7Nm3L79icEKmq1A/ASCFasrG7IvQd3BRn9rVZTWk1kuq9S9gkBcqznYBkg8DtaH2aNCrw8m9yD0XB0wUpDsLzV7CjgKKrNzL+3OrK8sszMwInxSQOltNaE1guoCOvzYY1rrsrdr67LwtwDmTq4R06cOi7l2risbaBoY12BikJTyq51bI441kpK76EQZqvF9mPeO3MC+y3GhzrDJvOA9qtzuMk9HH3NAipYJ6pcZoBZGRVPKDOIO3SAQEVJ+syuLKr0U7kii4srvM7wcE0AVGCMoxoVBlToHqxAhUpSlWRtbZ1OMNqWBipQoyIEKsoVZfuxDyZ14LaBHot70JYHD+/xXAAquMdtAVQ0mw2ZfzIX1ZmI7Qgtph0CFQo+dVWSEns4ZSm0uKXLOvkahPoqIVCxHaPCbRFfR31ddruFAUAJgIqgRgXuF4CKXj8GCuiQU1IB9keXGD7uOdhDWwEVvmcp6KJABcY6TKjQvW0QqAhBCk/C+PEP/+O3B1RENm/e6pi5g+3m4GxJCF2g1f7b1dmCQIVj1Ftl9+/q3HawZeaGHkNO+XD7Qh5Qktez7OO1G1mfeXAyTmj2fdZdnZ3uYXnH+RAOAhXmqxrz1W2WMACcHuIBmaUgWJW7BwcZ7joKW7EU/Ma7lZA3/vq5+gpJnztqRzh3eIgH/rPPGdlsQVCOMmHbvBLBdJ/3wdfCz1nk2oLTHjrIukYITGVePgG8JIEYH2P/ngfwCX5bf1gI2YP1OU9pt29+c84ywTZacgvBClgtTChxVoXboLHskQYyNdvfJWA8iEugICiaHrU/EU9RhqD+F8QnonkYK1pEwAXl/jQpgQHlcokFtV1eSDPcrb6hurXsF5MkCCzAjytRUhHSitg/cG2cgzZYYp4l54sm2MRgvr3hXuhBeZWUio8JfRdvc7lStuRU77MDLHGcxPc+JoahyDUKTBu4zgLdiEFYbU3KHzIgrfUxFDtKxXr4Vtdk9sM+5p7LhB5jYdjzguPQXiYqUE5bfWBtA9i72QydaIwMrPL566wDB5PcD2HPCTDY2BrYRFvEACRcD3M8yvi3xZRxBNQFQb/d3wvn9xbAXXqlCYEKnJfMAmMEAezwxDvs7bDfNMaixbaVSaES5LAL6cOjCDgUGkoohq71KVgI21gwEYjDNhrjwhg/zhbxhFA+ml4vxje4YE/1NcnrlXj8RwEGnwexP6xgWWohsMMYv6LygwIfXGPsnvgYEdzzIutWCJx1biKfGyBT7Es+BSq223Wefv6dG4FcoCKy9OItL9G58HlM/J56IndhbSeAigRbittwcPkdXCNgTJhwv+5zCdNM3yVrVPi5A4srfVf93FzQtJBsfG7LLUmALkF7E0BF2I98qzUfqAgvHBfC8mKhtlRGtTJCxzRucWKnid/w/nvhYs86sE22p9A4DRQGPsGmUEmHnQIVjp6HWZtqD3dpENB5tQ01BiqgG42MRTc0VCOQoAYQ6VY7koNCpqYv7g5UUHfRMlJCoCJ9exkEYQByhFn4TtN0IKCnRJAAACAASURBVCIyhE36yY2jMICKjdQzUN2o4/VNi9KBigZkjRqNSPqJFFEmssTZLTDupqenlVVSKsn6yooszi1oMe3JSeqQ75+e4t1qtjSg7xs/7pMWH9Nimwh0OWPE++1ORghUuIHo0k8EKjaUUVE1IAj3CwqWCEbgHgGowD8U00ZgfApARZ70U0GDciGFOwKDHKgwLdJOs5UAKkLpJwAVq0urBCoOHJySU6dPEKiA9NMAUFFUfUoHbjQ7QwEzMCriPquB6ZkX77/9LoGK02fOyOEjR5XCymLaCiJA+skNRp8LOrZqnjlQcfn3l+XLzz+Tn/zt3/F+DpUBGBloFeiQIiiIcVUoRuncv//t7/gTRYFHJ8ajmi6e2eXXpxFvzwcYFXgOXv3eK1pMOyjAN8iouCKjo1UCFaS2W2Yi56EV+P7q1i1ZWV6WP/nBD+Xo0SM0rClHBh30FCDhcyt8NqJAWM4umQYIwuBB6LSE5x5c0/K3YPSDznlXDfUvv7ghN67/Tp69cEKOHJmS9Y2y7N8/zexuzS7LoOwGp0f7tE4FZF80IycbZPFnOX6uo101FUzSLB53UpO1LeLx0BoVYeZSEthwuNIy/3mxONSSBkHyRszXoLzP47HvSyFiVOj6DKE1ABULcw9lc3NZSpUipYX27Z+SlVUEzG/L2FhdGs01OXbqGalWJsmomHv8SD7/9GNprD2SZ545JAcPH5NifUY63WF5/803ZGPhvvzDT/9GPvr4AxmfrMmZsy9IqTKpQEUBzB6VfuoXevLpjcuyujwrr732ihRYm6ImvT7qqXjWrQIVYBTd+fqu7R8NOXLksFy7fk1ee/VVeeutN+WVV16R27dvyyuvfE9GRvT7GM9ioSxfffGZ3LtzTb7/w5ekUt0rUkDx4pI8nntCJgYYggjsg/Ew+3hO7t27x3UFDC0E7xFsR5B9/z7IL+magzVRGRVDrE+Az9FG7G8j9VHL0OtJbXhYNlttAj9wTCH9pBmLCEhoAe2hIWhMd6XQ78mDr7+Qu1/dkMnJupw7d0ZlfIp12WhUpN0Fs6EsHUGNALWLMBdB+4fT6sF6PO/4XbV8k8W0dS1Qx9GBCq9RAUaFAkPtiOGA9yxkTemnqrQ2FajAXpMHVKSln1YBVASMCl/bHajQ+h1t7rvra2sK1gPEjhgVKv2UBirAkoIkAMYgLf0E9gUBmU5L7t27w3EYH0eNihKB8ehlQSXf55qb6wTAvCB2CFRgD6kamxPXhDwazqvAgALMLv2UBiqam5rgALYNgicAKlhQulwhABDaEuE6mgYqfP+lrAcTVEw/PSH9BFBa9Z0dLPDsQ8oPglEB6adeNwFU4FrcCywbkfrcBprreUoRUOGsVv8OAKGV1UXKPtDW83pjwe+wab5VRkVk0WesfrkAwPaB2fBsudnmWwAVeVcI9x3Pbk8mSuXvizv+JGRUGOMzplgMniUfJPh2gAqdv+7RqQemcx3JG8n2bAdY8HtObM8YkHSL6WOZeRA+R24vDZwi0irXBLC4dpRlLPPG4n+Wxc5uJaV4Iqggd/6lO731ncUe6b5iZFPZLwnN/SCQnWsLWCA/DSzsdG5F3zPde3eqw/O5JDD+FjPnBoGGPNsq+juH2kcz/L7d0GB8aQenABKC1M4isKBiop+QWszIKtfLapCdn9sainWzTG3/mCHtzCDtKxjxaheEdTk0gBnr5eP89B+9vkLQTz4dribhUw12jBUajtZ6BnI1kxz+KtigABp8LcbfsR77Xu4JaLBv1K4S2guMnpANrlny8Bsbm5vcZzWpyyVJg/hLMO4OuvgeQ7/Nixnrox7tH8qyg7Sigh98b4APvk+b2nwx2vQaiTZGjD52GntQOx22KuR3vUYiCziDwVIAwx/Z/GXeB9o/UCxA4oqeQKcBzm1ABX1/z9BHzASBZqsVyPsJlonVSYDf5bEC9I/zJPAHsp4lZ+RonUK1fXFPyGixexA/Dxrb5jyz5EXcK8wvJJq6DBH6ClsGwBj2YtwLggVDUGVQnxlsHth5rthAtg9AxC1Y6JECg4G7BGwMQfGkEIw7zunF0SN2gakroC84BgkrtE9NMcJ/x1huNDY0mWNIbQXEP2CHjtRHTIq0T9uIEsiURwVQMMT+su6JJZSyaTZ4Hkvz55LKBIg9mY2u/qKup17gOgZ0svc7ynzBVje5NgBqzuIgo9XWBwe7InAHIKD1m+Md1Y3VmN1ToGKnu87T474zIxADFWEwXeVIbM1NPKr6R+9ehmEUxfcDsdNdgBWDzIIcgCK02AmSppaUKLbuFGVtuJu1ubU2Igs3CVTQqYwuEeTX6G5gw6KB/GhjSAypvon34vSgaFBz16/kbdNrpO9YRP/b6uzZN2kwMynO3MIG54W+FKhoSRMFtSH91NhgcIWMivU1vl/f2OD7NhDzgFGBjcG1mZkpbIMEcwMbKjYrlT1CcVCMPQK8auh0Ok2i6DQY+iqTgw0Hkj0uBYVMDi/qxY3F609YFjokeABckBZuBoezAOpjygjwf25A0VAzrUOMKgIhTivXApgFgewVgi+k8EKbc6jM40CRJRmg22OhTjAqUOtAs/vbdPLRlDD4DYBhbHycQQsUtlyYm2eG6djEhJRqNdl38CCNCARVPODlRpprTuI9DA+cKy2h4JshfoZsFIYsOi1ZWViUxto6M/SRYYMgjorP2HPR7xOkeHDvPjOQR0ZHWUwbYxFmSLpBQuMsB6gArZ6FNM2QQY0KsDloTCMOVHRDUGtUgFHx8W8+lumZGTl24pgcOnKEtGKawAiOwGChYWr1KMxI86AaQTOTTvLAuv/EfHr37XdkcmJCzp47J0ePHVMDHIaE0Z4x5m5QhmAVf+d8Uofg2tVr8vlnn8nf//3fy9TUlNGCld7tgB0CjsjAFq93YqyiT377W2aNvPjSSzI8OsL5zvGhtq0XxmYerBouvZ689eabZN289sorGvi0TCway5YpgiJ4CIBevXxZxkar8tyFC/aMCeWe3FXGcbdu3ZLlxUW5ePF5OX3yBA15BOuQRQwHRDU2rRK6puWqU24Gc+jQJwEdXZfSwQQP5GUF/8OVbCuwIhGU9/lqq2Rrc0NufHpV7t65Lc89e04O7p/k8zM9fVSGijXKQEHACIHfrMxD3DPM7ZERPBNqFIfX83apJiqmgQdS4jU07Ic/g9H+EWb+eWZWvLskFvMk+ID7Zjc4kH6KDN3cQEc+w4NrXKCTG7bVXf4OMwP5UMhQH9n1XZmffyzNJgLEqA9RkanpI7K6tiK3v/xMxscRaF+XU6eelWJxj7S7RZmbvSOfffob6XWaMnNwUo4cPizV4RnpFmryzjuvy8LsLfk//us/yHvvvCV7p/fJ6bMXFaiQutaHwD6NZ6LXk/fe/zfZf3Bcnr1wUXpdrAdag6SLMTHHDkW0cc9v377L+Yx9anx8TBYW5uX40cPy+eefy9lnTsv8/BN5+eUXLVjgsmx9+fzG72XxyX155dVXpFAZk34Bur49eXD/Ib/TbDW4L26sN+XBgweyuLgg1UpZ9u6ZlLFRZVUUq2XZu3cvwQwFkaEHXVNnu1Qi66K52WI9Cjhb2OeQVQYQsonC2EvL7DeYd8oW04x3HFcpdaTXXpXZ+7flq1tfMiB85ux5mThwSPp97KNlaTSw5xaliGxJZKNVbZzcmTWqPK7BZIQUUIE9BXJDKDaOAD/2ajiKON7XRowpniGsNXDG0Y5Kuco9C32tViv8DLJYT+Zn6YDu37+Xc073QQU1atVhWV1FcesSmUwrK0uyvrHOsQDwEppQmO9LS0tR9p9KPYG9YYyKDa2HMDysbAjo/EJGaqMB5kXMqAArAy9KRFFSCYzCgrRbTbl392syeEZHsacCfVe6vhmEdIDJkgErpdEg0EsWibEw3Z6AIx22De12oAKJEpCcwDg4yME91YJbm5sq++dABb6L4zBGvs9nBTx8fY0TBNQGIogAwMFYR/gu7q+PQQHghzkBbrt5UgYdddgGnTZrjUACjgREK87JOW1BotAuYRFOiRkVaL+3C8etrS4bUAFbDPs61iM9F8CYaqUm/+EHf897S5AGxbghKUX2iwa008DM9rZ2juOSs34mZFIDP2C3df1ys+ZDnfVUECq3L1HwLJqSmr29xR6QdS4NKG0/YskjcmGVzBPlt2m3F96mNkLW1UnO1eu4Hc/AZcAKCGfD7ls0aN/Ey4SfGWNsMBMDilj3Mq6Uc/Es4Gu38lKxeZF9EQ9Gq6yN+bSugZ8xrh6I3OnMYR9ygp0JvzbI6IYfGsUkjC1gsejsecZ7mn8Hw2Cr2zaaT6TzyvvNALf7qgZq44LOcsgEvoI6EIm9aoBflQpw2MEaTLdu5a1D0ccKHHgkPq/HVC2wQsreH9ZXsMAzz2FTNDofExky2sjbZ7anJWXinK48YKqUyv4w5oD7m7pnqu/idTD4N9xe+HwEYtRXinxclyxisFftbwbvbX5oP7TxCpSr7cbjYN94kWUDOJl8ZnJbWA+wjzDRj8oPYJ4CeNEEJQLtBlhBZaDJPRpFp8vCMIYle8DWge+GcyMZAcmE6I/2Q8cK52QMhKBUzCIgGFIBK3aLmidgJBRVJcH9SLQ57JuCngZWWYAe+ySOZyIH5cU0MQMJAbjhjEfAx4mKtWvshPJDFvaK54NG1nR+6rxI77cEUgyk4DGwCVymSvpSLmKsNUmVRb4hTUeVC5XgVMau2vh4Fr14egRmWLHzMAbne280J1PUBgKGBIWUbaQ2kYLFLiGGpipApXXZyEhx2S9LLgrnnPef7eRAhMuNySdyfiqoAXsZNiHuGeINZBEzJjA4jio/F/tiysxR+TFVmeg/BSp2utk8Pe67MwJ5QEW8G9oOFVlp6c0pMN8SO2FgfH0joCI9hnnXsaRky9SKv5U+fmeNyA16ZfSNy4KvRDw93TADK1S50MGRkBGitkPMgEjzPHY+e6xRKRpewqCLrGGlyuW//giACm5yoL+pLicyw5lJAfmfdkulkZnJpUCFZse3pFRWySYvKIQNAhvKBgIMzGpEvQuVK3InmZuhbf6Q8gmBCjdUKVtQGWIGJoL7njkYGQMwtMwoirIRRfTYclEazU1psOA3djqR0hACByUtxoy9sNujNAWAil67Y0AFNDuVNhxKI8ABH5+YYDBpY21NFp8sGlAxKaValUAFgkRuFGJT9w0zZBE4aOCBgLAehxuAIYhBCZFuW1bm52VjdZ1FlJH9OgSjRv1/NfyMUXEfQMX+/czgnzp8TDXIrT6Gyy3hOtQutSwh3BMfU7VLjfZq8xrSTwAqsCmz3nSqmHYEVBw6pEDFoUNSrQ7TyKFhhCA6AhsF9EWlnnBN18VkkMWYKGEACV2D8fA+gIrJSTl79qwcPX5cjWwYEqAwW3HZ2BBSAy1hpNn4JIAKMCqYGarGN+6VMxmiGhUYXst++eTj37LdACrq46MMfCmTJQlU0OWw2hlvoUZFfYRABSVjWP/DsnoCoALaqNeuXJGxkao899wF3hcYudC/p/ELR6MvcuvmTRY7Buvi4L59cujQjGw2GzKk4lrW5wCosAJkYOWk19WdABWhsbtVYGUroILzKQjWaMjTwBNBgeI1uXr1sszPPpaLL5yWvXv3SLPRkz17UMi3Lj0Gt9VAD53b+LkvMGA6XIdUnDnuKUNd9Xa1po0mECWZEr4mu5MVvs/7LL2Oh+MDub6IbWFABcDaGDjJF+xIj3P4PhznRFtRmLDXIWV+mYDmqrQ312RiAgXXm9LuQNYG4G1dpqYOy/rGmty+9bmMjVWlBaDi9AUpFvdJuzskjx99LZ9//rGM1MpSHurJqZPHZHhkRnqFEXn33ddlDkDFf/kHef/t12XvoQNy+sxFKVX3SK+Pa+FeKUjRbTbl7Xf+RZ6/dF5mpo9Jp4fAuWZ0O1CBZ3ez0aQk0+2v7xDchPOztrYiBw8ckAf37nAtW11ZlqPHjsrhw9Pcl3p9ZEFhGe/LZ9d/KyuLj+R7r7wqUhmBuyWrqxty9859WVlZlnYHNZs2ZXFhhWwK7GVgkuzbu5dAxehIXQrlkoxPQLbJgIpCicAOTYkhABXDBPgBZOA5xhwCSwKBewAVyL7H/XCggllaZGL1pVRoyfLCffnqi2uUN3vmmXNyYOqwdIZQMBuOakkaG62o6GUHmXXQSbbsTGV4gFGhjDPsKwj4Y10PpZ+0+LMG20OgArUr4AxOjI9zrWuaTBGCyyhgjTUY4479DY4hik3PPdGC0wcO7IuACjiPCMSjRsTy8ir3UQCES0sLTITQwuS1AfMGY+PrMdriYACeX4BUWO/r9VGVQ+wPcT9ubK4TQNFCpiofhReBilJZShXUkijJZmNd7t35mhJTkH5SEL2SIP96wgMyZluNBlkGGLtQfhHjCKDCQQi0LQFUGBMlDVSo014QZVT0onuCPjvrwoNA6bXF10VPwPCB8z1Js9J13ca+g4QKjsEwmD4qpcFAgyWZoA8EHqwgZxqo0PNq5qKvIw5U0C5gogmKaSuYpECLrllpoEIlMdTM5vwcwvHVbx+o2GU0OgIqwsSlnRvz0ZEJWZbU97EXp/e7LYF8BoTik5iH8s2Aipy+5HlWu8RCtmjTLm/EdkWc0/1gB9xfi7w426stWJT6zm5bpFfY5iQJ1xrBOATRMq6UAqwSZ00dHnnhzlRIN2GXNykTqGDcP3tENFiX1QcN5Ga9EnJAwQEJ2yRMCIQNnHqfy1bShW9L0C1pS3kBecu4H1BgsBtrxZkR1EUyHfwGf9n04tvo3OF48RnVsUgOY+jJx7JMg8cN3FQ9lx2oAdjMGcjjKGNl8rxeN4gBT8vod1CKdgfrZCiLI/R5vG+uoY/3ek/C1aGgAXer3cCgMOFw9R/x8sQEtIf1IIx5733R+hCavMi9huBEzIZgzQIvFG11MuCL43uUr+wL9xqvgQFAhGsqkw0BgqO+mBYz9umpe5OxRcCmadu99ZqT2gB1hb0uBULwBm5hLpBt6TU3raZFLB2Ec6pPqn6FJsKqLdVWNgf2+oyFFpcmQ8XiTjjEa4Qg6I+/UwYJ42VAAc7Nug5W9NkD/kio8XuAnx4o1/ukPiH6qYXBtZB5EqhwcDU5H/3ZxDi4LRaCGW5juO/t8ZtyFbaU3W8DFzGO7r/7XEX/8B0WyzbAJr2u5AEVykAytqfdP9x7Z7Po/I3jE7gXkCB3Vo6zIVxOOgQpwjYQBDdQw//ujGSXtiJbimyJWNGAz5HCD5ZgoABGWKuV7CLYax4OLE2/9k32p/SYPX3/dAT+aEYgF6jIbWEaqNADfcOJvhauqlnG1pYjkH7MUit0esUm8qqgQPwKgYqcFT6jDV6waeCjMK0gEIvyDAEdBF3UdGEJTKU0Dzlqp7sNwa64q5kRjFN4DUOrfZHzU6ZrWqS2k8wr/yEYFZ1iLLnjAWrdbGA0qE4fM+UCoAKbKIgRlBUwoILFp7soQKUFK+G0a4adIfAtK+7daDJQ5s6vO+cOVCDgnmBU+OaA7JchBM0RJBm2QEVcSBKMCg9Y+maMcxOoQCCj2RBIOzHjp+dARdGACmVZAEwBmAFGhbJMkL2hsi7ePg/wA6hodzvMzNxY3ZDR0bGIUbEXjArUPLD+Y+N0mQ1nr7j+uRtBONaDAm4kYaONAR2dlwAqlgBUrKwx8B0CFdH3DKh4cP8Bg3AAKqaPHKdsCY7xsUdfCAw43TUopu3B6xCooAHSAODT0MyHbYCK4yePs/AtCtByvjtQwawJ1R5lxpNJrHgmqEs/hWwSPMdg54RAxZFjx1QfE5lTBFw6UdawP0BpoAI6GVierly9Ip9/qowKSD/BICGwFAAVeL8J0MSWLHwPBuUnH3/MufYy6k2MjkqxXJQh1KhIARVaUL3AgOibb74pY/URefWVV1i4F20OgQp1YArSaDTlxrUrMlqvyHPPPS9FUGEpbaIGO78jBbl580tZWliQ5y8+L/VKRWZmphmg76FysVegszo2aqWb4RrUXHFDLguoyFv6tgzE7Ga9tGLz5hqZw9qTtdVVuXrl97K6el8uvXhRarURkX6ZBbYJVvSQsZKUgQqBteHhqowa88qNbt0OFIxWAFDBabNXE85VtD4H2Uj4W9oRTL8Pu578bJBR8U2BivAaCQc+bCvANumwHsGjew8YvF1enJNnTh+VyYlR6fZB1a5JqTIqBw4eYk2Br7/6QkZGS9JuNQhUlEr7pdMryoP7t+TLL34nM1P7ZOHJAzl/7oyMjB6W/tCovPvuG/Jk9pb87//5Z/Lu22/I/sP75RSkn8pgVAxLv48AKgz2vizOPZaPf/ue/Nmf/4mM1PdKh4wKld0AUIElGYHx9fUNefLkiczOPmHm2HC9Lvcf3JXnn7sgH77/HgvHX7t6RX70oz+V4bpm7COgivsI4PPGlY9kbeUJ5aH6lRGyOuZmF+T+fUheNQhUIEv/3l0wLMCCq8v42Ijs3bOHPwkgFodkdGyMQIRS7YvMEGdziwAq6gwUw88EKKaMii7lCTdbLUr94AU5KdXvNWZPvyetxrLc/PyqrK8uyOFDR+ToiVPS6Q5JH3VlpCz9XpGFvnEtBOexPkZAhTEq8HewI/GCUwVGhQMVvn84UIH2O1CBtdUZfmibAhUtFuN0oALrrdZOqtEpn5ubldk5ABVFFhh3Bh6cd0gxgvKPYtoOVCwuzkeMijRQgfmKoL0HvL2YdlQ/owGgAswMAL+a/MBi2hGjYhCoQNACrIpKGYW3V+XB/TvMnXCgojAUAxXuAPu+297c5BzA2GGcGMSzpAoHKrxtOwMqsBkOyWZTJQu8bgj67AkCvs5yDbJMyPCZ9gQLt1+0zVqUGECFr0MRUEFmXj5QQe10BkGUUTGEgtwGKChIoUEYAhAWPFH7RhkVIVDhdtoAUEEJzRioGCoo2PWtMyp26e2HNQh2y6LYyTYWMi3SYEU+kB93wtvkAbW0f7CdF5J3jT88UJE3Onk3KP/G5fUB/qMHLDm2Qbb8bscpv7XZs4JtGnB5PUA+2JdcOyCj298YqBjwWa1XCNha4Jt5QCz4nK7HGI+Agm6DI5LHGoo96MHv5MkpZZ5/KzBCjbHcRy6WTrZaAiS6BJKc5r+jD8oO1DoMKn+jcyejvLIWn3ckInV5XTu2AiscxIi/uCXGZB9GR1tR8KxOMxBt4AMYlWo/wO/QjHpltzsbIby+R0ZNCtqzwD1Rx5hsHA+Tz1LWg9rD7jvTvzA5KLBaKXPYapG9Dz8RdhQBoCEHOpQxoQwJJPR5JjyUFTRojcQ2zBdm41uYF9fzxDzYMB4noF/JLINAestiOJ7tDpsF44GkRRavpm2k54ZENZQTwKRAXxnMLiiQ4/4AZRhLRdbqRLORcKjjrj4CbB90hjUYWkgyVMCBezGTBbKTi+KC5ip3h9iJF2GG78ri6iyKjqQXsDvRLg2IU/ZoCDEDn5cxG1/XGL3vrNdRQDIBEnR0rOEfKlM8HvsUdWBgqulcQlKb1WOw/gNYwphx/8E8sQQR1j7bbFiAHzEeMCRVliuZNhY/NyHbKds/Su5W0ZqS+LM+wyqllQTcOHfNF+ScCSSiQ5823Gc8RoIxDRmusI8RS9EC3srkc0lBJppZzJH+rxfthocDf9tBFXVE1Fd4ClTsxIx6esx3cQS+GVDhm1X8dGswyUcgz3Td6QjtFqhIYRTpy0RBNDc5c7I8tqRTexZumCXgGnt2wSCDQK8QZnqkgJPobQhW7HR89Dh3jCLzN0YV4hMFbIs/JqAiq0aFGgoI1A8CFWBURNJPlPhQ/UxogJfLKh0FaRW8PNiMa8DQgFQSCp96JiOD+ciqsMJE1PJ2NoxlRqizAikdFEJS8MOzMRFkYH0D05tUWSG9Nn4iAxZZHM3WJjNR+zCkkC07VGZGJjaWnkk/AahAEdGQUdHvaYakAxXusAOoWFldYb2GbqtDKShk4lL6aeqgaXOCOhrTQD2whHO5VrYHJxyU8P54QNh1R3WDBILflqUnC7KxsmqMigrrK9CUMXkmjKVLP+03RsX04WOUgHKgwvuB6zLLpFyKMktDwAdOYyj9tAnpJwuUeTFt1/jtd3qyMLcgV69clemZQ3Li9AkCFagzABoFgUcU1KZMhLIp8C8CKswYbzc31fg1FobT/9HOd996m9JP586dkyNHj8kQJD6o4y1kHQBoCtkvPg/cmIiLaV+VT69fl5/+9KeUqYJBhheMUBq85iBEQAX9KS2y5tJPCIjWx8c0+8ek0byOBQ1+Lk8qmfbGG2/I6HBdvv/aawSM8HcEh/AZHQUu2EMEKlBMe3S4LM8/fzECKmDouksHYxmFhRF8unTpBakho3m0LoePHJJOC5RVNcoVLDRWBQLzFAjT9TwEHBzMSQcOwgBMbMjvXqoibyXtoxC7bxfGLsH6ubqyIleufiArK/Py0ssvUQ4GUOnY6D4pFYchYEKwJrqnQT2KarUsY9CoR1a2OQvRTkigIqhRwW0k3is96JCVieNOgJ8rPVbh+0TwohAUddul9NNWYMhW1+9Km48k6skszM3JVzc/kwP7xmRyzyiD9cWhCguV79s/Iytry/LVl5/J2FhF2p2GnDz5rJTK+5ndf+/eTbl18/dy6sQxufnFFbl48byMjR8TGRojUDH7SIGK995+Uw4c2S8nz16UMupb9AEo6XOOAvc3P7ssjx7fkT/78z+TYqEu3d4wHYw+1gDcy56CkCsra6wloYX3+nQc1tZXCCTcv/u1nDx5Up7MPpYf/OD7Uiq5ZrA6tWDm/P7j96TVXJGXXnpZCtVRgb/54MFjeTK3oEW020158mRWHj6YZRB2j0k+QfppfGyU2s39YoEACdqEPQbzDoFXZqyXynSOEUAno4IArDIq8HfoPiOIjHsDMAAONdhWcCKbGyvy4N4teTJ7X/btRfHsMzJUHiFQI1a8GKALpIPwjJbL+F5HKtVh03/WfRhABfYxzA3f7NdV/wAAIABJREFUT9LFtLUWhBathuPlNSzIqOiBoTTJa2xuAqgAjb5KRgXWYfQVxztQ8Xj2IccBQIVnWMIpzAIqFhbnWagTAX4CFYHpCCcUAIrvO2ijSgOpFjAYFfi9VqtHQAXau7m5IZWqZkDiOIw993VINkFyj5JKIo2NdXn08J6UhgoyOjZC6ad+Qfde3UZUV9z3XewxWUAFxgtABc7vkhJgXrj0E9qhSRlaswLndOAfD12zqQkTlA/gnF6hreN7HO2qQDIjtFV8HY6dYQcqdA1xJxvnVNtGgQquYZYBG8k5Ym8BwIFgU7stS0uLUgqYD5r9qoEZD+Aw6MGkge2lnxTQsCLeCaBCGRjfKlCxS5Ai0x6P3Y3dGfZbHJ2XKb4VUBGGx50Y6MenPbWtur1boCJ3D869SPYHWwZkMwPO3wyoiMZkG6ACY7Z1EfGcnqeC/x5Y0kB/4LKZd0f/LivHLpQPSl8q1fUtPfFUYkTiVNsAFTq1zR6C9bpF4excRkXOjc0HvuJRT3QzHDvXvbegZ+adyAUqLMUwir8b89WsYM4PA2cimRiug8aGZsY6WAex3FBkB+oCEduP9oGdMuDzpMGKLPAisgizu5dxL9SVyAl2O3PC9glm4FMKN062oY+CwLvVB1JwzQpCR0HTQGqKUnsBeziQsdGvar8QDPb9iD64sdUBVHimPPwf+IqUZUK73J+ICkjrPaBcEIt4q3QlwQ8eo6/IV8UeZUls3gcPEuM7ZBJYIWvW26pUI/kngABkP8CEQk0JSCUVwP6AsoMqNjARjkWntYYX9mjWISmXtY2QVYxqm9g4mOwnr981NovLb2m0PBtaM4YIC3vz2vBt/acWxVY/Ip57XicFbVCARBNkPF5FEMOYHQSWPNEqkn3qq+ykSVv52MaLlc/Z5GJEaWCrTaXMnLimn9reKq2EewEwAi/IXqHxnL82/5Q5ofJUunZaXQlIP4G97n0NQNJ470qtLrYhMpHD5xXPa9KS9BV0XiuDB/dS56zPW691GfqufNxt0AHqoO3OBHFmjcdkIkaP1b5RdER9f/rS/F3nuN6bgFFhQMVTRsW3ZmI9PdEf4wj803//sS7iqYzRRFv54PtjrOi7fSlACMIFILUY7NboZ+qBtir5Slw4/sgjgYmDTSM9Dkv9O4bfw3XapGjrMwmPLGtSM6K94xbENucu/nPcHz9iN40MDcBkrg6uG4xdAIrknz/bPPxDMCq60H20GhXuqLoUQrfX0TuGIA21AU36Cbr9xZ7WdwiACgRWEJfnRtuLGRXoJzY0XIdZDP0ig0Gh/JPTR1UrUQEjgg4+vVl3V4GKyJgaGmJAAIEArSke13TwDZuyC6UhynIAhHCpWQAVDEQgkIwMLmScbjSoS9gFxRO1EkBr7bT4MwwaYnMDULEKDW1k17Z7MjY2zmLa5VpNDkxPM+OA42bGJA3BTpeZzi4F5UEb30g9mOHBFHyfxawQMCNzANkjbVmeX5SN5VWpDw8zcwRFvSEx5KkN2EAfPkA29V3WqBgdG5WDM0eZKYxreCaLZ/uClkq9bwR3nTJrk82BCgTuMQYAKZom/YSMaGQ3qZZvgUHyR/cfyReffyFTMzNy6plTlH5iQWSTmWA2OQIcgJ2MNuyFzVkDJSim7ffQwScAFe+8+RaBivPnz8uRo6hfQB0p1pHAvUPtFYxvOgDkgWYWt+73CabcuHZNfvaznxGoUKPfWQ6auYRXEwCBGSrM0Gl3CFTgWq++9prUR0dIL2fghxqpBcqIwdRiEW6AM70egQoENr//6qvM3MbfHajQumtYy4sMdl67cllGhiusPwFZLwSFmh3N9KCD0OvLzZuoUbEgL7xwUeqQ/xoqyP4D+2RibILyI9pfhwH856DOch5IkQYmwve7WRe3OraPNcT3FmsaZ1JfZGl5Tn77ya9kfX1ZXnrpIu95r1OUyYn90itUOJ8UZAgBaH3+x8brDIJmvVxvNEqSCfYkNYKzDXucKw1k+PnDoFEygESXzUIpSiHR0ysolh/QiunzOxnrxPV1lSCrcahX4Fr28P5t6XYbMlIH7Rz1ZYpSH52UvfumZWV1Wb787LpMjNf42clTz0q5fEC6vaLcvfuF3LlzXZ49e0Y++e17cvHiOZmYPCGF4oS88+5bMvvgpvxvP/+ZfPDeW3LgyD45eeZ51qhwoALOYrfVlPff/RcZHavJK6++Kt0OZJ80wN8vtKQroFaDSdSgjND169dlYmKP1k/odQkgPHhwX44enmHNhONHj8jx48dYC0kDMuokQYj4N796S4akKS+8cEmkOiqrq0159HCWAAgkn9bWV+Xrr79ijQq8UKthcmKcxbMh+1SB8wqQoAopJg1se/0GXAn1EKrDw2xrq9WxGhUqwYA1DmsPAum4HwAD0AdIADY31uTBnS/k4YOvyWo5iYLl9QnpSk16BTjUmFvUlpLWphZOhoQizjs8PKpavGbBoB4Ozou5GBbTDqWfAAKglhHar+cY5t6NtiWBiiadaQAVXpQagQCALtivwah49Pgh90lIP8VSfCgqPsqMSWdUgF0yv/CEAInWmlCAJXw5iIPPQ6ACbdtYb/A6ACqY3NAHaLtBJiTARw9soA8KqFS4Z6n2c59AxeNHD6RSGiJoSyCrayw+YyYgAK+MiiLnA2qfQLKLAQx7HtFvjKszLdAHBypcwknHX4EKtMX/jjWl1dLgigMVAGf8OE/aCIGKMPMvdLgx36IaFbDDjAmBsQJQ4ddFjQpGauzlQAXmoGo+FwhULC8vSZHyUZo8okEPzyJVSSm3n3ifRWtsYWzwT5+FIc6n1ZUlvlegIq5RQftlqMJ785ff/7tvr0bFbn0WjoVmoUYv//UbnCsbkEidMJAA2jIg7Q1yUuAW7dlqf9jJvpA4JicQvTXwkLmD5uyrvkLt/Dt5QDymc1SjwnxhjWfrYKXHN/AIdz4sGgcfeGnQN+MaVt8r/QU/ficXVjNyyxu+k9NEx2iAPq47pvaQB6gzTpU3B7LDrgNMluQZs+0k7snulwePSG6/c4EKI9kawyCSJeJzFiQqEgzxOglgiJtEKtgVKE7MQGLOE+kgQjQu1qfE1IjvVxhkzpg5mfcuWTsiCB9vMQ+cJYPnw1mROlnTk1b7lR7bBHARABiepIPAsso+JQO4lL2xGnDOusD50QaXXMTv7rdom+J2aWhK2wj/BgkNzgSB/4j7Af/JgXiXfFIZZ53LUUAZx4NBYHtY2EfsVW6LAKjwzHj6Arbvue/tz2cE9FiigderQsyCNSoD27/bUbYH60WwaDV+h+STsu5VRnzwBfYFAvw4FjaGfl8Z8Z5k4Lac7sPK5NBkEbVBIrkvmoNxQWwyRgCE0G/UDH8Wl0dygfnWWhQ+Lk7u1wzQgiDcZUCU9Zv+Mtk02je0H23hvbGEUQcJGH/s6zEe8I9YH1oES9UJ7NnWqa7ramLkEkovCt5FTDoyhwwAIciFsbD7RPbU/8/ee7/JcWVXgjd9ZvkqeBQ8AZIgCRAEaJrNHvmWWhpN97Q0q111z/66s9Jf0vpT9tv5YY1mtJrupvdwhAcdCO9dmaz0mfudc++NeBGVUShQ1GioD9miAFRlRka8ePHevffcc442e/JyUZsw6XD8DPM4jKsSd8qaVrBO+HiqikIs+eyrgG4FcQzrDFR/DhWXMT8WgB8G9MXAlzzxqHisHe3Jm78XIxABFVkdFIlNKaV3miiAZ4AIK8WSWSPkMk7ptTmqmgdm1owiXeMxDZBkn1MWNXt4gmAn4hImHrYmJKiMJmrXlD6OFjGDzuBI24UXwE+ptdDqX1GHRMSasCAiQIbtwHbQldKZ/75ABTo2sEE5HS5KqAcAKvRc/ilABTYNJP9kVBhQATmisEAQFZdB3bUOC/pS+Hii6zyviXf48sI7NBSxYbGon2BUVBkgNdtN6bTa7JDAxh4CFbj9CJoAVKAbA8U9ZVCA9oru1Rio8AAIRf/FpbrUFxbIqBgbn5DJqWkp1WqyDiwC6+ggUEGKpW6y2PxxbNBdHRgKgzO/NgctvLOToEIOQEVX5u7dk/qcMipCoMJptdiBr1+7JlcuX6G+O5gU6zdvpVnsMKCCEiNWjOASEdFg0aesNFZ+P4CK+pKZaYMcgYKoPfKAHro9uXX9lpw/d042bNoskH7asmWLVKrogjfjTho943jqUeHsDe9s4BgBCPOnBAwaGlQp82MZUAGzMY6xPs8IqDHPwuvwY3G86U/Ql9OnT8u50wpUgPWRw3G0YhidE95Pbwg7NpYcBKMJoAJyWpBnSgAV6NSBBE9fz60/kDffejMBVLicE4O/KBbKE6iAmfbYCBgVkH6CvEmRQAUTJdMr/frCN/Lw/j3Z/+J+GaVx7UBK5aJs37pdJUiaKEiHHhW++CcX8nTnSThW4e/CObH6VXGFd0IiEIwKRnugQ2shX4GKnHS6fVlqLtCEuZBvy8ED+2VsZIJSP7XRGRnktQM8DQwgKR0dU2k4N26Nz0IDbCYbiOkZlDuIE4MDmpAuT0b850MTw+BS4987UGHH+mcCKhKjDPo9A2yAy+Tiy8LDO9LtLkm325Bef4mAGBgV0zMb6FHx+blTMjlRke6gLbufep5ARaebk8uXv5Rr187L/ueflU8/fkeefXaHTM88JYXyjHzw/nty6/pX8lc/+3P58P13ZP32Gdm5+wUpQPopNyKDPrrdc9Jaqsuv//E/y74Xn5NdT+2RXmdEBEAFh70lHSQfkhd0z9+7e1+++PIrWbduvbRbbXZywcT5/Plz8urLB+WTTz6RP/z931ez5KJq1cJ4mt1cvY4c/vgdqZb78uL+/dItjsidO/Ny+9YdaTQgkdSQW7evy6VLF1nABlg4NjYqa9dMc42sVct8httkMQCoUIAQmvuQCsCrUC5LbWSU5wo2wtjoGOcT1iUwEeBd4Qn99NSUwN8G+8DNa5fk0lenpFzOy549T8n4xIx0pSpSHJMOsPcCurMwIHlptwBI9g2o6MhIdZxggq9nSMQg2cS1yaSfhjEqsKdD+xj7qgMVOG98bmpq0hgVLSbVIaMCsk/KqGgTGLpx87pUq5VlQEXMqIBHRUFqtaqAUbEaoALPLcYpZFRAzgpSUs6oAMjqjIoK7o2twQA4nMWAPUv31oEsLS3K7VvXpVIqysgovJiwnsReMPhOFGh8nwPD0hkVHjNgX8Z14780UIF92xkULuMIBg7WZ1wHuhoRQ4FRgTEOgQpnVPh6qutPbEKatbZ6k8MAcVgAVLiEFr43DVQ480T3Ci1a9GjyngQqXE/cz8nPRwEIgIdqpq2+JepRkQAqAEpg3xsCVGA8v2ugYth6zDg9M1cK1u8wZHxsoCKLN5FY8PX5DGKWoTuf7yl2Pp5pBPT3xMeyrvlb7b/fJ6CCkrIGGHjDjG7cvPTvBKjIGEQtdi7/JRtyHuM17N6FZtrDMrzMqbkSwGDPuRfRVgQqVgAkhl2adg1nPzDRkxGAdGjSiTrn4866rG92NGLoyEYyVsau9vg3AmcsT9TmE+3k1jVB9z0UdbUvafi9cy+G9P3mFWvd1l4OyiwHBay+Oxz1wk7uMkHpdSrjnqLYqeeNRoUOmwHAANCiswIDuhZrIZkF2ijfjcEd79SPL0GL0FFHOoreaPIi41tBHZf6wb81fihEXgju88GGtfDcbWx9viNuchkiLSDrsekzYIV0Z61XK5Bu6src3DxzU7wUxNd4h2xAXp8y3QECsDDOznploiNfUNaJ+x2KmW6rKTXmYq+rY6aAAOoEuQgwgQ+Yd8fjPLHf4bucocG4L6egA9mfWT4v5hnGJo9Wm9JMPgdxDwhaFLTBAteAceHeZXM7UmzAfXD4x1gTbM40xj6aEjjXI3DCPDnMG8FjCZcH41gaAyE5n+MVyGsNblTudSCj4TC+RYMMpdVsTDUeFcYIaPDB9ZKBY2wfZZ0Y+8K+mP9iymXfnZKNTxT4TaaX7GrktnaP8R0AeBBnapyih9PxU8Yx4uNkA0i8vNArDpLXaJIEA8fAIpyYmpWr7wb+I+vG2RdUgdA6jm1NtkCowgfVFkzOM1xvck88Kh5j13zy1u/FCAwDKlYKxHUT8k04DH1Sf48j6CQmH3YBBRtpIq4fuqFqUj30xV0/FdxEck/BkflX//fwYChDRdRqS3HxJwonHMPw4pOvh0PJwVnjpRqCUdHXDx6eauIyDJBYoUNi+DjFBbLVTs5ofY8+4AE9GAG6UCJwwcaChRyyNQAIlppL1LVGIQXFdRQA0P251FiSfgmSH1owpnG2GXlxZsFI2imnrpPZ7WghuDBgJ/lqGBVYyL2o4tJPkL9xaQXMcSb/kAEqFiKPitDskcSegiUqQfLixUoUmvE9KEB5hwUCHbAO0MHfgvQHCjzY2aA5aaaPLEK79BO68dttelRohyGAimYCqPBj43sWG0tSn18gkwDABYCKcm1E1m/exA3TOyS94ODFAHYbGFiRZmp4F4QHLgjgVA4KJmTYD3vy8M49WZybN4+KMhkVqHORcojN1IAKZ1Q4UAFvBO9G1Q1fO0TwP3anshgUJ//a+RKbaeNccf8gd0UqJOeAdtFQ67LTk9s3bsuZM2fIUti+cweBipBRgYtgl0leA1IPRBkYmvwXurCjx85YKSzMdToJoGIrPCowziyWaNEaeqi4194hqomLPqMM8AJGxdnTpyOgAsdhcGXPEJkQBlSwg8YSWAS7MNPGn2lGBZ49ZVQAqNDOGwIovYG89fZbUqvWIkYFgAp2JjlQwYwnx2f09MkTMjZSIaMChTCAUWAE6TFVvujChQv0qID00ygkQIxnNz05JevXbWQ3LORp9OWGEFl08+Vpc5x4xOtb2PG72jUr630MWk36iekGwQrMXV0X+70yYEKZn78pn3zyG6lW8/LSiwfoFzDIj0i5Os4iMj8b7V0KksO/AM+nP3fJc9CETbthfA+K54cG4N8eqEgDJxGjwq5Lt4nvllERznECWQNNdgBU5AjAzsug35KlpYfSas1zTtZGJmRqegP3gHOnT8jEJOjmPdm9+3kpFGek1yvIpUufy9Ur5+XggX3yyUdvya5ds7J23S4pVdbJhx98KDeufyl/9bN/Kx+8/7as37pGdu5+noyKgYzScwHP4P27t+STj/5B/uCPfl8mJ9dKrwsD6hpvySDXkjb2rYGwcH358lVZWFikJB/unRbRC7KwMC8b1q0h+PrGD19nUTwyyzVGBfyRjnwMw/q87Nu/T1r9ily7fkdu377H4j+6869eu0yDaOAbkxOTMjoyIhs3rpcN69dLuaTJRqPTJlABpgbWXDAqIIuEtaFUrkjZpJ/gS0Ez7b4mSWBbYCyxt2INHh8f434D6aIvz50U6czLnt27ZGbNGunnStLLVaWXq0m3j650lwMAoA+gAsdDkt6WkYpKSPm8xJoN6SfMed9TUbDGOWCfQGEDhtbwMvJ9N5R+wnHA9iA7rglGxXKgAoV1xA23bt2SGzevsei+fv06TfZZNMmTTYLvnZ9bVN+oalXgUQFZSJVwwj2K4zqcL0AGnOcwoAJNAio7pUxLADdupg2gxM2000CFLnx9AhV3b98kMFQbUaDCO/K8ucD9KXAdDlR4I4Am2b2ooQJj4B4V9+/fT0g9IVbBf/i9mm5XVG+6B98PjaV8DMGoCGMSv49Mak0n2YsL4XPMVcLYmIjDHKjAHoPCDhkVVTDpIF8Zx+IeP0Trd15lOSETGDIqWMiwOFnx+bgrWRkVw4EKXPfiwkMWyjjGBTARUQjyfR2eIWX5vVd/8i0ZFRkl3G8BMPxT9yj9/CqAivQXPUYuMOxqvUL62Je80gU/xjnpHF1h517hd8s/NXwvXfneZHzBkJNCXkA29Xdzs7VxInyxsIa9aoWCfWqdi+KH1EeG3uvgu/xzmhon465hlwf/vKE/zxiNod/vcrEp9ptNff7hEjGu9KD+D8p7j54Qi5m8sSx9XpHXRFiw93EbEm+FxfAo9V5JHiv1heFTiyZv5A5YG903QWP1IS96YKSngN5I98DwvcKfE2Wx+R5tn42KswqUeJHTi79ZsymLZYQZ7hJGXJP6aqRMXwMr6uObCYzQ9Fo78LWZw9h1oixRvAdNIBPj44y38ML6TWDAPAMxF1EXAMMSL5cH8mulx0FOC/BaMFZ2Hgq/KBSjcI2cTn+vuTC9LW2fxffRS4T1ig6L3bxHxuDAeaNpC8dBPEgejRWjfYw07jdwKhr2pH+J+3c16IGlTEL3dyAoMlAgBLEB/MvUW0v9ICgXBaCoa2zDfJ7n6Cx3VZgAo0PHDmwRekKZ35M3YrLQTzNuk1Dyors1T0RejcaMxHmC2asPVwwuYTx93ijDwjwqGCu3dJxwX+g9qcwiZYLE+YYCMPC5gHzu8rnqU99BMQdTuA5EYEnS8NrnR8XYJPqsoMFPYwI3/EaNAeOFfyNGQPzpjRGou3BCYZ5b3KPskhCYABtWx9GvqWP3BrGYzi9VRsjyEeF1BJJ0ZL4QiCmp/wr8S8D8MRYzGz2wVpiShzZWaq3BQT8CeuZpgbmFGJgSaZhvT4CKYavsk599n0fgV//bHyVPP5Q2WrYRa4gQU+/CN2QV4dPkwZiOFeMGjwqndMnSZcv/Hn+3dnGld3s7ZgCYrOY+ZZ4Jf2ERZHCgZIxpn47emw4N/Oh6LfErda7pSwwPE37scSNlY3WsZhwSdzYyW9JgltdMffdvB1R0KxXpYmFFgGNSAAgacGl9dhGR18BiQKfVkl63xSQ/h0QVplq2aGPz0A2oJKUKkGgt2mKx5ubYQbGoIYsLkG4oUaffgQqXOkIH6lKzoQFPsaidJZSoVNooaaAuicDsIZ7POFfMPWxYKAy4vJEXLLEpIshgMGEMBxpREynXYhOKxOiYjxgUKGj2FJjxjh2Xq0JAg0IKCif4/ejouExOTLHItXbdeqmNjRIA8Y04vIfOIsCfKGR48YbXZl0kXrR3vW98H7w2cNH3796TuQcPFagolXjN6N7vQW+TBW+Ra1evy7XLV2X9+vWU6dgwu5nyOQioMO7eRUEGQ1+7B5xJE3VloPhvxnIMnsyQFffR2ll4A1hEwTzoojB5X44ePSKbZ7fI9h1PyezsZpqzOrNEx9t8JfpKe0UihACXHa2dluQHBmDYoCHwwvch6AWjAuAN2AabZ2dpfsuOHQNdIO+FwBISWz6uHmRw/iCg7oucP3tOTp04If/u36r0k1SKGoiZKZkHHjQLM0aHPmd9OX7kKAGtV157lbJakEDjfXOJFqOhdvFdCL76ACrelrHqiLzyyiuRqTnGHQGN0uUBkuTYhX3q5GcEKiDr5B4lEYhjxuHffPONPLh7Xw7s36+FW+tgQaFudnZW0K1Uh14+qO+21sTU1UevOiFAHiXQQbDmAV8aSE//OwQ8Esdkodr2H+9iNMBLxz7H+Qwg/v6DG/LBh2/K1HRFDr28XxAD18pTUi5OSrEwDqoVjZmF3gx9KZTKlPVxf5joaoOuyOHST6ADxx4WYflDZbT05UFq1igmk83khpFORMMx8WKhHze7SWF5Mp04FwA+HhvAALFVF+kB9Hkg7daiSL5HE/ipqc3SaHTl5PFPZWJaE7hdu/ZJIQ/mSk4uXDwn165/JYcOHJJjRw7L+vVVmd0yK9XyrHzw7gm5evWk/K+/+Im89eabsnXbFtnx1F4ZlCdlkBuVQb8kxVxBzp46IVdvHJU//pOfSH8wJv0+QIqKRRA9aRhjCUbaRw4fEXjq3H9w34qcBcrc4GfXr1yR3bufkp3bd1ghW2UJ+0YPH0hb3n37H2TtTE3273tJFhYLcunyVa7PWPsh83Pjxg2ut2AoQYYNPhKzmzbJpg0bIy3eJsB5dmZhjdTOxUqlpgaWLA7XeAzsi0jiCVRg3ysXpQmGXQN76UAmxkek32vImTNHZGnxgWyZ3SRbt+2SQQ5rNTrhK/RQgIwbV3XryAK4oYmaFhngz+IeUg4uw8+BHXvtDhsQsMepJ0WZrKqFeQUq8HdnB1B2cWmJ02RqaprrGNZx1DEIcBCohowRWA3KqLh167Zcv36dRXfcAwIVRpEHIxLA6/y8+k7gM3P377HDDsAq1h8PD/V5VjDB5QRwX3VPQ5ciOvNaBGWrFcgZlkV6eTZYNJtgXqhHBcYIQDnOo1KC9JPFCNKXxYV5Aiu1GlgvACp0TQ6fpRCo6LS7NG4niIAmAIsBKafVavDcnKkC6SfcCzInivAI0b0lYoAUVTZRGRUaK+C4eB/mn3sS+TVo12ifTDuVxAgKE5ZI+57FpNpCVPzR63T5TCCuQvcmTSQDaRNfv7j3mXk2xpyMCisAKHCDogfmmUlAmFeSAg56TMwXBWKUUeHFpvm5ewTvwKhwEIg+VrwWgFQV+d2Df/wtgYohq+rjxta6Sj96k1vVO7KBiqza9eNAG8OLpXru39UV2Ka1qquN97istw8/K829hv3unxGoCOJ/fvNqUtfoLIecq4sBDJuCQyWNk00Nvl87GyR9mEee3hD5MB4rgzX0uEBF5h19BAAQxn/aGLKcWaDXnO28GIHWy3Jmmx+cQC5f653YOqfCcc0a2/S1hc+g76Va41DPuDjrH35XmE0GU8TzAb92vVw0nEEeB6bRgWdH8DkdO5fn8oKxFjuHvbKAChwHa6x3jus16c90bPU6PLfUYqv5RNBDQKWH49+rbA6autCwoV3ocVGWBs0mB+g5KY4RNbfZvUZc4X4Q2hymxWbEJogplAHa4j6Pn+G8uIdChnmADnaTPEKzh50nZanMawQ5G5kZxrRQwEflvkI2tN5a/bmzH3EmaMgsQ9oSPpZo9uoL93ssVaxRUGJJJQwJrHQBluRZvGb8YESusHhOqeSiNcjZ8+CxuxfBcZ5kAfTQNKpseIxpPI8sD7amRXwe8Q89KJjj9Xg+bJizpVWPbf+EDLHlm5AXhV8IXh5f4X3e3OGxJcYDc1VBDKizsB63AAAgAElEQVQl+GIY7DeRHJgCBs6E8cI/QRk7j+iabSLj5/gZ5gNqLXj5PAKQpSBXn/MQMQVAFB8TKmpg/lnDBGMV1gq05oG6DVYXfr+3W5NdojUPKhSY5BOfuYzFjjGUyUZx/KwRkl4cmKfwPbMx79CI3ZhABl55MyiHzv1GCAhqc6KykPRZpMzZE6Aia9t58vPv6wj86j+lgIpVRV7pgn1WOKQbSJJSEY+UBkTxv7PkmOLuXH9v+vseAVQkmBv62axlJVMSKgIfuD1FJx3FChqRhL9R8MRfYVSbETBEK50dXv/QhDtxdP/6dBvGoyZhRvC58sdsQ7FLCZHhbw1UVCtc4NmJQVAAXSfmVQCpJSlIQbRI0EbxtwsJpwZNkUOgggaT0NSEKTM2zr4aMWGzxX/9bpeJrwMVSOSR+OO42NDxd2wczU7bCijK7ggLDh6wUrvZYTJjE6JAyaDGQA4cH5vhxMQEE2/vHnWJKbwP35kAKpaWIlCCAR3mpjFIGEiYGSc+i2Oj0IOiFTa4sbEJmZqcZiAAdsXo1ISMjkMaJNaBjoJ1C6q0QxUdz0s8VojaYx7guG6ujT9RREJxAN2Ri/MLLCBVi1pIoHwVCrGs3g3k6hV4VFyV9evWy+jYuGyc3SSTACqi69ZuB++cYdHHAkXOb9vA9bnRoIVAQlvvj64XysZQPgXGqicPHzyUw59+Kps2z8rOXXtYNKdEBYMe9+wg2kRwzLsVVBOzx2BS+uoPgu8kQIQiCXxOAFS89TY7gV7Yt082bd5MySYe24zKaIbeB/sCBUPthInWGM0yqI1z7sxZOXPiJBkV8NEYAKiwJMZBKc75tntU6FFCoOLlVx2o0LH0wM31Mjk2+Hm3J2+/8w7NtF8+9LICFRaUEYDoqqRZCFSMjwKo2B/NfwcqaBo+6MtFSD/dvS8HXzxAw3h4lGiI2ycgtXnTJnqJkCFk9H0WoFa1pyQlNUKwwQM0nyPp9WoYUOHzOnwvZ1WUl5rcguutGk+QMwud452GXL9xUY4cfU82za6RF/c/J712TqrlGRmprhPp47owMl0+AzA9Bpi1zKcCYKYlOLH0U5wwUq82YFSEz+u3ByqSI7QSUBF+XzjOw/aElbYbslMMYIQk0uLinOQGPVlYmJNBryko6tfGx2Rmeqs0lnpy+uRhGZ+EB0NRduzcL4X8OJ+bry+ckdt3rsihQ6/K0U8/lfHRrmzbCaBii3z03jm5dvWE/PKXfyxv//a3ZE/t2PWs9EvwXqjRT6QoRTn80fuSK92R19/4HWm2IamkbAswZ9DT1YI0FQr89bocPXpUdu3aJXfu3OGeUK6U5M6dW/LM00/L0cOH5cc//rFMTUzqusV7BRjVu8y68tabfy8b14/Jvuf3y+27Pbl69TqLxdh3AFKgWIu1C4mdF9+3zc7KmjVruS6AjbXUa3NFU3BVgQp0zGM8CoUSPSrQeYdcGkV1PFs0ZyyX+HP4w4DJAimts2ePyd3bV2TjpnWy55m9ki/UpNWBhB/kByqUw1MDSC96YH3Vzk9fT0ZHYAquxW+8sNYDnMC+1W7pnqpABfwwADgUZZ7gtxYQsB6GHhU4NjxAoMNMwNmO6c0C2GPw3IRABY4PoIIFdSRlgz7XMBSk0ZGJY6Ko//DuXe5ZuHf4znjvw7IDeaY6zxPfBfmiBFDBJFHNtGnc2csZUAFzbmMnovAA6SeARwBl0MxQ0MIZPBju3r0jtZGqwC8jBClwjYxF6E+h/4FlA+knXIcX4XW9b0ujCaCiog0AvR49KjD+vhfjGvFvAEPVijJAisWysVRU0hFjhvHFvFZPIgcHdA+htrFpTnMvTHVlR2wwdnPrQon30yNibp7X7vtqCFT4vGExgjIi+hnMfT+m/okmBDW8x8F9r2RjBbpxc0KZzhCowOewPy/MP+A883gh3NvB7sR9/d2XfsznhuAZGFJsWEERwCQgwzzgUbHwt6rYf6sPDVlqHx+oyIIYhp3Rvy6gYuhOlQm5pPc7/zSLQcGh0mM0VKrnUflW8HtGrUMOwhg2o9ju8Ur6axKF8ygXHH4yqwUqvKD+yBggS9Io8+caw1pAnDjJrFnOfYc5FYqM2tXubGMeIKL56xFymd+t35sYIo/NzVcjkn4JDYftfNWjQkENZd0uf8VSVPHv9DOxWoADDSxAGttg+ZE0lk7OT91nWGjt9c3PTwuoyHcjiSc732g5D0Egyz9Q0EzvT9HcH8ZsCQAIHf/Y+FjXe83RWJ8wnXwvCmPtV7keLbr7HQBQABYkCvJ4T4WSRKrbz1gHBdscgAw1S4477LWJwueQ+gFo1ztztpwyOTx3xfm5BwN+pgw83W+omEAZJhS1FSzQOa/z1Pc9nA8ll9xAnPK9vpq62Y+eEuUujbnAInjgbYDJh7iHBXjLfTk3cmiYA0NSGzS0mA+gQMEesjACySswCHVeuckz4jhtOqPPI03cPZdQYITs4DIYD2i4s2YUa9BD/Ih7gzFXTw+93nCO8L6gcTIC0AxwQy2iUiaLn2M2gDpCkd9PcMSa7DBncd9cSgyNNrGqW1xX4v4Mv0ljhUTPhvuF2r33+e3gEBUVrImFHihowINSA+bFQPN8vx5cB6/VvDbYiMgmzfi5czAKdS3e12LRwAplv7Ap0DwlHZDxGg3nS+ZzpGoWiBEVQAoBLmXHaKOSjaHFRnp+YA4pQMbrJdMCNSqto7B+YPcAjxuajp4AFUOX6ic//D6PwK/+048f7/SjHSO1caf8GsJtmwWMIft8VIxKohXLC1t27BgGGAJULLuKEJDwkr8mSApTDE8qVgYq/HsDoCJM9hIXmZY8CT4bfTzFHw4C2fA8NIhOoBe2aT8yDE2OyqOSs4xQLN7IkxS27wKowBXAD8BNimCYDaCCWucokAZABcxsUbhxRgUWbQ1IisaoUGooNip2qmcAFTgui1IwtubOrxsAkmR0e3jRBn96YjwMqKABn90zLSoVmDBPTU0xYaY5q52jF6JRTNHCqnY4oujjxuIeifXNXNNReC9+YowcqEAxbHx8UqanZriZjYyOiZTzMjU9zSKFvxSB1wDEz1Hv58AMWrUg5Xqb/h4HbJAsgFWxuLAgjboWqBJABYxErOs/ZlRsUKBi80aZnJri9Q5jVHihys8nGnfWcZNABTtzcS18hLXIzHHs9QlUfPrJJ7Jh42Z5avfTlH5CIZ3dVmZqyuDGOoKGARVgsVBj1cbJu0oQ0L775lvKqABQMbuZsldpoEIDFR3rqKMlMrbWMTp98rScPXFSfvrTnypQUVaPCnbuBEEVAkwPPigz0O/LMWdUDAEqMFoIohTIMdZTry/vvfeejFRrcuilQzIyOqIMIbvXHowlgYoqZZ28iLYSUIEO4gECaQMqECjOwsS8WJIWvCos+dDulOGvNMCw0vvSBYZHfdaBikThPwAq8F2uGIghY9cRQQUNDnHtnU5TLl78Ss6cOyE7d6yTZ555SnoddG7PSKWI4rcehGOQLwhkzlggDNZZ/tbATIy5Jl8xUAE5IT9Hf1Z9HMK4N/27lQCGlX73qM0+K9jmE7nCdpMGKubnHsig35F2qyH9Xku6vSWpjY7KuvU7pV7vyvnTx2Vsoi/FSkm273hBCjLGufnFl6fk/oPr8tprP5Rjh49IbjAvTz29VWrlWfn4g/Ny9coJ+eUv/kTefvNN2fXUDtm+a6/0CgpU9Do5MvA+eu8t2f3MWnlq9zPSgpG21JAG8H47ULHUbEl9qS43b94ksIyEVgFnSPZhbR2X2zduyr59+6RI8ACJKhJdzBMFKnq9lvz2N/+PbNk8Jc88vVeuXKnL3Xv3mXiiA/3ixYt8dlWKIM/v2bhhg2yd3SLTU9NM0rHn1LtNgvDqcYICOfZDdEwOyNSp1bRTHh2Iteooky1Sx8sVAhVgJ0qnJfMP78jXX52WNTPj8vSzz8roxHr6frS7KBpUJZcvcq4S5DBNdgWCFajw5AffAaDC51G1XGUBn0X1FYAKFA3I8mg2eS04tvtnOFCBcfb919d/gDh4P3538+Yt3pOIUYFiFZs1BhFQ4TJEtVpF7t68zb0LaxZlsQKQHgUJjI9LRbjJNHWAB5B5cIBjVOOPAKjAdbCIAQ+iAKjA+0pFBXXAmLl79zaNtHG+IeiOa4z3UDXTbjbaBCAAVDhLEueL68a+jjFwoALST/gdmQVmxI25BBk6sG0IVBTKLFbg83gvzgFjHwEVSPSZ0Gr3HXuGwGDlyVl3oy0IYazD5NdCZQcq0KQQAhXhWqAa2xqLQYsqBCp8LwmBCl+bE0AF2IkAKoYyKiD9dD8CfHxsPV5A0QFMDwAV6kGyHKjQrux4AYv+njbbDBbIx4yuv0M+whOg4lH7lMfKSUZ7FPU+NlCR9hRI3/vvAqiA91r4Co8Zfp+LAzwKqPCGnaxGQIYnjxpI6wTm++z5SMcP4SEyvRdWCVQ8kvnDnh5lxqs+v3ZDR0CFFy+jxuxIT3P5laYmh9aitcCu8ZR2tmtFgL/k/6m5rrM4rByfgUHyOGEtwQrebAizjnPmHmBNm3pA+kT1++OCYwwCqPcFXojvUXTGS+UpregaHSx5glFR3djuvG8Z+X82o0JZGJov6WyKc0mNlZ1lodNHZWzV1FrZ3m10pfe1yQDXhbiFckI2boypGG9rkV2lmRS88GMTMzd5HcZfgaefyhlakxv8vqCyYFr/+A6X5wEjAQVzvS/wltAiuu8lzo5HsZzfqxiMLTOq1hHf5+RTpXGjGi+TZVou83xRNCZQge9iZz7yPWyRXe7L6tOpzQheiMbco7QTC9TIF8D6QL6pQATjG5MIJrDBbnpnzWjhHcfCdeD4WldxZgVkPptRAyDeB4AB94m5KzsTtDagwIqCRQ4Yct828A5jtDC/IAUAH9bA4CwOxmPmH+H1BFwTvS6iaZpsgPVp7EAemwxMDknviUpj6b0xMMTyXVyxjgUYLOrLgZcDaA76UBK5L4x/+YzRfBvNoCGIhHXB5jmkwwgaaf3CnwMdT/VC4ZAZQ9TlUtPPt8aROp/wHr8ujUF0ncEzjThYVyG9fzi/SG6LIZvOGTJXAE5ZrEtGDtk52pj5BKh41Kb35PffuxH4u/89BirifT1cpYdtq2kKYSLMSn2AKX206Cc4BxFEGn9EF8LgFWRE2UCFBRmJb9ZzijFwP0ecOxblDO30jNAORfLlr9D9yjK76E1Udk+Fig42mH574oAxBzgBliyjvIa/fWQYmv6Gbz0/tQDAcCQqYHw3QIUusCh0ctZBOxu6lgGjog9GRafJggUknLyY7AV2bIpY5GnCbNJP7PQw6af6Yl1yuRILGV70xwZPVgA2A+vUwwarZpraoYiNxDUfcVzFvW38Wfjuq2eGbYoe9KDgAONPLzZhg3N0X00ulS6K80eBIpTZIOWw2YwCLg8CfDPEuaHgAv3L8fGYUTE+MSF9tMnmciyI4TpDyizvXHA9XvjEOaCw4RrYHjjFST025RxBimajwWJsDFQMpE+tc8hVDSLppw3rN8jI2Lhs2rI5YlSkgQoECBFQYd0rfo36qGmw5GMU3xOV7+H9wD3o9mTu4Zx8+vHHsn7jJhYnt27dGut+0rtNgxwU6bTTwlgwxi5pd1pksTBEsCDQrx/35p033+RYU/ppyxbe87T0kyd3+BzuNbqHUERSzjrq2QAqTsmZzwyogIRUAFS4TiuWH0iE0OfZJKOgaXrs8FHOiVcp/TSuvipu/EbKpxlfe+A0EHn/gw+kUizJywcPSc18VKhNSp8KdMvg/+Uj6afx0Sqln4YDFQO5BEbFPUg/vajdy9aNAlYA9V9BPS4UZWpyKmJIpYGKocWiKB9Yng36nOCMMNAt/JkvaOH4+8/8uyIgIAAqeAzmrJ6UohhqHUEFdDdphwzG9esLX8nFS5/Jrl0bZc/uvbK02JGxsWkp5uEjgIQCHevCZMwN+uKFFnuAZl3aHah7a7zXqr5tWBzwv2vzXTwm6b9nFRTSx0sv+it9bqUNYkUCHyubeq1gHsw9vCe9LlhzXel3G9Lq1ilNt34dgIoOPRRGxw2o2P6C5GSE4/3lV6flwcOb8oMfvCGnjp+QpcUbsmfvNqlVZuXTD87L5csn5Be/+Im889u3ZPeeHbJt13MEKvoAKvoic/fuyJFP3pcf/uggDaQhCdXrIxEsYkdh9yV2CRjWY/1h95/RrrEmQ84OsQHW6KLv+UzWijTPJigLRgUT0Jb85tf/t+zYtkZ27nhKvvjinizWlamGbvJLly5FzxKOt2bNGrKONm/cKONj40xOliDl122Sbu6MCq7TRdVpBlBBs0SaWKMjEbJM+gwXS1Uak/fbTZl/cEMufHFGRmolefqZPTK9dpOaZ0tRYEGRy6msVE/QPdeVEiX2tNMrBCrwnejYR/LjBQzILdUbdSZmnXYvk1GB8QuBCoxtCFR0O1pUxwv7qks/OZMAv7tx4yaBCmdUYG93ZW88X2BfQPoJYwT5udvXb0S0enwmTk41AYR3Bq4P6xNAIXgsoJCAdbDZUm8LSF3R4LAPv54laVD6qcQkHC8U6TFHnFGBogSOBzYF/hsbH40YFZS8swqIF/99n2s12wIAAntoCFQ4YxDNDbgmjNv9+2BU9GwfxxqtMQnkrUqlaoJR4WyLUPop8suxzjsyKsjsUylCdnQEMlXe8ck4AfGJr5X0CeuxUYHST8ZU9LXAwQIFKvB89KXAPbCrHhUma6DvUx+KNFDhgA6OqeyjpPRTu92KGBV+nuGflJasVOT3KP2E8RkGVCQZe0+AitRKH7FAv3WKsPyDw1GEzC94zLdbwTnrcBlmxplfMiT2MN9AFwUIvymjbp19bdxV4nPiyuIHCQ4W1UY9JhqSdvI5dk/DiF0w/KsfmSEOk35aYQo8LlCRiM98PFecYi7RausU1yMUEpUN7YBKDC4AfM3yzQi+yK/TgYW4PVsBzGBeKFAQ1PX5z+Ej6XtkEqzQXBlrIIqk2uRgN3nY/IsY+vYd3s3vjVYwuWYjkxWhCczHxen4KoNY0aRdo0tbQZomG6hQmUCAAT7NdH8F+O1AhdYDCFA40GWd6nrNWqB37X82W4zU2JilxuV6vEj+lnGJ7jl6POv0Zyym8QoAc2/8Y1GeBXxtUHRAAmOCPBl7LfInxB7MJ01/FfuY+1rgvS45hT0R18PmUCv8egOaV15StXYDI5RF4mAY4jn3CWGjAJrgzIwa8yKPZgeAGWSluieFNkwpSONjjHsAVimALmX6uyQyzpnyViajrWxP9eZEFOv5P84fwBaO600zPscJQkTPgsWEBgyS5YDmA4YN5gllrCBcT5WNnsbUzCsI4nLKHt/wuo3hQtPzIUAF7qU2CWpTm8pga9Odzynf770hIvy5+5IAyKOsc6ohwa8D14n4gA2PbChU7wo3dQ+ZQVyeyTJRgCD2zNE+M5Wl0hoF4nEygDL2FgV+IPME5ozeP8/R9F6rX6o/03mCdSorTilyjom/T2WhfQ4gfiVbhvmJ+bs+kX76DoOYJ4f6H2IEHhuooHHu6oEKBQTSQEWsC6mDkKTSJTGELBAk/jmDhKg9xTd7H97w86haelfFykCFQzXRupoJVCQTIL8eXnekaRjeaj+fdOBjC3NiVhj3PkZbkgHTCtFyoiEg4pE8/pSLwIkA8tFA+Vt4VJjxZ69WZbcBi7Po5ESBEx2k1G5UoAKMCnajslsQng1LLAiiK9Qppt5Zgc2iWC6qCTOKIMWSdgh0uyyMQD87lysqG6BaVU3DSMZAE3bvhsRGR83oZjPa9LQbMGeG24ZaI6BBB3ZwG5MbJDS0a1Ywt1lhEkjauaqFAwAj+E6Xp2DHAKRzrKvBN08/BxR+VIe6LmNj49T+hnYz/j4oATzRwBDXh2KygzFefHZZq7Do69eMnyHI8c/gephe9XvU6YZcFHTWa5RX0PsFs3FOh15frl+7IVcuXpYNGzbK2PhEJP2Eq1fJq7hzAQEMihi+aUdPKws9LJNEmzHGyDueI+knn/u9PoGKw598Ius2bJTde54lUOESWxw3AlzqN4LvRWDBORMCFezoCR4oa+lBYPT2b9+UyQkFKrZs28YgMA1UeLDvcwABKLuSrVsf+iVnT5+Rk8eOy89+9jOVkKqomTY+q2aBCmqgsObSGhGj4vBhBjqvvvaajE8aUGHdTs7I4HNpxTV8zoGKVw69zGInO19BF2YF3Ls2NMA8dfKEjNbKsv9F+AVoMOUdPJAI6QiAiovy4O49eWn/i1IdqfHcQbYFUIHn+M7t23Lvzl35Nz/6EQuxOsfiHHAlgIGBYdAN7f9OzIuM5St87lZa4ZgAmcQDPWi8oGhEFA0N45WTnTV9Nef74osjcvnyOdm791nZtGkj6321yoRUymPSM0F3FMsgdZbsrNY5h3N06Sfv2NFrTCbZIcjg7xsGLKSTy5WYEOm5mQVUpMc8PZYrARV6GQbKDHpSX5wjUNHttKTTrku7uyQTU5MyOTlL6acvzp+UsfG+lKpl2bb9eRH6SIicO39C5hZuy+s/+KF8fuYLuX3zS3l671YZHdkixw5/JRe+Pir/8Zd/Lu+++Y48tWerbNv5nAyKM9IdVHnnvvnyvFy+eF5+/Ee/J91+UXLFUekPIKOEuAU7S88K32H84FcKa2/OaGUYGCjvoQVADgLM5GUoUPEP//U/y3N7t8qWTdvkzLmbUq83yKaAzwL+dM1kJCjr1q2TLbOz/HO0WpMODLebDQIVuNcoVKMrDAkbC+cDkVKlynUSc9CBCiQxKDzni2BUzEv94W25+OUp6XWX5Kndu2Xbzj3S6uZlUByVXhdJEBJcdODjvDU5K7l2bx/MIQU5vTN+dGQ8If0EXwywTzAmaUaFmk6rrwfGDesuTMTJqOhjHtQ5uBMTUwRgsXcRiDFGIz7r0k9qpn1brl27xgKDSj/lhSp1+ZyMjmqjQSz9VJFb165HHZRJ6Sct6sCvQffWAvdMFsErZSb+YE+GZtpQ9sK5LzUWpVItc7zwguxRBFRAZpJSEkKT9IcPH8jk1ISM1KosIjCatQ47/B2f8zkAnw8AFe6V5c8hzg+NB0ii3aMCElFYf/FvSE1hnmBzAGhUKKi/R6lU4d4RAhU0A2+ohwjlC9kUYYUYk36K5BxMzsNji/DcAUKH0k/1+QXOD/qoIH6xxydZQOgwo4ZPhUs/ecGC3wH96xwYQ1qIiaQisBcj0RZlebphuB+b96Q+HyX5UTxm8QT8mnBfCVRUM4AKeBENidW0tjA8kM5iV2fvMY9bvs460hNGRXpkhjWDr3TvsgvqWfco/nkiM/PO+9QJPe6d1shC+ad8zsIDPCZQwRnrFT8r5jl4sWzcVgqILObyIr3G+3EcNvSjGcwJlyfO+n4/rgMsK56W3eyo0G9NHt7w4WAFj0FZpuG5fPgd8fdbjGdFRcaO4eQK/MJCWShtNV9+1mHcFT+1HvSa1wUKnlgXrQg+7NoZw1vXtK/Z2symxUoWhK2TnN9pRXwbguCQxtq1/CUGZLPXlKzY0aVwvZiKL9GGu9ijgtI5Ls9lY8lCvBXlvXarxWjsCz3u7YgDwgYReyqsiVT3K/cJxPE5N82fA/JRziLUQq3G0Gx2tGK878UKoGgXvvULRdUQByCcmUQgiJ3y2giiXerqcbBsnAOGhcb2aHgx9jhTCJVJclNvNiNaU5TnsJr7oonRG2HArvbmJP1uzQ97lF9WZpHmspormeQU5a4V4OG5+r0Hg94K98qOV8lr/XxfwS/LP21TNgaNXgv2v1anLcW8ynLrPdDv0FRVATnukzCP99qBrU065srmgDRWrqDHSTyX+mAaewSykdoEiPhW/Tz0+UznLPg95aYgg0Z2UdJ82s9X75vOH5wf4hemyRHop2wEX5d8zinzokc2daGk8bePMZsJwdzIF8ywXJm5WYwKNn9inprUF+RINUZUthJAJJ//vNeFonStscSfEZ07+r0uC4vroWQqDL3Ny4X+GU+Aikfsek9+/b0bgb/7mz8Kgidd7Lx7wMhgukhHP8UjsQJQka5mMCIbFkikwIlH+S24uHjGCCdq+bwEMyWKrsjZDIzyoqI2v5bdoHoELgxk+mnHLX9qidXQr86IWHVhNUZF0GGnMdWys402AkNSQt7hCn/XzUITSjNA5D814Ay7c6ixCZmexEvfEW8C2f03sZFU/H4WWEm9VCkKILtI/mlQTVCiIfXGErsqUWzG3/HzHnQqzaOClEjTTdQbEAMVqq3YooRIq1VngQiJbhqoYGG+jERXNZixKRANB+jQbMr8EKDCCyWadGtxXwMOZTqwK77ZlAYKKzaW2LqZPBvCTr/vDKBCAzSlDKocgdJONVCItUeRmKvMDDY+LZ72OwoWoNiAgCyS4DH2QwhUzMysIVABqSUpuRSP3mQcz+UkvIMVPw8RfQ96PBhzuSn/PLuM+9odic5SdHQCqKAuJoLUvHWEG6MCQMXGjZsEDI8NmzbKhHlUOKPCN17QLx2oCIMJbuAp6SeMkQemejNMvoKP2EDmwaj45BNZv2FjglGBxy4EKvjUo0veghoEtgiG6HXSbScKFtoBmmdH/Zu/+W0CqOCjhGKV+22Y8Xm0cpLi2ZdOr6PBIJ7HXl/Onjkrp1YEKsy/wzwqOLXsGo8eOWKMCgMqIqNRLTK6R4VLP+G5+vDDD8moOHTwkBa8qPmrzyrnJ4NOdHo05eSJzwhUQPrJO4C9gInSbWcwkIsAKu7clYMHDgiMba1/nh1LOODly5fl5rXr8mc/+VOZnoa0jQbHUcPOsGrDkEU16szK6FBZCZgY9rtofUOXG5M90yx3iyRbMxkQa5+5LcO4c1hL8tJqzsvZs0fkytWvZO9ze2R2y2aRflFGRyG9Bu1/LbaBUaFUbn/F7D2s/aH0kyZvKwMV/mykA/UQ0MB7HgVUhMXTld67IoiRvT1wq2MHmfbDSb2+ID2CFC3pthel1b/zhTAAACAASURBVF2S6TUzMjGxmdJPX5w7IWNjfSnVyrJ9+wsyGECqTeTsueOysHhHXn/9R3Lxq4ty8cJJ2bN3VibHtxGo+Pqro/Iff/FTeffNt2X309sUqCitkU4fEk99OXb4fckNWvLG6z+Ubq8oXcHPAVSoP4VCa+RWLJ95mB/GqGC3lBWEsoCKbrdJoGLfCztl4/pZOX36mtSXGvQhQLEda5aCxSozuAGyT1u2yMzUjFQrZem02twPFzpNNcommIukJUegAq9SpRYAFW16VGhhAJT1kjy4e0sufX1S6vO3ZNu2LbJ159NSqk0RqJBCVXpdyC2o9jEL7zk8k0iGlMrOQndbWQ4sFsOUuaYeFT7HSoUSpZ+wHgKowH6OYjvWB4AM+ByBikGfjIVms8HrxjHAYsALXkooKLgvUsiooJl2pcrzuHXztly7rkAFGChIHLsw8CzkI6AiNtOukFGBIoAD81yDo3gL4EQs/YTzjoCKfleaBCograWeEZR+Wqoro6IKBop22oaMCnwPCvH4ilu3bsri4oJMTU8kpJ/i79e4woGKpXqDQIV7WfkE1MaITkL6CZ4puBdgWOA8cE540fi7BKNpABXqUeF7I447HKgIPCqsiEB/igCo8HHTwoBKQzGGJKOiS5mHhPSTbXYOGkSMCgMq8G94gjjYoO/D/IuBirT0E4EKSD9VKgmpSMynpfocx9LjNAKJpgeOOYLP/M6BP8qWfiJQET/zqwW3h2xPK/zo8cvXmQfL2Pse73yy373SOv+435G1LWSORmbn6eN+swdIqc8xb8vosl+h63XYt0fP8rKvWC4fnGV0HkUC1KhZ/i3pexFno8PHI5QGCt/hBWUtdMesi/A9y77+UXl36hRQkI2O4eusycGwU9nzTmvlz+oyzsAGFSgJvjNsJ/AirgMVGh9rk+KwsWfxEoVdrjvKYo/jptU/qxqCD/8OspKtvM77Fh02dfx0Qh5PCvu8MYbNf09/6GwCZWnjP+ZRvB5hHI84AEPtzH80OSV9F6Iv0jXdJXOdRWCj7eftzTtRkZlyPQqWKFCghVQWke26kWvHRtja5KG5dGjqHdcanC2AM9N823wOrNvc4xJWMqzxyq8i9OXwHDueLsausII8BoY5DMcUDQNFZVfCDwnVgi4Y9JqLQ/0AeTV9C405iwuE/4V23KMmYMbFecQJDZM30qI/ARuTQPY9lACLAVxgPsC7C8VtgA7ImbRGr0wLfJagC9j0NLlWbz8CHD1lVgKowGdQL/EclnJiAXjhfi7ajKZsJLwU0NGufYwB2ReQo+Q1l4xFCWYM5JDgYYjaS0fGJ8al2dD4UPEIZbY4gOIPPH7Op5/sCxiWI5bEfNFGR36yiEZFZWeAfQkghnUEK8AjZ0YTiealKOCX6FfCOW6xCk/D1h1v4sS4IO5ko6UZtEegq80t/A73XxskAGrYNRjggWMASEAjCO53qwlFBLBD9Vkj2IF1zmTByHSIfE9iMMXnrsaJuE/GqrJ6goIlKvFEDxQDIHy1cKaSL7IK0uH7XXZNtT38mURcpawVBWJ6T8y0h2+aT376/R6BX/3tH+oKZF2h/vd4m40eIVur/qlARRgqZfw9K4bIiIjjooO+wfORuOMm+XOBAXA6UtJ13RbB5V/kWpGrvdss7Buy7dEpF9igwzha/e2gj5c8eYfEMNBj+LjquGSEgYkxDz+vvwiDaf87gwwrkipQ0ZFmG1raClSgaMM/63WpLylIgf+6ZmKN4i2BCjOj5uLNiBPsBeug6HSocd5sLbF05IwKD5qI7hfy1O/kgs2CS4nrfA/n0wBQAakIaFjDjLMaBQUw80I3Hil2AaXSg1n8ietC8kwDLxpRFiKjsFwBkUwQJiUKsXFQyG7Mihpl0syTQYhuUi79xOOzSJ+TnAWkKAZ5gIqxRdCCwksIVKyZWcvAEXJAg5LRZi2o9U0dmyaOhW7vUHIC38/ub0swHKTx4IHFG+uYv3/3nszDjHQZUKETGgHO1avX5MrFK7KJQMWkbNi8kTJUmNeR9JN1fnSgk14qRRqarm2q56wVZLIgYPzdaPCaGZggKMO4e5HZGBWfmPTT7kj6SaVT0kAFu3poAqYdOMqw6EqnjWKhPQSmg4vzRgDz5m9+EwEVs9u2RYEh5JdwTrh3nrCE6wO+B9cJMAXm1mBUnDr+WcSokHLAqGAC4EBFW5dju0bIaoVAxcTkRCQ55mCCB20KXGpy9hGAilJZDr100DpzDZhh8OvSWjlKep04cVxGR8py4MUXY6DC9DARHncHA/nm6wty//ZdefngQRklpVp7BCmZ1B/I5UuX5Zuvv5Y/+9M/Y+e4Fq9SuswrgBXe+fIooCIMVoetx+E6mli3CB0bUOESbn7LeSBI+qhBNrueSBmC3w3062F8PC+fnfhQrt24IPte3CubN22VQq4m1dq4FIpVzvPR0TEyqfQcLO3mMVUf1ZqMLKFFIK/avP4KAQhN6CyBTclDZX1m2Hg4MDFsXNOgxUp7ENgomS8UAv16B/D7mSebgh5Dnbo0O3VZu26djE1skvpiRz4/+5mMjvWkXC3TTNsZFSfPHJZGY05ef/0NuXb5upw7fVh2P7Ne1szsNKDimPzyr38q7/z2Hdnz7FbZvut5GRTXSG+AQndTPvrg17Jzx2bZvfMZyRdGpNUDMwFsO9xLgIbsW5RQyjEcA/qU0KtkQD1/zjWfI8aowFHYuddtEKg4sG+3rF+3UU6fuS4P5+YpXQTpJzd0pFxetUKgYnZ2s0yN6zoMoAIeCvUePCKUgef3HGs6XgAq+F4yKppSrajWc7+LBoGOXPj8jNy9+Y1sXD8he/Y+K938iOQr09Lp615JoKKD44uUCK4qOFHIl9V8EB4J5svkDQCjoxNMqlmKsy5OSA9RVqDVYdMBpOTQzeZAxdz8PJPLarXM81SgokOgAnMKzD8k4W6mjb2QyRxke+BRUcH71aMCIA8AvxCogNzemDEqIumnalXu3LwZsRGxt4YgAcYSLAr3qAC7A4kw9YYHMVABM20CQ/28LNYXpNlGV78ae2KsFucXpcjzxDlj/9fnGvd5aWlRpmemlnlUONAdMypK0jAQy4EKJtMwVKf/CIAKZYxg3bx9+zaLGPAnyecHClQMhHMEJtqIcdgd2O+zMQTHwT2BnwYZFTDsRjJtEl+ItbhHmTYzryAwmfYGgmhtxR5rzToYP7BK0ACCMWbRz0JE/5xLMsCjguPW68n8wrwyUQ2k0KIJGkKUUeFABX5PLW3zqCCjwpgbmHMA0usLD1lYGQZU4BrxmX81QMU/M0iRjuezF/XV/eZ/PKAiW9o3C6DJ+nn2fvi4QMXy94d7/upGWt8Vm/omPxWlcEOQjmH99JoOrtR9kD4r1cznGqELRRi4WOFV4yvvgs4ExDJyfJU8jQ+bOLsgBorZTp79Lz8g93WXQjV2pO9pQ+kRGTfBgQr/dQiKRMydFECR9QgnxyOosmjV2orqdtWRv6DJCCEvZpe8do+zpcaagSgb44VTl/Szk/BzCSsGPq6UtEEx2d4UdXBboVuL6NrpzpybQLSZ+prSALvmzWfC/dhSRRhr0OGE0zkcnZuxTgImYtJUOQArIrZLXPMIx9mZF5rTqqeDduXHPnnU80e9gYxV3cfBVMf+wX/ncC3uY6B7JkBwxD3qcYActMA6AI6jfoSQ41GvhkiZgcbQauCMOEmL1lp8V+xCGyK5P/J3aDxRFjvZAhYbeU6O/BFjivPGPhhKHGn8qmCMggVqCk5WhN0rHhvMUpMKwtt4rvYMIwdEs6fmjjnWUxCv4cXCfoiwOlAQ5AOsj1muokV0jK8zUeyeW9zkNSMFtFTemQX3vsqlafFd5wX9TExiyWs+jIvhXwNWMUAF85fDcZDTe60uCUxqbc8lr5QJpE17iAcxrjQYN9kx/AmmBmMmqwcw7o68bdDEpqBMyJTSeDlmpjnw57UWzBXE9sl6mj4X/jNKrUXgk94inAbAHdaSymhWUuASLzV9N78SPJNPGBWPs50+ee/3YQR+9bfuUYHHLgAsUhtvkgWQDm6ywAfbmJY5kTlw4HTK5PGySYpGMwsG1koJUfk9ip0sWIu7eYMPERkOiy527cvisuC8HieeizZiLbprTBcb6ujXDBvDxwv5faNNHMuYJysF2Mnv9u+MzzU5DCsBFRq4ULvaGBUxUNGIwIkkUNGQLswsrZtTZXl0k9cARjv6uA2gqNxpS78Lfe4Gu5Zdo5GbhmkbYiVHEu0v77TDxkxPh7k5/oqSCxUAFUKdahRTdFPV79eNTAMI3zQYjHRVsgLFGzdD4vmymGnF/kQnp88nHVtuXiYBgXNQ01T9OY5LEAKAjHWuoKCGzRPvZfEIRt9gXnS7Mr8wxw6HxfklGRubkOmZNZIvFaQ2OmIBkBZX/Pzxd+2CycvMmhmZmZ5mEEINRDv3OK9Rai42ewYslE3CZtyVh/fv0wh0pDoiIygygbWCp85ok7gf165dl0vfXJL1GzbQ6HvLti3sjGUhAj4gJimkAa/qa3pgFxZTrQEquh/uG+JAhTU5aPDU145XFOXXrt8gTz31NKWftBNVZZ80IFJjURZU2OWgQR/ZLN0OmTu+xqlxm3YuQEf+zd/8N5mYGJf9+/ZR+omBC2U1lLrbaRmIEkh+WBsE5w4Lgv0+gYpjR47Iz//9z2UzPCpKMIY36ScWD60A2m5JP2fmp0xMYaZ9jAEZpJ8mJseMBYTuEF3H9H5qAIxhQSfIRx99JOVCSV4+pIwKJjkGYpn6kyDWofTTiZMyWi3JSy8d4DNGc79+lwwE3wq+ufCN3L1zRw68eEDGxsc4Nzi/LDi+cvmKfPH55/KHv/8HsmvXTt5bjKv6b+jzlVz7kuIamUlt8Gz5Mx7uEXHaovfZg0N/9qKkKFh2fT121qCeCQpp7i1k3UhM5CE/o+NaX5iXz44fkdu3rsj+/c/Ktq3r6QNQqU5KIY/u+TEZG59UQl8O3YeBLnXUZWYsEzNgj64pSN7Cnyl4kQSL03tIWGzX9CtIgkOZiFQ+v9KYL9sOg6xQE/7wbuA6C5SFBKNhqX6fng6NJdz/JWkBqFi/XkbHNsgSzLTPfCYjY12p1MqyY8cLkhfMp4J8dupT6Xbr8sorr8qNq3fl1MnDsmvPuKxbu1U+O3xBvvrqhPz1L34m7779nux5dpts275X8oW1Irmq3Lt3Wz47/r4cevkFmZjcwp/1CVIgceVKZowK7VbTl+4j/tLZjNlvHamWzOIPdMGpJq/u5fBO+vv/9/+Q117bJ5OTa+TEySty/8GcXLt6hc9qmckmZI8mZGxijEANwIrx0XHJ54pkFcJDYYldfkVK/3iyqfthTopgVBRgUL0k3XZLKrUR6baxhvXl9tWv5NqlczI2Niov7HtJCpURMilKtXGyENg91gFYqHINTK5t30GnIJ5LZ5RhrcTzin+PjU6SiehyHlgnIT2EZ0b9FJYI+iMBR+Ef5wd5RXpfFAsEKLC3oqACKSy8pqYmpdsdEGjHcUZG1Hza90UYdoOBAaDi6rWrMjExJjMzM+zCa5uO9Tg9KqqyMLfIa0Gjwb27tyMgwuUF42cjJ4sL9Uh6DUV8shux/w3gUQHgR+WWCFQMhF4MzXZdylVtSEBsU19YVH8GJLSIE/LazXrz5g2unTPTM9xvaHBoLFrdc7SwDilKSG9h7O7evcd9HYm2AxUuNVmtVfkdWKNv3bzFOQipRUwiNHhgjx0dQQwD5o12I+L5BesTSTnei/mE5oyR0RFtqnDZEIuXKJWirZFRMSDaH23/4mcshEHojvhk/uFDggfuUeESgxjrMGZSVhWejR6ZjuisJEABUIQFtDgezgIq3KPCAQzEfgvzD6LGBmdx+JzFsXEPf7T/D/51MCqeABXprecx/60SfcNej7PfrfSlur8mN9OVGRXfHVDhcc3wC9Q9TbO5OJ/0budg20vFYqsZ4hRQkfqIF7s1drY2DV9vUu9lTJNuFox25AzRNe/yCOJBHMeyrMz77d+jrRTp6Cj8mEsoJA/lQMUw83POgOh5jWOilQGxFEBhmI9enjbvaWgSvw/xvevVY+/xdZWMdytYKngRq0KlSziKScXSUIyBzQA7GiOTuOZ5GAsNx/dirOayan7t63DU2W7ngW9hqB8AWQquBdetpxJ4E8RxWJi/chYnwCtnCtkBOFCeZ3sjkH+XecFZRzzPnXJLkOIpkxWBuAhxGJoQ4vwIpl4ikJjC3oqX+iDgmnVjRKOA1jBUogrjQfAAcRaaHvPKTvUHQeM6bVhCQ4abWOPiFKBQ8EnliJVl4XsrzrcAsCUoD7lEEL/DvF+4HxqghGN4gZ35P2R/kYeZrBJZJTp5eU4EW+AzaJ4kKgkVeOclpSNsevo6E99rzntj7WDORo0MVpNwphtiAc5XM1h3phAYFF7L8TFxo2g1CNfcnesHmDOsZWjzDV6Itbzor2uMPUcmxUUptaJKq9ILwxkNxhbSmoiyPmNpSo2jNA8jTcUMvfV5cxAKX8XaCcAdexYwnrhteGY9XvP57bWP+D7o/KV8E2VHlQWm80CfHX32dH9zk3D9uY4Jx+cJUDF0L3jyw+/xCPzqb//Yzj4EKcKCuW8uYVA2rMjug5D+XegfYe+xRS8q3kcrsIccK/tHpIfbygrxvhhQKiJSQ7SfWaJkC7StqvEhE18dFPGzMISMex8WuuO3hAfJ+vvqJ9PQYBzBRUSXHHIvlh3eqHzBhq+7UOwVoGt9GFzp31mkNH1KAhUAFNotZVRQ9gmSTw3tGo0YFQ3pldHN2Y02l5gCiI1AJQLQtciFF0VbAhUtleOyYneUHBvi7Ym/Ltraoccu1EaDTAAm/UjywagQTWxrI2O6KdDY2Y2cFKjwa/ZiCn6GQkPolwDtaJyjgxxhwp+WR/PxU6kJmG3DVDsfeWF4ZzwDIUPHXasZx1Uz6b7cf3hPWksAKmBsPclijpQKUh2tRJ0jahimNzrqdMwN2LmKosqatWui6ws7KbnB0qhNOzE0ENWN8+GDhwQrMG7QV6dHBZ8pHQMHKi46UDE2IVu3b42BCus28Q3fzbQdoCJN2wEFNoLGIE9ocO76nmSf4H8oLs0vyIfvv69AhTEqMMZatNaAiPMCxqwOVJjJG/6NAlm3F0s/ocBEsIJARUfe/PU/yvj4mLz44ouyZes2GVAbG0U/BC89aQNEs3sWPV52LRybjrKNzpw+I0cPH5af//znNOWGxjyO4WCSnyfkcgb5JFBx9PBRAypelcnpcZZSNcBVgCIJVJB7JB9//LGUzUzbzdUdqMBzi45aFF1RhDx98qSMlEty8OBLUWGJ5+UJf38g31y8yE7fAwcOyPjYWJTkdK04deXSZTl//rz86IdvyI7t2yn/1OmAjaSdIPpMWAUs6FT3MVupiJCep2Hc7IlSdJ/DBD3NREhRyZnoOsAUO73pfHGTZTwXA8gIFKTb1jXp4w/ekYXFGyxSr1kzLd1uSUZqU1IqjcvEhBZYURgnQ8MCdwelPODVYDsoJmSYaofvj8cqubaHY8cOmzApTBW+ViqorLaQEwXtXAMG0s91ZSAlyfcBVrSkUb+rQEW9rXOgW6eHzOjYegIV504fN6CiJDt3PC95AfOqJMeOfyz9QUNeeeUVuX1jTk6fOiazO/Kycf1WOXHkG/nqi1Pyv/zyp/LOO+/Jnr07Zdu2Z6WQm4ELjly48KVcunRWfvQ7r0i+tFb6A9DIUTz2jjokbwAN4zno+5iOq0kVkAGjL08q+Bzjf8wklGXRaS3Jf/0v/6e89oMXZWxsSo59dkkePJiXy5cvUV4SvgXINwAOT8xMyjTW3jXrWKgGUIBOvkV4CjRVZxdeENq1N+C/8ayUqiOU+YEkUb/bIcAOlsq9e3fl4pfHpVLoyv4Dr0ihPCGDPHwh8vwM5iumL7riABgAKNQEjEiFJmIAx9lVFncZYu8YgUcFJAcp75BjYRzghHYfNvl3MIeQuKuvRkGBCsr5Yc3sUd6o1+mTVYmXAhU9AhV4rgBkADzHZ5H0A6hAknrj5g25ZkAFPCpw61rWeTg2Oia1SlUW5+pMqFHUv3PndiT95Kw9v3dYv8GoUAmQPNkGvqeCUdFoA6ioqEG1dblhL2m2F6VSK3ANxfgAqADohGstoeuQxohgf9xkTIA9GPsiu/wgjWKdgthHkDiDAYHrbLY6cvfu3WVARbvdkqVmXQhUWBPH7Zu3uFqCJSG5AscRazyAfwIyMFRksWEgDTPaBlCxsLjAWIFNDixcKOsv3Xzhczta+5x9aPs+mK0sYURAxRwLCPCA4B4eLD+6/6v+vib+A+m3uwpuUFYir+wNW0/9O73A5vEa9hrs9RhHZ8cgPgBQsTj/kI0NKt9gEpyRR4VKXL6x7/efABXRyrXyX1a7zq/mcFmpUQoTjw+VAcR8O3xmyLdw//vXDVRk3RcWhG0gPR4KC2Hpzw2VQMy86WqanMVGYHnY46nMd9lOuwJDdHkTn52QT5BIviiUJ1g+DxhvsbHA/R/j+sLwuZkNVKRZLMvmfDh5jWk8bBi94Jgo2isJ2uRY7R9ce/UsMabYw6Nu/a7q2qvkC9Z3ZUZ6LhY1BCUaS3RtdokiSgZxvY6BETZoMO+xnxOogJk2WHKIGzT+wZrsazfvedQRb34QgRm5F4rjJqUkY8bzJpUJisEP1/tPkXaWzSq9RDA8dN8t5NULwL8PxfkC1BasmI0YAblYvP+h+VHZzrgnNG3va0Ec+bL6OSFWQr0CrMWayjNZfK2F7ZgdGPsd6N1HzAU5IowRxg3fjxoJPsPzZOd+KZIZgkynXoceEy+CIubnSaltA/+wTyJ3ZZ5CwnBcl2EjHX7Gce3xuxFfOduJebd5UuKc0QDSpvwxQBn1j8J+jZ+j8UEnYnJGD1wb3XJxf/7dqyMxZ8EwYXytc5Uej8YYR+ygcxtNobh+AwksJokAMTJ/AhCHTB+N7X2O4rPRGAVNay5NxjENgFTOAxvnyGMsBELt+cP9c4Nv5LHOpGAmYeOF69D5peOI+0Z5VKt3Rc1AkF5O1dR8ZBlD4XyCPFWZMVqn43OCtcAYN6xncD7H5ulPgIrVRC1P3vO9GoG/+9s/CYpHjuQbEh1dSQA2DN3hrfjPlTG1hVPGZdkKp0fGWyPJKf8yrq7DxzBDNiRx9PR7wgAi+F3iLBX+1+9MFavioGm4vujj3ezvGKhYFoybJM6yzmUfbF5g6pRdu0iR9fiW29+NrjccqHBGhUrcYIFuttssZqwEVAzgUQFfgAh1dq1CnIMXiVUnBUVbFGiQfKPyEgIV7MgzoAIbRFSotO5QMiEMqGDhyIAKyH6w4D42oQZ30G60pN+7/LwQh83HgQhKIQ0GKmVVr5OKh4ARAYN3nWAziouy8XDG6LkWiSAFQkaHMR4wHrph5wlU4OXeFjieovt9uXP/jrSXWlKfRzFiXGZQzCnmpDpWk2KhFKP+HuCa/4WzFHBMFDtcfsL19D3BcL3v5UDFA3lw/wELOwAqfLzZcW8d31euXJVLF8Go2CgT4xMyu3UL5aZwLH9/BFTQIEzHDr+PqawoQgzYUcCA2TS4IWfB78H9Aj3Xun0cqPjg/fdlzbr18vTTe5VRYTIgPidYHIFUU9CVwQ7iIUAF+TwrABWYh+iQtUhQ2i0FKtyIS9e2mMmBNQWalydPnpBjh4/IX/7lX8rm2S0i+RKvk4mIATX4OwMdFEs9EOz3BUAFnoHXXntNJmcwb5W6C6BC2UX6/NIvAuMDoOKjj6RarsjBlw5GZuY+35jPkvYt7Cw+deKEVEsFOXTwoF6HUWOdLQHpkIsXL8qt27fl4MGDnENeeO/iIPCouHhJzp87L2/84HVZt36dbN68SRBHomNJ149vD1SEiY5iHfFa5UCFDruCV1Hgl65+PAZQESX66IhBAZLdMUUZdHvSXJqXTz76rbQ7c/L6D1+lbItISWrVSZmaWS/FUoUMAYLJ1LSPgbcQCH0UUOHrbgIY4HORvfM8DlCRLlittoCVeN8QoGIJQEW3LY1FgIBLLP5u3DIrI7V1BlQck9ooGBUl2bHjOSnmp0QGJTl+4mPp9xvy8ssvy51bC/LFuVMyta4hW2Z3yqljl+TLz0/K//yLfydvv/O+PPPcU7J129NSyE1Jv1eSUyePS6v1QF79wQHp56dSQAVTA/NoSBpjxtdiiVSwR4b3ikAF29dyku8NpFFfkF//+v+Sl195XkZGp+TY8Yty8+YduX79mtSqZRmtAdAtyKaNG2R0YpzyfNPTa7jug1GB5xmF2UYLQIX6WPgzxe4r7AEwT6Zpdkv6nZ5UKwV58PC6fPHFKWnVH8qB/ftlfGKdQEa4VJ2QXh/ghhpZQ0IPSQzWiGIBJshI6nS/R8KItZDrTVcTd3aZhUCFrUnVWo1ACd6LorEWwkdo0o1kHt2DCwsLbFQA4A+ggh4WlHpqcdhhOI0kFNeLPUBZhcpkxB5QKdUoQXX9xnW5fu0aWWMxUIG9T2XVsPfUF5bIGANwcPvmDWXnkZECsD5eFwAGIQ4BqIC1Enu276lgzhCoKKscI4AK3GtIHIFRUR2JgYpGfYnm45SrQqE8n6PcEgzTsW4DqEABX808zQCS3ltqPg3Ta3z/UqO1DKjAuAOoqDcWpVqrUKoPx0wDFYt17DEKVHj3oWptDyLpJ+zp8ArB/cH72Nlp0grJLlWXQVDpiWjdDACAlYAKfCbtzeXHd2B70OnK/IM5KWOfBPhmQIWDFCFo6wk8ni0HKpwd40BFfWFOOyGN+eoNJIy1jFHxBKhYfTay2nV+NUf8lwMqQlZfeKYrFNO/HRqybBj+pRkVQ05I+aDmC6DNXtZ5nMlcwNKcdfeG3fkYGIgaIXw8rdLOKDRoFMyaP1rgzoQLsqddxKBg8cCr+0Pf72sMi/HWtKQ5hMUCqU95UT19sGHnmg1UKNgR26Ynj5bMo6MoKwZLYQAAIABJREFU1bqn7XqYO2gtIoptIdVjvgVaCFUQnfmi15ANMPaCqwNWPsra1W2d9FYsBmMwvO4wTtUGGwUqvFNfvxNABeRRFV3B/7RD3YEKPSb3CQPJE7lRgiwCj4XYPFlZgDl2oCdeLrnDBkbuWPZrzXsUp9ExoQ8FFQzKjGfA9PT7jsYBMOoRFyF+wPsBVLSa2qhGIKHVYvyChgzELNhX2QxmIAIaTBjD1Koq++tG50HdwR8LvA8NHXjxnMpl1keQx3rOR9UE8/kggGT7sNciCEg02ypF5Pm2ARYomHsOr+bnKnul8Z/KgeHkeYx223wKVQ5UfSRUDYMM2H6XbFjk+NrgaDKhboId5lU266KqUZTfhAyGmJ3AuYHSBsEuawS1nNVzOfwY85n1AHgtGPuDdzs0vLbmPjTRsDnG4lZloWhNCi/825kG3qwRPXHGrsHYoAGE96cIF1Jt7uT9MPaMNmKY5B39ScE8Ni8WfE9BfS/wPsSACh7Bm6zIZiRPOXFMB/mUzJT2+tWz4z02Tx3OT5PO5Hkaowk/dzN0nT8aA7OO84RRsZqw5cl7vk8j8Hd/+xM7XSvWUyQSPVEWCPimzn1heMdBSOceBlQo8ro8IIof1OTvsoLoRLEqGOTo/SkgIhF4eELm25utsEqDD4AK7jDLz1U7dIYHVo+63xGV02MrDuWwAHF40Dh8QQu7htLgkC2AqdPVIci4vsTmH16RHmQ4UBGaaUM+p2Nm2g5UwFAbXhXmUWGsitzICDdNFKe5oRgDQmV6FFl3RgVkdeA1gc3dC8S6MKu3gHfLhN2Unvi6rjc6+xSoGJFyFXJPIii+TExOadDqlEgDDcJNzRNrP0//bhQ/5ucf6oYfSBhFcgQpw3kPPjTQUPMjbCyua+n0RWdUeNepf7/TTO8+uJsCKtbJoDCQkfERFkTCgqYXpR0EiEEUDeogSQIgARsq5rcDBl4w0+9WbURnVMBsagzjCMNgdiwpUIFNGEDFxW8uyoaNm2RiYlI2z25mVz1eaTNtAFtepPLv5X2nbrYahPm8S3hUcHlS+QqyKoxR8cF77ylQ8cxzCaCCQY6DBgFQEXU3AKjoous7ln7ygvpQRgU9KsCm0IIV5lW73WDRjx2jQeLGQN003rvttnx2/DNKP/3FX/wFGRX9QcEonjp+DuIgEYHvQ2QSOIBHBRgVbXntlVdkYnqcq1HIqFB9VjdpUxOwEKigDqcFMpxLCGZx1yn91JITJz6TaiEvhw4dlDyLpGY8bkEl/FkAVKCL+OChQ9SQx/WRocGutX4EVPzojTdkanKSXdQzMxMM1HWOeHBmxbE0fv0YRYRhy2f0rGYkwBa9JpZrB+i4t6z4OTPiBvhAWjWeiTvyycfvSqUykIMH90m5VJVSuSZr126WSnUcveiCJifO58hgMNndvBqgIgQr/OS1IBFfSrg3Pg5Q4YX4MIB/1H6W/j1T1TzucUnymNN9SD/doUF9fRHSTw1pdRZl8zYAiGtlaakrZ08dk+pIR6oAKrY/J6XCNIGKI8fel1y+Temn+3fqcv7cSamMPZAd23bLmRNX5avPT8pf/fWfyztvvyfP7ntGtmzZLfnchDQbPfns+DGZXjMqzz2/Wzr9UaSdQxkVhqsNvUx0xA8zYuX8daCiL5LvD6S+OC9vvfn3cvDQXvqUfPzJl3LtGgyW59VPAey5apkG2jANh9/AxMQUJXqQXDUaTTINm60eKewR+EupPhSh4VGB57YiS4s9MrPyubacP/+pzM1fkz2798imDTulL2WpL/WlXANDEIwKJODoTtSElF2FBCqUUcFrwTNr8n9IrDB/KIXXB8igHhW+bzhQoUUAGD83CfqTUVFSvwT4RrQ7MGZUOboQqMCxJyd1HUA8gGsDUO9rMAoK1bIBFdev0aNicko9KgRFhH6HQMVIbZR7T32hQc8IMFBu3LjGNYhgRxqoyBfpC4H9A2sfgAqCEib91Gg1yNAgy8KkHBSoWJTqSDFiVDSXGgZUVKVY0jUbY4DzxFgSqKAck0vHaZcdwCiMabmsbAuwItLST5iEGNPFxgLPrerSTzduJhgVS0tNrrNgleBYPnaYIwCacR4OVGA9d6AC0KrHBA4mhGtRYn90oALruoXEEaPiwUPOT1wnO3dTIacfGyUq1tiGABUoVoVARSytoMwaZPRueO73EtdKRsXCHItszvYkCGPSYTgXFI3eeOEJo2K1a/f3C6jIyrsCaZLkrp45DI973Znvj3KpYA9eMT387qSfss4JMZoX/xkb4zleoaOBqf5qJ0z0vmS1cpmsEhkVXjzXwvvjAFm6Nw0/Kx1yzV/jMvXKYAXXJdO418J59n3Q8sbw71Zj5CEvZ6+kcuQsoCJZQvHcOoq+rOBu/2ZdEoV0jTmZS1iRNpZq0hzM5U5ZQA1OM7wamgOz+1+lY6iVb0y45Swc96dyE19lfkdABVkW+k3uW8FY0sZYTcxN1tbimTjGDMdRY+MQYAule+KR8XsfX1E8TfQ8HNxw+UTKZbFWoEwNymSZj4H6dpnEbw57MPwbitq8QRNv3eOR59DroqtjhxhG8zytW6h6QWwa7ueBfV8Z9ypRxO+n8TWYFGqqrQwOZUOgMK8m5ZpLOSshjv2dPWPNBS4RhD0bDXcAFQb9hKk6GYhQljC5JMaBBPr1+zDuGB8HMBAH4pesB5ApAgNwjQ35sqGP74ABUg5K2aPo1+tFdnyUpCYYaRM01GMxvqSct64XaHDBnAFgoCboKrkVj5MCX5xzFvNRYrVcjqRxyYhxhoSxLVR5BHNMwQbWLVIG3dF9wrlEkrx6pRrLOehr8mI21wkcWD2KoIezj+z9PrdpDE4zdZ0TWhtIy8/r6flzpMudN7kZ5SqoVTrQRXaVPce4x0+AimEL9ZOffa9H4FcAKnzloexOaKztq5O5ulqr6rKtnEaazpBIo4RDGBWRpqB1DiQ6+YfiBLpOZhWyUiBEchsMYIcAyCACT5DC3x0uxv5D/1N1y8OgLF6349FIGg4NmxZhZJgOewKwJPVRUjKjn9nfuG4FC114HRkgiJsUR069ugwH35Y+pzAoWP53FsLpUeE6/zDThvRTDFSgKwHyFpR+CoAKLNq+oWDOeWc9CiqKjSlCDZkV/IegAQXUtPSTdx14Yuubrxe/8Z2L8/MsKKN4UixXiFaD0jg1vYYd6DkGBhbYG0XUJXJcmkj3N31PlJT3u0ys3Uy5gAKCzTFIbTgw4AXr+Bjx7MHf/Np5fFL/VCoHhQeVpIKGJIo1yqhoLDSksdiiD8T0mhmRYl7GpsbYNesdOP6dODd8FoGPJ/Z+DQgUIGk0MzNNU1QvTruRl2+m2ODnHs7F0k+1kUhH0hkVLv30zQUAFcqo2LJta8JMOyosGDU6NB8LC6YIaELpJ5USg0a3dmXQcNymI/5Ex+tbb70l6wyo2LZtG7tCwqIIg0biCgpwsTBnHSUI0BA8xguhekWgIxfv/e0//n8yPqHST1u3baf0E2VU2GEPOZQlFgM9MA3nii1cDFJPnzwlH3/4oQIVYFQUVBbDASUPYlC4krwZATL5BKPiCFkZYFRMTMPIWoM4r60jyGOQgwQEskP9AaWfaqUKGRAI5hCk4lnl3EbQDCmsLjpylVFRKebpZ8H3+ViZrBMZFZcuRdJPzqjg8we6ba8n1y5fkbNnz5JRAYAKgf2mTev4rOEeLgMqkhZt2et7sPb7PU1LjySWzABwCAv4fOqGZJvRMU3vNfp3Aglw93bMPQTDHZFBV27dviHHj34kU5MVeWEf/BLyMjE5Ixs37KAcVD5fIrDmrxAEZVJusXP4+2HAhP/ei4708gleCcCB7TrxLxO/49q6uvJECHquFORg3egJ1qcigYo8pJ+W7tFfqLHUJlBRb87Jjp07pVyZkWajL6dPHpFKtSnVkbJs3/aclIrTEDqSTw+/J8VyX14+9LLMP2zJF5+fka5clmf2vCCfn74h588dl3//Fz+RDz/8SJ594RnZuhVAxag8eFCXkydOyLPP7JLZLRuk1a8mgAodU5V+kkGslZ+MK5YzKhRg0+Qwkn7C2tAfyPzD+/LWW/9FXvvBPnphvP3OKbl48Qrn/ZqZKTIqxsdHKYNWKKEQm5fx8Qk1SM4VDKioS7sDILfE5w5rpIPfODcA6wBOOw2A9XW5efWiXLp0Wnbu3ChP7XleGi0UfyGbNJBSZQyprybcg64UC+qB5AaQmBSk+Lc63Eu5/1Lax6nqmvCMjI6TiRhJD1ix2Jl9AFggrYfjqPRTUebmFqTXa0mprCwvSBt2O/CkqPMph+E0gFaABrhG/B7HVwAVZtpoXmjRn+La1asyPaOyhjl6VOAhycnoyAg9khYeLpIBgX3z+vWr0VqeBNhRKCnIwsJixKjAd9OPAtc+AKOiQeYdwHcAFRj3YdJPSwA4AKZU4UNRIHiE9ezSpUscL6x1/B0L8ZbcspvPgQodo8X6kty7d58ggjMDcI+7vY4sLM6TUeGAya3rN9iBiRhA8kWpL8VghDdGOEtzqalswxCooLwYGkDoo6RzOC40qVxCem30n7EAEwIV7Y7MPXzIPZVjnJJ+8niI8YMl1v1WRxYezpEhkmZU+FrisRtBF7JDhPPDQScHIxBPLkD6yYAKj6ui+KqgDJ0fvvB73z/pp9WsxavpUE/J/ay0XifXvOXvHDYvhh1vWD4WpyFxUWnZZ4M8LPxdZoc985ygYKNBlYVWK4AY9h7NabUIneF+kDlcw/ZilsqTW6w+T2Gckjoit93vWI4qLmLplwGoYBe+F65T88YlUfy5IYiRAVZkgQt8P+aaD3uMGAwdw9hsOpY0GlYUj+KfwBPNf+ZfoRzr9MBqA0HcIOREC2128nP1Oc1/W6FU03+9kYlYx3ML7xLHzHGAI6qVaDUADUHexe0ys2AoevHVz9Yfcz0fBUvinqYMaMHSe8o1kfkAQAJeB6ncPxiSKD70zN5ZD9alrf/U7+bfLVZW+CcJXPHf3p3OfST2w1BQPh43jK97VxAgM7amFuJVygjfC/CAcssmj6inHo6F3kq/Xy7phGOjYY5znl+tQIgeE/GBN2DAc9LkgPhzNcdGjAHGJoGz4NyRt4FNgDjJWQe5AnJ3Z/mrBJN7RCjwp00deCnzoMOYj2yJZlPBEEg+FgqUW+L5oDFs0FcZoJ56g2lzm+WhvYF6J7JZU4EQb9ZzOWauYcjHIrN0ZU644bReq6oGIL8DyxP3Dz4bOBfElyHY5c11HuchT/GOfzbKMO4FkNEyOW6TPFI6ANnyBDzMh4GsE4JSNjZdBSU8x9X4wNhN5lHBlMueCYIZVgvCfUe86FKPeAvGGPcJ98tzeI3N9Rn0tVoBqNgnwkHb+L0ApmBqbT4Zwze36PmMahH2PsxhPBsEEBFX2YOsXhUKOOHlrJVmq81zVskxjHFJ5wyZGcre0OfBcVhjIhkw6Ywbb2bF9YWS2frAGIPpCaMicy9/8ovv8Qj86m9c+kkXfyCcsRyThld8Kld0Cgs2WhYBUq9A81l/o1kQVTFSUhwZDf/RpjhsqFcbWIdyIctYE4nCTxo00EDZA80QYQ47MJJAxbBQLwRDwiuxMcuIDnXDCMATP8wyoELPe+VgPB3YB8dNDK7/PPZriIMuPUYaqABtEBuzAhVLNICECTQMHtNABQ2kjVGBhdgTd3Qhct1fBVDhCzfOJeymVKqcBksAEmCQCR8KFAhKlQpNuZFww4iamofsLtFuP3ZP9BCQqYeGB2SctSmgQt+jwVBYhHGqHoIGPxe/f74hhSGhBnnaVcjbbIEcNjcfF5d+unX3lgIVdQUqZtaslVwpL+NT49TCTp8nxtm7R9wkypM2bNYIzlA0mpqeJFiB70Ew5fRhDQQ79Pl4SOmnqkmaqHm5UhRjRkUMVKiZNhgb+L1KfbgslnbhoDjh4+7FVI5PCqhIMCqsxpgGKt5++20CFXue3isAKkZqtagbwY27KGdkhXp8D4OxwUBanVbAqIifIQRpGLs0UIHItwDTLgJLqwEqNOA/c+q0fPTBB5R+2rR5VqRYjjqkNMDT80FgCDNtBnkRUHGUQfAPfvAq7zVTbo690p5JPbVVSj83oJn2SKUqhw4eioxI+cxYIDsgtVYILsKjolrMy8GXXtKA1sfKM9JuX765pB4VL730Ep8lXwOQQiWAitd/KNNTUwwEayMV2bxpE8cRYIrGdLq2pFeqTCA66CyJEs5wy0kXe741UKGAcCKptUXPC5BxgcSSNBnI1YsX5OypI7J+46Q8vXcnE5Z1a7dIrbJGJFdRvdFozTY9d2cipYCKGIjI6haNE83wsv+lgYq+dKQvRcn3AVYAWFTpp+YS1nn4FT2U7bt2SaUyI42lnpw5dURK5YbURisJoOKTT9+VUlXk0EsHpbHYly+/PCv15hfyzNP75PI383Li6Ify8//wp/LhBx/L3n17ZcvWnQQqLl++Lhe+viAvH4JfxIh087XvDKjAmsh9gPifpvS5Xl9uXr8qH3/0W/nRvzkk9Xpb/ttvjlL6qVatyNq1MzI2OirTUxOyY8dO6YmyirBmVwE+DPIsymJ/7HRhCgiJoFLU4cZEBIB6dZR7TK9Tl6uXvpRvvjwva2YmZN8LL0hldEYeLIKZNiLtFo4xwvUYBd3+oA3bRgIF6BZEkRnJdQX+FTA5LBRJHUehAkkTXs4WhCSiAxVcJ80nwPdHABVghSigUiUgAEYFvrNY0sQe6z2AinpdpZ7AqMDnnN0A6SjMWQcqKuUa1z2wFOBRMTU9QUZFrghGhcoYYE0frY7SDwMFeMg4gFGBccXYOWvPn18ABYsLi5RyQKGksbREJiWTcelLE0AFGBXVKiWKcN7Y51rtulRqRSlYgQhAeK1SYYxBMKkEf5GWXL58md8NoIKyUJTVMEkAAypwjmCM0HB8EUDFPY1DAjNtSGZB+gngD6Wful25AaAil2OCmyuUBNJP+C42WxigpXNEWIjAWOK9kH5yRoUDFXFjhXfE6j4zLG5mvILrtmWajIoQqLAGgDRQ7OsWioaUC3GgAvtkSvrJ40gvZhGQMBYf4kZnbnhMBEYF2Esho8JjCcYPBlS8/vzv/usGKhhwDS/MZ93PYfmSHmZlsDorp4qLQTFTJ5G2WLPNit/xLYEKjW1DqdrMq0sUniPZkIw5n3WU8BqWjVcmUMFPLSupW8Y09KsyoZZH3KOhQAWLmfb9XmgPQCzmNM62gAxLxsVnAhXWDMOCL7uGUtXt1PEIVASF8bgap2iPSt2olr/mbF3pplggmUAFB44iOkngxMeA5tIGqgTxV3hfKRdj1xDLWelF8BkIQQy7UV5Y5Z7pjUbIZ0yixcEZj8d9SMLbqfMpvvPx74LZoAQFzbO0ihsNd5ZZvMfkDjwwR3DAgcCNjlninIITi37jXd92LzQ3Ub/CNIPD76/KPipTAcVdSvL0e1Enuf+cY2vGz8621vHWTUdzTo25vLsc/kja0OU5N4q1iHPQ7KNsE72vWvD1/F+L/wAqtOkskscxthH2WsRjqFm4hFK7q1K2LOqzmK1MChSWsZY4uwIFZjR5EJSy5wHn50bblITGOeN4lvUg7nKJTEr3mKSRAyAKvtg9t3ugzHmNH0PKDeYEcmiME5vP6EWmE4YNAwCXrHaEa6PHJhoBAiUHfF6ljwbS7Wvtw58P9dVAjqp5psd/CvyqhBMK7YhxHPjS9/QprcXmSANHcEwCbibNpLfaAGTL1zxt0zhKjaG9SI/zw7HA9GVsyTFd/vy4X0sUU1A6WusceGbYVErPtCnGuJQJM3/S9FLoa1PUgGj3AyCQX7AzkjgXzcDc1w76opg5tzdI4poBGqkShco2O+jhc5ZAJ6WjAGjgnuBZUPUNrXmpHwXBr0iSKj77J4yK9J188u/v/Qj86m/MTJsori5G2npsl8YVJWRFrFCA51uXAxU0FE1J4ShQoV0PXljPol0+apBXCqoSnw0ZFclfBP8Kj+bXYsFW0KHDEmVgWpqQd4q6GVjJXXZsvc7l45QFMKSD5LhRBnr97C3IOP/wu6NWkNRwWmGWwdrykXRwJjwH/bvROtkZoIacLv0UMioAVtDTYQnG2gpc5EdV+ilMVL8NUOGG3NioKUlgCRgTdAYEHRYnFoxRARonzLQhx4JOUAIVCMSw2ZpJozMpQhDEB2w5UKFgi+teY+MDe4SFLRgyQ5qAhXecT9zFqPcv3GSVAsr/2H2i3+gGnd7Jis/cuH1TmotL1H4fG0cxZy3NtCdmJqRkhW8HV3BtuCcYa5yP0knjBBM/Rycv/BDKlSKLILgW78bUQjgYCB1qdz+AmXYKqGCIY4nI5ctXBEDFxk2bZGJ8UjZvUeknL6IkgAoDhzRw1ADYxzcEKvBZByosfFPpJxs+Z1S8++67snbtetm95xnZvn37UKDCGRXeQYLAB1/eajcZPOo9sY4WA20xRmmgAvcVtFgVn+xLq5nNqND1VIGKs6fPEKiAmfam2VnJ8X6ZjBk6Maz7td2BcbxpnVtQdAzST2RUvKrST6Qeq7Ypxs8ZFWo2DiguJx988IGM1UaWAxXGhEKoR+mnTlvOnjol1WJBXnrpgHaKIKg0iRgOS69HM+2bt26RoYFniQGxGW4jKLt6+YqcO3dO3nj9h5R+wrWjTgUACUXbVgu+NNqRxGAulaGvtniC44bU+mXrY3DcBMDLJS75pZ7s632KOy517ofvRReNfSvXSmOzYFJ1u3Lpwhdy/otjsnnrlDzz7G6pVCZkamKzVGtTAk+cBGnQusD43ARm2lGCEPm+LC9hxAlZsmaVBCqSnXH/PRgVg1yXQEWhX5TcoCn1+h0Z9DrSbEAPOAYqyuUZaTS6cvbkUcmX6jIyWlXppyIk4kry8cdv0x8AgFmnlZevvjwv9+ZOyTN7npeHdwby/nu/lv/pr/5M3v/gY3l+/wuyafNWyeVqcvbsV2TOvfLyQcoPdXJgVJRM+km77XRUtPsuvCHxfV7OqAA4eOfuXRbaa6M1AgF5yH91u/LVF+flxGcfyh/84ety595D+Yd/+FQWFxsyMQ5/hRmZpCfFpOzYsUMgM4RkFJJ4YDXguVOgoimd3kDKlTJllJCAeHcfgYoKnvWOPLx/SU4cf5/P6AvPvSgbZmal0S/JYgeFngpBgSIQHnT7lZDYLkl98Z5cuXpVIBu0bdt2mZqcojlztwsPoCL3KezdDlQ4wwxABc5NJaMKXA/AjERRB80Izcb/z96bNsl1ZFliN/bIyH3fkVgTGwECBFgECZBVPVKbZGM2GnXXdKulaUkfJJPZ9A+R6odMz3zRJ1V1cS2S4E6QLG4AQexrIrHmFhn7Jjvn+n3PIzIiAVSxuopVGWYwAJkv3vPnz5/79XvuOQcazgAqsEnVOQxARUNg9q1m2pB2qpRhjlwIgAr82+4tYFSkkpKIQbZpI6OCQAWkn+j7AKAiI5lUF4EKMiocUEGDz1iMfciEl0syoegB5t1GufcZFUjRAajAegdgPun8nVaWl6VUAaABoELHTX49R6DCCgcoR9UEVMBMW1kT6lGhCVVsLtE/AKEQj6yurcvS0hLnTot38G6C0ZcHUJFxQEWtJvfu3OXygiQKgArIRqEtYE34jArEzwAqsGFF/6yurnK9b/WowHcNsLC5rTUZbesvEx+uQMk30wb7hDILbUJFnt+tFxgntXJZsitrfE6sbPY8KiyesvYYcwLnRbzoAxVoC8ZeIb++AaignjkSSQ6oOHHglS2g4nGbJff7x621raexMdOaHPdZEE34Q1Ae+oQN6ozBOJ8nZ/prW5SNS2PThTQm1YN+CKDC1ubgIi0xfLt4ZuOddzD47tBFmz2j4N6CzaDLt1sy0xWyWLU/mmvJZlsLN+vCjntxV9XNSDkw0d3kTAzu3XNwiX8/t2AeCea1wARkc7i0IU5s3aXSOcoBxNaVYZwUti2Y95yngY5ln1mmiEXY7/5gs9/pFVAIZEl/JrRdFb/5BNC3wBUOhW1qfdChv1/4G68vfwCgwpAO3pPJ13gJb/aJyT/pIPca6dikrnrckvc2B7Bow5K3TLorK47nc4l73yNAQXAXi7X0H/vUA9ZYyOaACkvMoljImAhkabg9dZDY9+RQLbkO2Sfbx9o1OMYAjjkmAOIbBUycvBKT/CpHxdiZQ1jZLPhPuaznVBWGKAsaEENxX1KHz0WC/lzcH3l7Cus3MCvCKn2YI6sHF3IQYCjgfswz04o5IN9kc204teoYxBqoewnHVnCgkoGCzLM4UM3YLfiZSkLpI2fyXOB7oIWKSMbjepoc14Q6chPmzcD9ut4h4x7zTWFcQ1NsxI7wL9OYkVmqONhAIbuTmT9jt7hnp++S5kLs/VHwSxk7TbhoG4DN5gEFtVCQE6X6A+OsctmxTPAM1a+Dn03Af10/INvlQAWO0TA5aoChL89uY4EgC+THEsq0IUjB/kS/u2dm75AbS9pulTLFM8EzIhgWieuY4LvFVjnZsRAAshd3C6h48phj68gfSQ/84j/9tVt5ies50KBd6r8JuWi5O+/4VqCCeTpNADZ/2gEVwZLetvc6MwUeE7UGb3DYhuZvbAQTXKe4b7op0y06wYJq1RrB+e1bzZNZeDOdrtNygseMnSCQaovQmJyWTmY6EdtflqwJr9e0Wd0AqoR6nn7QbP9WRkULUFEpMaFKNoVjVaj0UzNQ4TMqmNB0JomQStFaazVyqpa02h0JDix8pnOMNvhABZL6dqu4a5wPv0dyAlWS0J3B5j1F0ygkhlIyNKyMCkz+CVYmaOUCK1hZee8oxS6AYm96BmG4d1QOINmR6UblqwIDYHAgAYVFXRccLLwOtHDsCXsofv/rv5F0UVorqj2pRw0KKapeIxF5cP8uEyf59aL09vTJ8MgoJXz6B/slARkOZzhpSQDfC0QrXAzJR1utwoR1DkyUY3GFiWl3T7fb2EDaq0ygYunhQ8pkUD4MvLqxAAAgAElEQVQDCQtL+rq9yK2bt+T6FQdU9PXL5PQkZaUQhCGJhEoTyhU5GrUxKvxNpVUuB1uERp0641joNdgOBzTng0ZDCvmiAKgAaLN7zzwTg0gq6eNy4KtjarAKxJg8AEmc7nqlUnTVehp8aiGYSm69/eZr7I8jR47K7NycalYG0k91amgbRdmuqRfXP5AKQmLywvkL8sHp0/I3f/s3Mj0zzedKUMDpdRp9mUAFDMV5q7oZ+PKL30qxUJQXTrzAZ83AGdTRmrJZWM2BDVgE742a373//vs0n33++PMq/cRKDq2qpVGaAxwh/XT+3DlJxWNy5IgCFZR+QkLdWFtO+gkeFWBU+EAFzofr37p5Q77//oK89JIBFSKwnMEYnpme4flQnWuGcToOgm5y7304+flghEmq+ZuZTqtF8zrhAAiaAiKqD2d+f05jIMzXT6tVwjFplFznUaQ7dDfX4NxRbqRr1ZJcvnxOLl76UnbtmJX9+/ZBhEeGhiclnurDjKR3GhjKVRxIqjTh4F6CyjClebcmKwx0aJV+apqfAyq9bmSaz9GZqeGvFTr0mo9tTVLZMfw7WheoYWEc1KtZKZUeSiIWkXwOYG5J8sV1mdu+SwBUFIt1OffN5xKJw8uhS3Zsf0aiSQAVMfn4g7elrzctR48+J8VKQ65cvSR3F8/Jvr27pJpLy9tvvS4///u/lvc/+EQOPrtfpqd2SLWSlG++Occ5/ZmDBym3VW5gHcHGUkEJSyq0VGDoLTdteIgqOn8Y+O7ckDsLt2VmZkompialzqq6lJRyefnum8/l2pWz8tO/elluLdyV117/hEUDMI4eGxuVwf4+6R/ol22zs5LNrZPB0NvTS+N1SK4hcV8olqRUK0kqDVmdtMSi0OQvcT3CmEwme2R9fVnOfnVaisWHsnfPHtk2tVeqlZQ0Ej2SqyAx7qoFE1pdh/5eergoiwvXZWl5RRKpjOzcuZugDphgZQIMKScniHdSdYgNuMVahnUTzxJzAZLsmIPxAWMSusUZFhtgUwtvBgAVq9jmSjIJtkGF7IBKGYxGlXrq6+8lqxLrEc6H79drAFfiBGhSCRhTglFxm6wKk34CKFBxSQ8k6dPJNMEHrCNgHyzcuaMVadEIAQFj6NFIUaKSc0AFfo57MrABbS0Uc5wXYaiNhDoGycrKipQqkIhSGS7MUAQqurr4R4EbZcMAmMdncGBImQ8Bc0orcdFGsCnMx2MFayiBCjAqQjYdYhswKgDekFFRN6AiokBFFEbcIVCB8yE5j40snhsYI/gO2oD2I4ZBrIM5U6tSdc3HONf5QyuNNdFoC5VOa8YABSBHmQbHqECxh0k/4UBNtjTLf1jiCtetlMqytrqmEpFcezUpwaSRm+x8E1IWLACoyOebpJ9wPIGKXI6JHK6ZrqCDMRWBCuG9v7D/5S2gomUtaQWjWteZpsXnMf/hPOkW7ADINwmZNluwDsSJTdgcnfadbeSD/whARVPf/S5ARSdVgg6Jsk5eDf6a1bx/c3vtQKXSzI615X7aXZOe7VlVrWtic3wSRmV+LNZpnCGhz22ysVnc1hjzEOcfV1FujeO+xSviYrtt/9rSTxaF6Z34qgPhmr4B0AmiTK/Q0JMaMhDHeiz8vh+jWZuc1J1o0lzjagX3Levh34vGYjr/2rvBuZmStm6z4N/77wpU+CCd629/529xnSXbA0PtcIDbDO3WC9RkhQVuaLz5T9h6gdiG46au7AWMXdtnqUSOgkIBe8UDKuyyOqdYH+lPNdFvIBv6W/c32ocm7WXjCOuc89TAuuB8CRSIcUxTJt01gY02U9KJYwdJ4YoCFLgXrm3KFEdMh/UJxQkm60M/QMr+YKPocgiogMfxzBFo+9HXWK8JDDBhr8AClRzoeaFJeK5/dfWDVOaMMhsJkriq+TCGdSPfKwwgW4Gyb/oe6F5f13yORwdI6P3oOk9QwMkX2V6VzA4AFzCCLpZUWcEpJqDY0fxe6PvhZLABMqoUE0Abx6ohCBTm+CCToICJt2A4g3t7ziZJ7jA1jWUdyGLXQrtMytoHGILspKW8WMinfYJxh/YhPlSWiD5L5HdUWnvjJwTcHBDkpDPt3SVA5OTC+d4DXDBQx8klmweKvhs6R6B5JsFnc6Y9J4JrTrrP5ksrdMV44HizedOZ3KM76cvhqatsARVPE9VsHfuj6IFf/NN/69qpq4hW59uKwqk2WLTCcKc1oPT+3xaoaNcVf0pAhd++TmBCqMvJCaaDVufmskudzt0Wceg4fjoBFRuDRf+5YINohuBuexpEDkGo4F3TIhzdJLQCFSyU2RSoKEge4AQ8KgBYGFhRKEgE+tWktDlKpFuoFUVXqiUVwbG4l0v8g808aIhWRYGG2jnwPSTP/fs3uiS+B31lVPWQMdAFRkWDG9qhkeEgGWe+DApQwDxLgQq+CS07LkO9VZ8SyZlkUMGIfkLiN7sOuasckz1YwAgCuI16kExx/+dC7WSmUJGJ+CQWESYtWGWbSkoFgFCkIY/u3mfyJbeeJ1AxMjrKRNHA0JAk0lq9iYSTBYk+IGRUQgN5SGd1Oo2abK6x+gGbfjAhaLSdRFVAWdZXV2X5wSMHUiQknobXhxpkRRpqFHbr5m25fvmqTE5OSW9fn0zOTMrA4ADvPU7T1aQDKup8Bibl4I8tVpqYvz0BkLqUCkUm6a1iJJTh0UQJKobfO32aoM3uPbsJVBhwZYE0D4y5ag437ujFgCADHhVlTcQRrGXljM5P6KO33nidiTUwCcyjQpMkCDxU+imQh/Erg6iJj3kDZnhRuXTxkrz39rvyNz//G5mdnVKJKwMqaG6moAWSgQAq3A6P7fjyiy+YLHzxpRdlcGiQgQmC0WpFKz3QTiQQUX2NYB4BzqdnzkhvV7ccO3ZMZVFc5Q3GrQWgTHQVi3L+u+8kHo0QhKCmqKP4B9vSWp2a7Pfu3ZNnjxzheMd3+Q67yiP8/sL338uJF18ktZa9GVcewtDAIP1KKjAUY6/RMSBggxknjOGtmbR7m7ZOG+G2K0vwvipNO5vNkQ3EKqGoGRKq5A3f8YiCKbPTk5Q/s/cE5zagqxUw8K+LOQvBJ5gDVy9+J5cufCMH9+6WffO7+IL0Dk1KV7pfGhF4B+g8zOeE6v5aCFR0BiWsiiYED1qBiqb2BGDHRlDCdOQ7Li6ebFZre1o3/T6QgUqs1eWc3Lp9TXLri9LfH5W52SlZWynwfSqWizK3Y5ck4kNSLkXk7NefSiS+Kr2ZjOzYeVgiYJ40ovLJ6bdkZKhPnj3ynOQqFcqN3bp+XvbtnZRErU/efP1N+bf/w0vy4Udn5PBz+2RuZr+srFTk7LfnCf7h/RRJA3ZtI8Chd93pvvg7bBK5U6pLrFGXc+e+lpVHD2V2dkZmtk1LPZ6WerRL7t1dlMtnP5dH967LyVd+Kheu3JTfvPUxE8sAZyenJvh3X1+PTExMyGo2yzkCc3ZXV7djGxQJVBRr65QkSiUz9OnAXIeEP5MdNZGL57+Ve3cuyM6dU7Jr57zU65B46pVIoluKoNjHIlIu5cleyufX5N7dBbm3eFvKxaIMDAzL6MSUDA2PS6Z3kMghMM14RDdrmB9BpzegAn0D6Sx6AtWwyYUXRIrMRHQL1jZ8D2sp/gZwjfVsdW2F804iAR3hivOoqJFhgmv0DfRKrpDndwBY4/v1qlYOYp1LJVJNQMXQ8AA9KrDGVMj0jZLFgXkMDE20F2v4wsIdTa6Dj4O1z1VtAqiI1YXt1iIHBSrU9wnvobIYkEgHU4CMR/iOrK1JGUyLLp0v8cH1fKAC10b/AJgHa6K/f0B6enp1E+lM0LncQLcaa7iT9QKI4AMVltxCuwDidGW6CJpgTr3r7guAD+YQtAEfY1TgnjFP4cYBVODaaOPy8jLntJ6ebleFGG5wLc7wAUeb3+y9sNiEck1IJoEtC3bEWlaBilSSz6IKMDyoaA3ZGhgkeBp4zuhL3zuMCS7P3yLcoGsiCNfzgQrTYSbzaF1BJXzfj5/wjKJxke7uLjk+f/IvFqhonc/bJWjbrREd1wHvF8F8aT4PVvzh5lKuzR7Abl/94YAKLMRhItoAk808J/y16fdhVLRbL9wqsqHrtM5B98ttIZenBCo2w2L8NSxI2PrXd89IjW21NSo1E4KLnSqJO9+zq5a3+/Mq4DvtYK2YiHOOU0+gp1VVE7ow/KVcixd3tApSefVQTewK9ndEk7EGCLQDT/z5jv/2no6CuCGzol0y2JfbCca2eziaDEWiWqv9cW5dX9ozKkKgIoSN0Ibw4/37hwAqNIjl+4k9l/aPVssH8zFB7LCy3FrAVL2XAFUQSUELxv7OuBv/VhlnzRuZAbjPiMBl9T5Drxn9mbGMXEGZq7gnO8OB67ZGMcnOwaBoKfcQLgkcICBO6cGSxMbusESxnsNV8jsWIPbIJjekRUp1KVPuM0LWJu4TDAn8XFmTZhgfvuuoelcQQ38XSEUBtHcAhcogKcDPsUITb/0eYiLzJkMbWdBBiSb8vByoFgRIsXvXET/RANybf7XYD89Ef47YRvd+2l8KXDgmDYrHHLMCazvaBakklYHW4kV9pmBUAIyDrwZiihoLKilTxH2rvkPYlyD3gPcaey/cC/0vUfBQU5YJgRgDFLgJ1P8oY0XHhPk2wEtM4wBlrVg/qfSRV3QWvEAh+Go5IBu3iDmxD0Qckcl0s+CFYIN5fnhvIVpEeSaCiK5d3Csqk8YUN9Sr0oFbru2IQznfVnC/mBfAsoGkp4JVJqttUmQBaOTeI/P5snmYwBKZwiqNp2CJF9f56Vr8Nj7xk8fg+E+y7G8ds9UDfzo98It/+m88YMIHKlrbGGCWbcKwpwEqwmObpZ+cniQv+3Sv2ROn+b3Iublqo3OYFQQmrgpNg1APqGia3DZrif2uE1ixyZjwNgJNQaR3quZEXjNAYWfWe3aLq3Je3a86mXyHx28EKnRz2p5RgSSAx6gAYGGG2pCQ6Ib8hAIVFkSaZnPdGboTqMCCBd+LUiFIcBjFlguBO0cnoALnxya3HVCBRLYPVNj1N0g/mR6g93jsGAMBsAihwtwSD+gTJPzLkJ7KaT/EI5pY8DfZrM50lQ0MBBzVNRqt06wVRm1YpBPpFOWdECYuAahAX67npAdAxcgoA52hoWGJp5OSznS5QEirPKyNODfaif+jX016y5INVg1kySskGFD5OTw8KPF4RHKQfnr4SLW4k81ABTLOSGoRqLhyTaYAVPRD+mlSBgcHuKiC7REHFdSxOqCHqYGYJudtfGmVgtH1tWKpCMkQmoma/ncYSuO+1tfz8t7p99SjYu8e2bZtlvIqFuBaHwOowHXM+No0HwGE1ap5jkcNkK0CW4O9t954g4GNARXC56ZAhUk/GVBh41nBTN1ARSATVI/Kpe8vyvvvvCt/+3d/KzOz086LQyteaUrG6p6IAhUIyCOOblutyW8//5zP/OTJkzI4MhQyKqoa1AG4unLlqiyvPpRavcoEHDTUR4eGZfvcdgZbGH+oTkVgOjc7K/0DA/w5nvn5784Jrg6ggka7VoHr0r1IWBlQccTzqGDg70zUrl+/TqDiRTAqBgZ0pkEf4D4kQoBtYnyCkjjcXDLBqEGgD1TYCtDk/9Mp67HpUqoyhjCw/fzzL+T27QWJuapcBI1gwqBSGRXeo2Mj8m9+9oqMjg4HQEUTyLXJdZD4BQCB4px6OS/fn/1azp/7Un5y/Lhs3zErkozK0NCEJBLd9E3AHGfVT8xEu4+fXLF5PtyAhKCDHqcrkf9dv4ntvteuX5tuy9usNq0zXvtagRtrM+amUr4qN25ekVvXzwqUwQ4cmJf1NeitRiRfyMmOXfMSiw0QqPj2q09EYivS252RXbuelUjXIEHqT959UyZGh+Tg4SOSr1Tk5u0FuXb5rOzaMSADXZPy1utvyl/99VH59MyXcujoPtk2u08Wbi3J5ctX5cDBg9I/MEIpqDq8jjo8M38ta71Prd/DZkeBiq++/Exya6uybW5WpmcVqCjVE3LtymVZuHJO1lcW5dRPfyZfnb0o7733ufR095BNMbttmkAvEsYjI8OysrbGjYqaaStQAbYBmHelOnR3uyRJvwfo8BYllYSJYUFuXbssC7euytjYgBw6dEgi0aTkizDm7pFYIiWVKkwgI1LIZ2Vl+YEs3r4uKyuPOJdMTs3JyOiEdPcN0L+iLjF6VGATjTePkoDRaMCoUNAUPhrdXGPA1sJ8nUqmJZ8DUKEgPOYLJMzxfQMqVlZXOBfGExEpFspMuoM1gntEl/YP9PJdwx8wR9Av1XJdEskEpZ+QoIdk5MKdBblDRgWAikFuuMtM2ChQAQZHdj2r62IiEQAVeI7GGrOK+1gd/aJyk0iaWLvJtqzDL2OdIAn6HgyWRhXASpYygKkMEvK6Qcf6jXgB92xzQjablQXMJ7EEgYrubkh0qaa1jTusrQZSoK2rK6uytKxm2hZvoN0AUtbzCoYYULG4cIdtNsAdQAY+2GzbdxWowHrRDFRgLffbinswUMDeV4sX/b8tBrFEDlevmsYK66trbIuZaWN98GPOoNrP8bINqDBwgbOVSxAZcdeSVOjTVqAC7CgUeHDMFYudgQpooScjBMaO7XlpC6jw5mrr83bTYOscaMf4id4N64kb2Ew4e9KIrqRJD/cSZp2Bik0X7ZZfWiW2l5SyKv1NzLH9tfT3BSrarYXcR/n7L1tcXetbd4K6k+rgCNGBUbFZL+lSrfFhsK57RtStz9H6I4iFzV/BFe1suFaHxdOqu7XqW/fsmvxv/wlcFTS3HH7HyT7jW1gX+WuXRG/q1w45/CDNzyK6kIXhxyeswm7pW86FLuGoY1i5D7wbS+J7vt8BkOHdnl7bMq16MI2J8VMnWfMkjAq7vo4vK0b5AYGKgMWiQAW8P3T9MtAgrKxne+3SHthmkrz+O2B9HIIMZqKs+xffp8LYF6wid7I1QZKa13G96ZkJt7JOuGczc+6Y2x+6sUf/BxuLzoDanm+QYCfzXJ8PJaXg+QBwAmoFTDo7lj1ll0ErhCmy+j0gea55Bt2foy2Mn5wHhybR4YNQcvLOOo7AHDf/1XIJMbDuv838ulJTY3Cr+kdPWCFjBe8DxqjziyKjwVgyTZ70mpQ3NguLLVyuyLAvjneAIyjccD4K9jNjzOIcKKogo8QVjeJ+sIdWHzNjAUV174z3Bsbb7LuqMvDN2wJyUWB8ur7Win/tfxb3GksmMH92S4YbC9bHxoQAuIa22Xto7A3mgdoAFVQTiKEYR+dajA8FSvS58VwOgFDGbPuPzR2B74efg3NMVPXJ0IIUfJRVYvOIjlPstVHMgmeLvkQ/GGMf7w9iHEpmunFp67KtryEI5dioNLQ38DnMmTbtlbeAiqcJMLaO/TH0wC/+yUk/BSyKMORoF3w4u9GmWws8Jhi7tUZvLlll3/ATLBqd2FLlAq7NQAo30z0BMrHpIWay1TG8ssY+HsAIO6IZ1tRvtvPm8Luu+fztdUG9sCiIzjwoZ0MT2wAhQZcaSOECLR6qFEeXVWwZsi7R2iqP4RaIEKgAKl9mgAJjXpN+wuYaiVFIP4FdQUPtQl5iSFJ4QAUmZ2M0RCJAqB2jAkBIuSzFopOMiCc8M73NgQpLQhtQgYXfGBV4Kj5QgZu265tuN5K9rLbmQhuaQNuChONMVskHKiygQvUAwmfcCSWwsuvsHzUP1QoB3xzSFioyK5DYpcmSk2hAZSYAiHhMVu7fZyUATEp7unsJVKDKADJWADS6e7XSXYEHIPjqBYJrAmQwgAKBCOmQNJlSGS380YrXeCCvAA35gYFePoe15VXqV8aQXErDlBwLptJ9AVTcvAHpp2syPTUtfQMDMjE1LqOjI1rVEXeMCladCIEc0DiNemlVRVrhoFULRjllVWwHoAL3WiiUlFExPCrz++Zlbm4bgyyObpObQNAedywgVP+46k5UixZLBalWctwsICmytpplJSyqnFFR8v67H0p3T48CFZB+isXV8wOZ6QYS3iGjwoAKY4boJgiBXFQunr/ggIqfy7a5GVZCs7qGVaugBauUB8ZJTVC5ohRrBIfwqABQ8dLJl2RwaMgxKhBw60YRVTBXLl+Rxft3ZHn5kVbBrq7J6PAIQTSMGVbjJvV5T01Nyfw8EsdqDHv+/HcEKnCPqPypOokoSyoRqLiuZtoAKvp6NTFHqrsL5q9fuyYXLlyQl06e9ICKOitpGtW6fPnVl/LKqVMyPjqmgSSYU66KRqu31HtEQZ6nhavDqStMwigFGxI1t27doixKxemt0hTQ0WiZUEwlZNeOORkY6GvSj+dM+RiQpAHGjBLNJRZpSL1SkK+/+q1cu3xRjv/ksEzODkg83iXDQ9MSj/dIvZGSRs0ZqkVKAXhsyUR/EvYTLs3/bp74/U1jsNR683TTOTdbHDdhVASroldJaX1NYK0Oc/aKLN65KA8eXJd9e/dIYb0ilWpJsrms7NqzV6KRfgIV33z1sUh0mYyKXbuPSCQzxGr/j37zmkxNjMqBZw5LrlSVhbv35Nqlr2V6KiXTI7vk3bfflROn9snHH38pR48fkpmZ3XL92j25ffuOPHfsOXqDRCMZKW8SRjwOqGCtXqQmsUZDPv/sY3rQ7Ni+jdJP1WhSssW63Lx2Te7euCCl/EN5+Wc/k08++1Y+/ugrJq3BoJjbPstkPJLrAwP9sry6yvcc3j0APcslJMWxHhal3KhKqisjyViSUgTVMqSfGnL75lW5feN7SSUjcuKlUwQaKtWklCoJkViXIE9dq65Tduza1Yty/+5tKRVyMtjfKzNz8zI0up0rEBxrkkmYi0clkUprIgGOEjQ8DOUHuMGr1cgCAVABU0RKLKW6OPfgA6ACa4gBFfAsMkaFAhWQRSpT+glsL5N+6h/sJbNS2QkZrsXlYlXSXWkaY0PSCQDN7YXbcufOnQCoAEG3zFxEM1ABGSCAKHfuLAZVwjS7BssNVfeYdRuQHlPJSTJHymVel4mKWlHyhSyBAdwL/SgIVKxLrYF2JdU4s1bj941RYRXJ8IJYvHOX6xoAKQIVlJSIBVZfG4AKsBKXlwlUGFsAfYr5dz0HjwpIWymjYvH2AtuM62K8Yr3HnIjvEiyIQNMa8mbCmKuZUVHjfeKYcOPvSz/pm9wKVvjrJasmubCrnvO6MSocq4FSAy7OsAILzqdtgIpg825V3kGOT9cu9JMBFRgfuC81J9dYwYAKK/SwNd0KPWJJADgZObrrBNd9HIdKWDyLWBSxjALW/jz+uDlde+jpCqaa2eeWvveC9mC/4RJ0v0OCuiVA7/jfIOGxyRfa3Z2/NLT7fZCUDrONmrjy++ox3fZ0t23oiAMsbC/yuGsEexoPz9/0O0/+rHnkJswJvlsbdlJWjGPX8fbZHdbjTmCSjU3rRxtpulvTseWPOpN54s8pL+K4rMG/Nw6Sds8I5wRrztRbrIq99dimcEkRmqAgzY9NLBkXxsyqYW8GsRv60XtEPjkFVdd2Tc5FXiW+Pwz0ldakL+/BMU3C+9Er8j6ZKHbsXieh47fH7tk8KWw+ZYKW0kGhxJ29GgbqaIJYWejKHjdGUqjaoE1tRWn0qVocGM5h4XGsmqcUkSbW/XfTvydjtFg7gvfXmqAUC22DmXh77Qlk/tw1fHaFJZWZiEdi2DO7DhO54ZjwlRVsfJiEVrC2EJRzeXg3xtW82MlCNcWtepxeV/tXvRX06WJtM08FM1lWWSJliyChzfU1mWABmXlgMR/g5Hls7NSr2gZU+2NdZk7EMZe4f3ePxqQW2e+BRKS2DcfgOtgP4/fmhxHcu75Ayl5gLkJZHzpuI9xLY1/uJ8oJXtDz2tZXGDNXuM8EQGNjx2cUmRwV7sOYjThelQM0v2V7JlUKMEk+x7hwHhLoaAI1AEcQUxKIVDNsK2iw52zxlMlTonDNmKw+tKsglwHkLs4Ci8n62sUW6CMNbjSn44899ROFETfkvdUnBLegQIjz4XCDzObPVnaDMXRMMsvmLlxS92DoIwXPVOYa4AQY+ypFboWqFnuTGdFQRlnwXAl8KtASzqWh9Jo9A4BP7i11Hp9qYr/FqHjSKGnruB9ND/zin/77TdvaFEO5SZUC5l404sWsG14u5WraH7uUd9Y2Bs4bG6STpC7cLnHfxI4IA0dr16ZARfMMsMn9u7OEzGZ3rH/29kbWXpjyxGOh1ejVN7fWheVxwEbrXbfrBY/6akBFEIBsDK810eoFTTYGzEjXSQaZ6Y9WXCIJkFdgwiUnQo+KPKWfjDpnnYMJXBkJOrYoGMNzV6VUVBNOVC8q+q+VnwZ2cGPqNu22MTfaHwyukVQw6SeYaSPiwSJGzXEvWYnv2iJmiXskYf3KagY9DhnHMbhf6I5b8sDAGwYKSDS7cVuv1mjqjf7AOaxS0mdYWPAAgD6q8Y+rPI9IA1pQ0IIsFHgeVNAj4QVfBgAVwyMjks5kJJVJO8MmRe+RZECbqMWdTrMf0Xf4W6sm1IScyfEaku4qk2GBd70Bk+eGZFIpqRTL0p3JSDKdkjhooqw8RsCiCWEAFdcuX1Wgor9fZuZmaSaL1x/a6DEn/cTArKaBGSoKeH1XjeAzKuz+Uc0LVgU+9nsdNxpgQBMdQMXo2Ljsmd9DTfhUOh1sjqxfowkDcJSCyjFSLkuukJNCfpnSI5BXunLlGvtrfHyCFdCffHSGCchnn31Wdu3eI1UkV5AAIVABcEMN1G1cWt+hb9T4G/rnMXpUnH7nXfkPf/dz2b59VmIJ1aysOqBCAzFNqNUjOgDYB/W6fHHmcz6bEy+ekAFIPwWVQVqNUa2oDFmlXpYa6bgiH3/8MUGEnxx/Xqt3kBByGp9oK5JefI9qNUo/JZz0E9AnMqVQeWKVL/CouHZNHjx4QB8LADeszEHA56qoKP104YK8+OKLlA4j4BjT80OzHO35Nz/7mcxMTet1ubnQ4LYSCxwAACAASURBVDPm5nOf5v9YHPlxM6tjxnBf6v5AssQ+tr0zLfc4ZMzgDeJJWzzuEvi9yjCp/AyZYBgLUpePPvpQFu9ekxMv7ZexsXHp6hqQwYFJEYFPDvRSI1KPYFxrS1qBio3gg9Lqw2uGrfOP9c9jwKm906R8b5KA07vQjw+M2P879kcU1deaMikXHsry6oIM9vVLMQewtCBr+VV6VKTTo7K+Dqmmz8APk550SnbvOSqSHoBOmHz41q9lenJMnjl0VNbLFXn4KCsXvjsjQ4MV2TmzXz5+/yM5/uJeeffdT+X5F4/K+Ng2uXzpNjdr+/fvl3i8Txq1Lqk1+2U3Nbs1AeT3HVc7bsCqBCo++fh9Os7v3DEnw2MjUokm5d6jrNy8cV2Wbl+VSGNdTr3yU/nks2/k668vMmE9OTkpe+bhxwHZn5jAFPregwesCoOhdToNP6OIrCyv0o+iWK9KprtPEmBpYT4ow4NoWS58/6006mty+PCzMjIyI+sFbLIzUgTFAHJ6sbIsP1qQa1cvy8MH95mc3zY7Izt37pRU94DUY31SAgDaiEo8kSLLAsZ+vN8GWH8llaxwcgjGCARQsb4ORoWaSwKUhawc3mcUHjDhn+nmxpnShPG4ZLNrEsUYEKwhauaMSkJIP+G88JzIFQFUwCw5TbYePCzIjPAZFQsLcmdxQYaGBjiHMAmAeb4BH4I0GRxgVGBNbpJ+op+HSkNyM094OMJKfBQr4Of42xgJ5QpAoix9oOhbgTWvBpm4LH1+0l0pZ6gJsMWxHZy8JM4FWaPbtxYIVKCdXemMSgSw2lATCGiHn3R/9OgRz4/roa32wTps0k/0qID0053FgFGBuR79hs2ueWwoC0ErWPNFXRvNowLjG2u9xRY2TwegolfB578YNu+x0MEkOgBUlEoEvXFOAidIxrX45wTJM1dobowKY3+wP5ynBvqHlaoAsB2T1EAJ9LWZaduzRJ+V4dviGKmtQEU03pCBwX55Zu4Y2T8oMtgAVLQAzr8XUNE2p20/fPKEt06yT7LC/B7HPB0qsOmFgqb6laxM+Hb4Wsdrt9+dtT/cgIoObIROLfb6tR2I0qrCtGHvZefttJHEhNQ2m7+5k6KCBC3FD09JPfHXr6Z/B0DFxk55yku0JMm98wUmus3X8Iex32Uu3/3EA5jSlN5L0fScvP72r4GiMtv3Yb2ilJSXK2i9OMdDh3dYZYdRAKDntOpsX5oqZB94hu0tcmhg2Lb76P5R2eTc87hiKmWqNI+pTkDVRqAivFI412sCNkjSM77Um0Yi2CrjzSjYzy1o/2zsoHbtMbCJMYXzrghkcJmsVSajJaS1pWHfKEbj5HocM8XuwV+/7PvMGzigh3t351cEhgRlFxnbqPwSfQM9WR8ritL+0/eQ1ew0L8Z6rH5/+LfJNZHp7hh/BAK8KTvwQCA4pftZdBtloJC09xQrVI7XVd57EmyUV6I/lgNUcH8O7KCsEEGWGgtAbI8cjF13fsRjKBhhQUYMvlgAJarOuFo9NgjIOJkzxGsKJCiAg9gH14CMGtrIAgU+JWWQ6GU2jmeoIgQKF+4Z0nTbsQdQdINrWLuZ1XFMTL6vzqsSnWbsBibwzQ/FXTbYj9k+Ds8JJtUsrFEJaQNhUTDbnAMMZcr0vC6X5aSveG3nqYJz4lyW4zFQRY2vtU+ax7E20B5zs4Rb+E6qvDAKDvEcTcJJY196ZnqsNlOZMR9HvguOOWdgV+v8rz9XTzTEVFtAxRMvN1sH/lh64HFARcuyonPkHxWosMnBS6jgR0F5iQMyHvcAOkZurXOyyTy1ntBADPd3ixH1Hxao0CBiYyjx4wAqIP1kyX7r1QCoaJV+qlYCoAIJeSwaFpQ+DqjwpZ9QEd6LasSuLgbCuJ4BFXZtrW7XBL8BFaj29DfwPpiB4xCEoWIdSZPgu2BTYOGORZkotmQugihUbGLjjQXZkgkWEHMD7hZDWBRo0QIkchxQAbS8VpFiPi9Lj5Yo42FABbwqkpk0E/SWcMJ3TeoJ7cMf6FnjXUG7kfhuBSqQzAmDftBKIb2Vl2itLql4gpXykJgywMcHKm5cvynXLl2VmZkZ6esfkKnZKSac8FFGBZ6fgiBIXrcCFUa1xY2rnq3eP6p54VPBN58/D1LMDnQpy3vvnpbR8XHZu3ee14d0hCWLLGAEo8KeEStmoKOJZ1gE+AO5FLBfcqzORmJ5ZGSMybo333iDki6QRdqxa7cbP1qxiSriQh5ARaUDUIHnCEAjJhe/vyjvvv2O/N3f/wcFKuI6lnGNchmSXBpUQfoJOr30/yBQ0ZAvznzGRBuAipBRgQocrRqiOTYqiGCmTaqv0Ewbz+zUyVMMihCQITDVYF+1RrFhwbO4fPECk6QAIVhx5BgHlnTDWLx29ao8fPiQx8Bw109O4X0BUPE9pJ8cUMHgEybLkCArleXDDz+Ul0+elN074d0AzVJsKnTOAlDBoNgrOPz9czhmaqcQAv5UG67ixk08rLLiJhPJTZMW65SdeOyiQn8DvMXUH41G5cyZ9+Xhw8vy/AvH6ReQyfTLQP+4CIAKiUu5Xg5mctug2VVagQomEF2io9WjohWoMMDVkqOzs7OBbMsfAqjAJgeMCvRntbgsa9n70tfTLbksmHZ5yeZXZfuu3fSoyK1X5ezZz0RkKWBUNFL9TL6/9/ovZXJMGRXVSFLWsiU5f+4j6e5ek307D8lvP/tS9h6YlI8+/Eqe+8lRGRqckLPfXWRV+575eZF6tzTq3VKDdnWHLOCTARVgVNTlg/fflkQsJjt3bJPhsVEpNWJyfeGBLC4syPLiNelKVuXky6/Iex99IRe+vynd3T2Untu5cwff73Q6xSTqvfv3Ob77+4bIUKhWG7K6ssakfklqrKbHuxqpV2X54R25ffMy56SDz0DKbrfkijEplWGinKDPS7VakPv3rsuNqxclm12XwaERmZ3dLjPT2yQNaal6hP0HNhFANG76nSkk7z+ilfIEDF1SxuZ9k34CowKyaGA50seiBagoV3SDjHlwbW1F/ScjdTIqwCYpl6pkjWDuGRjskzyAinyBVW0ADABUsMjAARWQYqP0050FSg4CAMAzNKAC8j6ZroysZdd4TiS0b926HSTkcS783Ob9eF0oWWXVgfhbPR7iUq4WKP0EfwqAHwDMI/UG12Z4x9CjwjEqfKDC1moAFZA6hH8H2olnynXGKvLaABXwpwCri6bgKJhwHzIq8jmyS9KJFJ+HARUABhSoyPHeyP5wRR1kIcCjqaCyUOZRYf+2RI8Bl61zhL/p5uzoeWYF4axjVKytrLKvwDLEVGpSFBuSpp5HBQpEDKhgbOOkLCx5xGSKS1JYWxEfWaxifY2foVDBByq0slSrL2MEKgbk4LbntoCK1iXqDwFU+Put5g1i89X/HICKTkv+Jv26WfRgUkRBEtNVrLe9TIdrtAJGAQDZyQOjw26x9TE2taHT/XmeBU9yfMdu8uRem86DuYVyqeFPrT8ZH7bpKCSBNTZCAZH6hW326QRUWMIcyxhBevPvcz4IzQWZnlSSsVh4gIIXnYAKtAvxOZPD5i2Ar5FdYeX3nUECPwZsd4+Myd2DtWO1GM+8STTBawV6QYV8U8+G1+8Eitm1LWZlsZGT3MGeAnM4fmfGwQbQtbYZ+1N8D1X+PJcrmgjjXL0fSvE4RgOOUdkm3a/b+sbEr2O/EEBxckoGOvgFSBiXABdwDM6bgryyk5jyhw/iH2P42Fi2e/E9/2wa5B6rWmPC2JL+mpDXIjtL+JvXhbJfwFzFdfC35gssua1eBDVpRBEroSofSgmOrQBJJXe/lFeqwnsw9HkInj8L6yB9oNJX2EFjv4h75jzUACsDRuGa68K6jI+CEOGeYwNYQWljp1pgUk84NySW4lrgEuwRHdMIxwc5DpNDckbXymZRM3H2J2WttB/ZTr5eWmiF9qNIxnxP0F+MvXx5PR8oMpNzBjZOxovPXgFJFpg4RizGAdpJY2uab+N94U8UYKTnSDPYxve607zTiFKe04pTCIgQ1NIiIWNP0G/LyYupwb0rmnPFrhq3h0XDCvxwBAcAFeLXLaBi0+l/65c/xh7oCFS0BFBBsMBdyh+TUaFLgl8RZQuzm930r8c9jM2Aig0naAc7/DGAivCm2heM/PGBCibAHaOCZtp5mGnr38aqiPf2BECABYe2+Yahqkk/cRL3gAokBayajlXkTj6qHaPCpJ/yeXhULFN6BlWcKbA5nNTU+OSEowCqRrIi9CFQQVoh0jtuA28JEAuOKP8EoKKvj4kH84NgkhCLDBYeBIgIFIDK04xM/QiwoFjywTbgAbsCSQ6fUYFFlIwKABWo6mhIqVjmYp3JqN71yOiYpLoVqLAADqOFbWk0mGQgUFHUhD+eE/7Y4mltp5+G04bGwkxJr3JBGkhmNSJMhiRSScn09pBZoWgKdxdiQAWSovA/mJieZMIJ/dYKVDAoi6MqWIMZ09HUgCQEKvCckWwKgAoO8RCowP+Q7Hv3nXdldGxM9u7bS0YFEirBxsOqapyZtlUQW2BbKhZphIzzriyvydpaVqanZwLjrtdffZWa6zCl3r5zlwZn8NtgJUddioVcIKNigT2DYlfV/TigAvENqk4gn4X3Gs8FjArVViaXWz4/81nAqDCgQoNT57uBwAYBMYAKJNwbDTl9+rSk4kl5+dQpjhG+E6SiKhDHaiqAWeWyXL50CfUzBCHIqHDST9QixzsQiQRABc20HVCB52iJ+VaggvRYiFg16lItV+Sjjz6SEz95QXbC7LwrTaCCDGYmt/TzQwMVDGyDrFtE6lEAA+5aTfN8hOM7ALU6rQ9t1xUNFt3KxAp2jNsENEkaZfn0499ILrciR597lkyUnp5+6esfkQpkuwSAhX4eB1T4wfBmQIWdC/eC9x0Jw9HRUbeZB5jVeXH0EwS2yXjcUqoUbYw5VLNHpFJckbW1e9Lb7YCKak6y+ZVA+imfqymjIrIkAz3dsnPXs1JP9gE+lndf+/9k985Z2TN/UMqNuOQLDfnu7IcSid6RQ/NH5NKFKzIx1SMff/S1HD9xTPr7R+T895dkZmZapqe3Sb2WkXq1W2pRpZu3+7RuKJo24wGjQoGKd95+Q3q7u2Tnzu30NFrOleTKjbuy9OiBrNy9If3dUXnx1Cn5zelP5OrVRenvG5AdO3aoNwklBlPS398nd+/f4/s5MDBERgGkn2DyDjPtklQoh5ROxKS0viaXLnwry0uLsmvntOzee0Ci8V4pV7okm8MYa8ja0h25e+ey3F28wXdzcmqbzM7NSyrdJ41oSlLpbpVbizi5AMjUkWUQSuygbT5QYYkG9AWACmNUAFzGJrpQKPIcYFRgfgJwC0YFPCMwjxCoIAYNtl4IVJj0EyTVciWABgX1ewCYUmkBKgoFWVgEo+KODA8NEBQnoNlQijuACoAKq2urXMuwXpqZtrEXDKig9BPYBjnITxY495mEEzae1TqA+lzAqCCzr6aFBGARAqigSaIDCegf4dZW+k2srsrNGzf5LAcGFKjgpwWoUFaNmkADpGgFKtDflFbKqaE6pJ8wN8OjAmsjgAm0Ibu+zvs1M3CLl7DB9oEKgCH42HE2Z9immHOUgcJNrOjmuc9nVJAdsbIqGRi+O4DFRGaCJGmQxdEkI6QI19baARWKvjMJsQlQYX2G54Y4CcwYP04yoIJVw7EGpcIOzB7dBKgIKx+tD55kXus43W/4RTCLP/60/hG/Pxq/+fV+QKBC327vExSHdWjCnzNQ0ZJMf5JHaoU3PNbkdHSxbt+BHWKQJqA9+K5b7dqAFZsPgfbXbmYQtL87Tfm5j+ePEfzUpKDbXILzR5OJdHgNzj3eJR8HVCD60Ap6mP9aRbgpMGzs2s2ACk7h7pFQGsYZNmtcqHOI9qefzLfcqrYU1dedgAqThaFsi8mrmtdIc/ClDXdjgKa+WlXjpLtapaH08Kb52B3LQjnHZquBeaALtZNlMp9IjcBb728zoMJ+p+CAJuI1wes8DVyxGc7bKebyi+qs/b4PpXmiGFMG+xCwZy1eCQEXM3M2SSLVJDa5IW2rWwPYL8qqsDxBkFAn40XvBedGUQWY9gaCqdwh+kw9JcghdQwJ/M04AjFLuaKV+riOxzahdBQLy5SNgOQ0wRqwVh2bAM+Ho809ewATNQELR/fKuADHOmWVnDk3C88cQ99JLQWghZPewldtT4zvhaxOsB7KEgfDH0AFOoCX0cHOa7bbNERDJQQcinslsMO2KbuEiX4AY/SFUCkwFseBSeLYCwCeWPTnrmUSSOb3YnJLqu7hwB7iFlAf0LHAGhHHDLHJw4MSAuDH3l0r0qDvJUEcZdOEHwXZcA6YYwMEArBlhukbM4wKarT7qME4WLrIEVUVmIpBxhUSrCrHFwCJxrjDPsp5odgYVSKYY4OFCVllwESE8l+FYmELqOgQjmz9+EfcA5sCFXZfTQHT0wIVurlu/nhhyFNLP3E5/YMBFZzI/TDJNVXvoE34FJRZNGd/HguUtBkzj5d+CmNattM0NoNz/QkAFWUHVNCPAibaG4GKRG8/J2ksWKYBGGy8dRfL6maCEeWylEuofiy6KnlF140eiQV/M6ACibqV5WWB9BIYFQAq8IRRkTE+MeFojkDK1ehaNQXDZK7Jwlg1hlXAY3HFPUASA0n5JPQsnc8DFhhSHB0tNRhTqHTnz7Tqh+yKtTUNGp3ZFuUOWN3tzOqMekk9KPSLBhGMHViFAxAgIWNjY9LV003wAG21ah2rjoBsRjqVkkKxyEUdyRF4iYB5gA8WfBxr1acauMGMGxXRRT6HeqXGpAHa2D84IEPDQ1p56ionTPppdnYbGRXTs2qmjdAfiz3MtGEsxWqWBqiP0JDWoJn95UAhVOVqAYU+Z7SpaIwKDcddUI1gXzWsT4NRMTYu+/bvl9mZmSbpJ6tkAZkD481ozxbEglFRgwwKEizol1JZenv6A13zN177NSuejx8/LnPbt9MEGsEUAy1pMHlnVS4WvKtEVRgYq/TTZTIq/uF/gkfFNINoraBwfius4GjovbrqFgveAFQArHnxxIvSPzQQeFQg4FT6stMgF/hvIOEfkXfefodmsa+8fIqGYrxfV8WBChQGyzHIupTk0oWL9FcwoIIBODdc4cx37Woo/QSgIqzQ0fZvBCqcXjDGW7FEKaTnjx2XudltrIBFAEeABgGhow77M9hmOZwmoNrbiVsSTqfEsIJJA22wk1AtFJ7ZzkPZLbcW+ZVX/jTd6ZoKUujmTEetGvQhwZtJpyWfXZZPPv1ApFGS/QfmJdPTpbr2mT6p1nuD1oBRw/ca73gEAS0hsXDf7wJ5LycYNK/ThpJyYJUK50iOtdZlrHUdegKPio1LlwdUoCqquCJLy3dkoLdPctmqVKpZyRaWZff8PpFGrxQKdTn37edSl0cyNNAn27cfFklgPIi88ev/V+b3bCdQUaknpVyNyPlvP5Vy+aYcPnBQ7i3elXRXXD779Fv5ycnnZKB/WK5dX5TpmVkZGBiVRiMj1Woi1M7bkAdyGrIdYjYKT3C3jVWiJm//5tf0fNi9a5f0Dw3L4v1luXbrrqyvrcjyvesy2JeQEy+dlLfe+Uhu3XpAz6AdO3bKFGUFawR2e3p7ZfH+fT7Hwf5+JlOLxYpkIUtUrki5XpN0OiHpaF3u3r4qVy+fl9GxIdm7f7+k6N0BhkRMlh6tyPKje3Lj6ndSLqxIX2+PTEzNyfj4NonEYCCeFIkmJZXukVIVwEJddY3ph5RQQ0UDhutqpo0Ry2Ow5jjTwr6+XrLYsGFNkAmHJL/KC2GuxXwB5ggYFQAqMK5WCVRosqBYqBDIBJsDkkb4fcioKDoJoYyUK3XOT0n4JyWTPPftO7dlkUDFINdVxDg005aIZGCmnUgFQAU2d/fu3nWAcYuZNh1/opRIxPyMtQbMty6TRqyXpVTIK6MC0k9IKtCjIkcJBEo/cfOtskvYZOJYSivEkwQqMN8BoICcFz2RnMlkGCvATBuylABVorK8vMLvgW2i7EJNHAAIANiAdqA/8b4SqIgrMIHxiMIG9CMktUwSCX/jAWJNx+DC9x89AlDRIGPFvLCsytQkBvx5LAzxdea1tnNDzA5Qmci1VQAVGWVg+vJxThOdq7JmQpQVWCwxtgmknxwDwpJteK4GVOC+TPqplVGBn+NnrUBF2AdRicQbjDP2zxx5DFDhV0E+yUrTYQXquDBx4ugws3T6cZudwg8JLvyQ5/JuwUvTdr7fHwyo8KrNn7R3vcfw+0g/tQO7ucpv8pg7/aoVqNBQtvOJNjtPGAW7DkFldlMRT9hRvxNQ0Wnoe4wKH6gI/u0uZv2GmKqdGJZp7Lc+Tu47Wt6hzYAK/I5FEq7yHPsJY1Q0ATpNY7eT9JPrVVUxckC1SzR7Ei+utNuLvUKgwvZNYelN8x1Sxsclbuk/R6ki3e/YWGjX9YFkmCu6suRtu/7Dz1q19XF6Jke9anAzFsZe1ub+TucL5ncP6MY1WKnvgAgzKbbEqsWbxpJoHu6aAMexYQW/7oUs+c/jXeLW4hb0DWSeWNRH+SDdU7PYybER/IJCK9prBfcYWXPvqdK0NDV2bHPIOMLQGgVcFhMZKKH7bhUn0+vant6ZiDuzcpXN1HYZUGF7Oe5RFAkIxi2T8yAlO3+DwKPAFatRDQCJbbdWom2qPodnAMkfBS6490dS3YzTnek03yo+ZpUAhlSw5VFoUE0VCE2g61EoOLCK/c5AheahVAmCiX4D0tgOleGy8WBeH9z/15xPpGOzIx5Q7zTtVwAZ2seWyFdwSY2nQzNpyik5U2zd27RbmfS75klhbVZwwr17Ln5RwA3Fssrg0XGlbC1jYnSSeDJ5qI3vEH6i7wnyKQBzWA8FH1IWNDpQ1TWd70UizrhQizyh/KDMEpsfOae6SZfvi5tX2AVbZtpPGiVsHfdj6YFOQEWA4NuNeDQq/ZEf9OtPLCAKcQ0LX35cQIXenbeBaGvs6jZ2QS2w/8R/F5gCoHVLP3kgTphQs6oJXZibPy3XbQGBLJAN7o2HK5rc+kzdE9UFy6vU4ELkDufC3uJRAYobGRUGVOQLrBb0GRWJ3iEmdnWjqkEeFjMNHJwWIGiFqDYsFqRSKrIqEkagvuakAQOoDKBJsEPs8bctjpjslx894qKDTX66KyP1SIQJgZGxcXffNX7fAh1jTHDhdGZdtoE3EAD3jt8j2TM0NMykgv89q9q35xPQU2Ngbqg+I8ECJCmcl4dVX6LDEXwgOGLy3rQRXSLE3j30j1IT49RBR7V2V3cmCEAs8MIz7MmgIjQpMKaOxuKsElGgIilgsSAws+pRtAPn1iRnmbTQcrHIPkTCANIj6BgkB4bHBpl0xS7p5s3bcvnSZbIRkGSa2w4JKPWoSCaRrEFlqWNQUH4rGmh5YqE1imeEWpl6l2gTTFiRHDPAx6pCLCmNPnz3nXdkbHxS5vfuDzwq+B477Vg+W0fLtmdj70+pVJBaueTYBniuVSZlEJvg32+8+iqTZMeOH5PtO7aTUIZgT0EnrVo3cyy/bQ5qIm233ojJpQvX5d0335X/9R9/LrPbJqjJT01c8z1xgTLAPXh64H3Fq4bg7PNPz0itWJYXX3hBeob6CCJokK/atgiMESjBCJaBViMub735tnQlU3Ly1AnJZND/cfpCKKvCVQJB1qVclksXLtDE/ehRSD9FyDpC4Eqgwk0r8Kh4+OChPHvosPRkujm0rYoEY+XmzZty/vx5Sj8NDQ3pOKSJWkxy2XUyKgBUTE1OsloaiTXzULHKqCddN/1km7UhSLJ12plzb+DPsX6VrQblPKSNRwWesz+7WnttDOpzx3c1mLQqq2QiJd1dPXL37m354rMPJZGoy8GDuySVikh/74Ak09tAwHBzKujyMalHStKQvEQw0Gx9QVV54LURaiO36y/dLHsBewBw6M/8ZWFD0rJDlaP/rDde07xYUBUVkWppRR48uCkjQyOSz1akWF6R9SIYFfskGumTYqFBRkWlfl/GxoZlduYZScRHOH7/5dX/KnvmZ2Xf/BGp1lJSbYh8f/YryWXvyDMHpqVcykkuW5Nvv7kgL7z0jPQPDMvdezkZG5+TZLpP6hFsOLHZMOAIGwLdaNi7phuKtukAcMgIoOE51KoFefvtX8nwUL/s23tQMt0DcuP2otxZuC/F3Jo8eHBVxsYy8vyxF+XNt96XBw/XZGJ8SrbNzcnY6DjnBPgIdWW65c7DRxKPRGUQMoEwKyyUZDmblRJYg424pON1yS3dlssXvpTuTFrmDxyWTN+wNGL9Eo0lZenRHbly6Zw8ur/I80yOT8n49JxkeoclFstICVYUGEixiKQzSfpEAUC2JIABVTZnYD9skk+6zplRYUP6+vqdmXYt8AuA1BE+pQLW95L09PQKpJrIqKD00zLI/ZzTS8WaZLp6CYDk8+uCfRlYJfliUdbBqEimJdWdkUqlTvo+vRdSCSmXi3Lz1i2aaY8MjxDM5Aa2pkUZYJ0kYymyC3Af2MAt3rlNUMGkFK3SnutHIyqFXEFyuSy9QvK5rHRlUpJMwGRRva9wToD4xqZcz66zIADAhI15gPNkgWS6CLTHosqouH79OuewwUHIeTlgIwJNaCclFwVQkeIftBdAxaOlRwQ2rJ2YR7B+FQp6DfzBnLi4uMg24fyYBbJrWZ7DzMDRNpV+akihGEo/QeoNHzsO7cU1LP7w1ydbB/05oN3ch9gLQAnb54AKfw4gO8+xNKx6F2sigAoAUZw7uSE3CQfdnFsxhQEVXOvX14N+wM/RBxh7Jv2kcaL+PAArEkJ5tX3Tz/4JABVPuoI176Gav9XB/+BpTm3H/pBARVhuretI0J6OWe2nanFnXON3AICeEqjohDx0SnZ32uHxsp1uxKuGbyp66NRLHWSWmr/r32gnDmFnhYFOYEhntkP7quEATHD3/zigsfNMrAAAIABJREFUgknbdmswgU/MoW0+XtFM0/xjkjlMGscoH2SJ4Lansarkll8GNYeUGHJG1N7cqf3usyqs6NySziErth0YjMshXqeET8D+0HfdKviD19ZvmxfPGdCLIMeKiJoP1eSnxZ9M1HOPrhI2uL4mbF1i3xVucTZqYfDYnB5OJTparDAK/zYfDFs3sHapQbUeazFG03zB+9GfmCxTqKig37MiP1u7tA3q74HHZzK22nfKpsE1/Sp09DHWHvuwjdZ+JIMBGIFdXqsFUlX4t4aHSBYjp4B+9se8JZU1JgELPhqzRLYCDWbYbdXyCiZo0ZYl2dEWJuMdEIP9G66nDHAtIsNHC0wiUhV4SMJvUscK9vBQZsCH+1hnDk+wAkwD/M4q8En0DAviTDwZ41BZA2oujncGz1NfYR3TYf9vfCPxndD4Wp8P2xfEkuHI5PmcHJc+B/WrsMIG/I5jlpKZyKVoTIH9I1Up3OW1iEiBFMplOUkn9iXGAowG9Q7cfVi7FDiyX5kpOvbCfKuNVeHGE0EMV6xpoJOCVf65/f91nmPJ/YD3ZKXMZvlAiBvW+vwgnxYHmFjVOLCk7H/EPHivAuDLMUv4frqqVfiFBPPTFlARDrytf/159MBmQAVfcZvoHwNU2MJjr2vzmvdDAhXNbIpg2mhBSR4LFbQsyvY0/cDUT+i3D+isWqT1ao+9etvBsxlQ0TwN6kKvleKtH5vRdYL2PxuAimCWtKNaz6fB5FMBFU8g/ZTsGw7Mm23jHDIqNgIVACuw8Y07mQlrrUnYWILfr6qwxENboEIiDExGxydd0SBYGaH0ky3OugHXShR/A+8zLnD+kZGR0MDKM/nmQusCEb96kPTQhrIafHAjn8tJCdUi8Ri1vxFIYeGmjIVVS7RsD62yBpWX8A2AV4V5L9h9wEeiu1sNPFFVioAIFRmoxNTEA2iImsywikb0MdqGxbVYzAvkkVhxml2XSrHER4ANRe9Aj0Dqqae7V27evKVAxcw2JqInp8coiwFjS5V+Ut1vjF0GIDA1RxbLXQv9pT4VZuCFKpKaFGDQ7kzA7fZtXsLYxH28Q6BiQvbtO0hGBbW03ccCA8Y4Loms19LABWOrVi4wcELAA3YJpE0MqHj91V8TqHj++edl29w2AhVMkjiwAobtFkj4c6Zz2RABUCExufT9dTn9m/fkP/7D/yjbtgOoUEkQu39uKOrwvEAVcpzX0bhMgYp6qULppJ7hPgZRNsbDRBRqy1xAVo/JW2/8htImJ0++IF3dClTUCFRAA9UZYUe0cuPC999LLFKnDwcDf5wJwVoQ8DVopg2g4sjhZwOgwqp08bcPVJiZNuePWFSKubx8+MGHcvzYMRkdGWEiDeAaWVOOVdEpKbBhhmuZu+17NiZ+1/PYdkQ3g81XVcgw/Ni85a8b/vWtDRjzfb0DUG6V2zevyGdn3peenqQcPLiHVVxd3VPS04uxhocNubKk1CMVpB9ZaaeogurI6hKnG6VWMKJpnm9JlPjHu1O0XX949qa8R/OqZ3NZ2y/ziwDIolIpLcv9ezdlbGRUcmtlKZSWJV9ek93z+8moKBUb8u03Z6RSuydj4yOybfawJB1Q8atX/4vsO7Bd9uw8JNV6CqNZLn9/TpYeXJX5+XFJJUTWV6vy+effyEsvH5b+gRHJrjdkaHhWao2ENPDesIrTTNPDvgt1ms1ss/VOMFoBVKCXE1Iqrcvb7/yLTIwNy/z8AYlG03Ltxm15+HBFCrlVeXj/mmybG5JjR38ib7xxWlazZZmampapyRmC19iEd3V1k9314NGSxKNxJqlh1pjLF2UJJsGQaMJmubQmV85/IdFGQfYf2C/Do9NSrsXIKHm0tCTXrl6U1ZVHMjw4JNOTszI8NCbJTL80YmAIxqVUBuCB5Epdkl1JKZeKqtftNnJYE/DBGkA/HAdUYA4hs8KbD/v6BpiYxntpxsb4Pz6lAp5nkfMjwBAwCfDd1dVlkYhW9ZXLdenu6uV5YViN+gMAFblCQXKFonSluiSd6Zay0xnGewCWDADwGzdvEqjA3IA1BBtIgKutQIWyKJOycPtmE1ChyWuNEaONqPOoyEoiAUYFjKwBVACEUtlGzEPmFYW+QlIc1wokjhqNQDIKoAE20RGJCySWMN9h3QUoq0wDAHYqF6C+IPDRAFChAD2ACkg/9fX1aTLHyZ9g/QHroysN2S6VkEQfYIPKa0YibBeKF4wpgfszicZCqcD5APcBoAK/M6DCgFMfrLBYphkc1gRcu2SVD1SYp5X/5ti8YIUriF/ACnwSoIIb95gyKnygwqS9DKgAm1DBKQUqDKwgyJHSoon5yUM/MqDC78Wm1WXTSvuOk3e7X/zQQAWuEVTNB6tf+yY95bU7H97Bc2CzbdYfGKjY9Bn4RQLuQL5XnjxSU2K/w8kaTNjrkX5Sv1MS3D//k46RjrFSBwQDMX+7jybN3Me7f7bf/aJlhLcd4+RmBobILQ/YAyr8dlOe1BWImEcFJV06uLxr0tTaqn9rSMmdrjQcMM57ch4AOlc2FwaG19Ckrn40vvYT5H5/qXmxSrCqubL1WrN0jN/9rf4OPoDQWpBic7ut+7ZHYBLYmU0H33djksdahbbX2HbxdGuRGP5v6wiuZQl27Ql4AAAESLNin/tz7ImdDFDY767nvHNhH2bSt3xcUTXm5n7DmXZbgUUoVayyuT7wHRghG2MbjIE6WBSQ8VFWBmIB++h7qkwXxCVgfOuU56rfncQRDlOARKvu8Sf0MhA+YxRqkK3C/aLuc+15meE75Z/gCVipMIYAm98q5y0m04r5MmuWqEJRb5Dhb0CFjXnEdSoP5QoDHNCg41GT7Cx8jEWZBLdxoDJNunfUIgsHUNS0n3SPqu+xfYd/c59uOQ4FFLBnJjhFsELlnAD+MF5JaH8qcONM753/CPqGwJvrS+v/aBzxJKtw2H/oL5wH8YWahodsIL8YMZyKtECJY9SYRk5uyZ4bwRFXPBqysfR9N3CAxaVkgmDv4GR+3T7UAEN75ylDhwDbjRnN1WkbfAZR0EYyUUKFDBTxptPwcVWwiZ6RzqDd1gIzZuc9uCyBzcFbjIonXf22jvvR9MAv/tN/t3lb3cvor+s6EQZTe7BAO9DU/f9xoZgXhLRU/m/EEFyyJlxOmtrcqSrEQo/2N/gEYILfxA69pPXu7kp+wzdrVIdzPTlQsdkj8+9rI/CwsVTFP6aVoWGb7nCB1cVWr48FExMyqjWwKGOxLZYLrNRX48w8k66tHhUAKowNYQGAbUBpzszFK2RUGFARS0A3OmwjJn5b4M28yxZOq7JoB1QgLEOCfmxiSg0z65BGUaYDTYldcKrVIJrQZrLbVQrg5waSYBMP/XcmgECrDQy5Qu1I3KPpgXPBhkGp+Uc47VELVpCQyBXyDMqgx00AB6kRlxRnkbX7+FWS1G+Ox8kaQeLEpBRY4RhF4qJLEsm4AAyBDBP6Dcl/Jh5YmaBV4KgeRXLFjESxQELCC8n4WqWqQAXYDQz2oJ1Zk4mJCZkYn5TFxXty/dp1mZmFDMuAdPcCHEnL5MQkK4v5jF3ABOknBCvWTqvKNKDCoWMEKsjSAVDCDUyYTLFAGs/gnbfflrGJSTl48LBMT00FZtoW7KnepQbVWkWh4A+eDRJu1RISwyJleKJQ+qmP4xyB1Wuv/lq6u5300445cn4CoMIxKizZZ23iWEHiFuOZjIqoXARQ8fZ78g9/9+9k+44picRUNgUfBnCuSgp9jag0BCpEPv/0U2mUq/ICgIqh3gCosI2BjgVw1pWK26hF5U0CFSk5dfIEK4mRQAIbl31APwyAkDEG99+fP0+5teeeO8p7g8sKz+nGG/5tQMXRZ48QqMD3rWIKYwdJxvPffScvvfQSDWb5rmrcL+VCkebex547JiNDQ7wGximSawbiddyAt5nu/GMtUWbv55MCFZy1vTkbLBL72Ya2dDBybN3M+ZtIrX6KSm/fgKTi2NSUaH78ySfvydjokBw+dFAa0YT09vdoYFoFuJZx4BCqaZxpG+N3Jwvl5t7WDepm97wZUNH6PSVx62czMKT5kRigrYyKSmlFHj68JaNDI7K2UpR8aUlKlXXZs1eBikK+Lt9+rUDF+OSIzG17VpIxZVT86rX/KgcP7ZAdcwelVktTZu3G5QuycOu87No1IoP9XbK6VJYzn30tJ08dlv7BEanU0tLbOy5FdFcUnh9497DB1M2V9Z0xKur1cGPafI+YXHQjGIum6Cvy9rv/IjNTEzK/e78UijW5ev2WrGchhfNQlpduyr59M3Lk8HF57bV3pFgWmZ3ZJuPjE9Lb28cNFir2kVBfXlqWWCwhAwMjEk2kJJvLy0o2qx5AhWW5cvFbKeWWZO/8dtm+fZdUalFZWs7JnUUwDBb4LObmdsro6BSlnWKxLokkuiQSh3QftHqrUiUo3qDMG4GKWFhZifUJ7ygS33jfG3WnjRzT9x/j1mj//f2DTIzb2op3FAwCHFPMlzgfQ/rJByqWVyA5pHJ+lXJDujPNQAXkpMCmAKhMZgQqxhyjAgyHLgeugFFx+/Ztgv9g6jGR4BIV7MtYkubhWO+wTvlABe5NAX3dGEbr6t+Qz0GCCIyKdcl0wTNCqxGxtgFwwRqI82EeAZCAE4BpaO+2MSr0/HH2HQABtBOAgJppYy5XGRLN+SD5rm2k8WckKktLywSAsEYbaxHP1YAK+JmY19XCwkLAoMBoRtIf92Rm2owjUPAAoL2sbEO0AQAKfmfH2QYZv7eq09Z50v5v77SfjOAzp/TTGlkmBlS0zj/4Lgs4nPfUkwAVNm8b6ID/W1+jf/As20k/tQIVyXSMHhW7xw92BipaWHLB/O4qe9tH1E8ZxD9lYt6VhuqlOxRObWjX017jaY9v3xGb/rRzHX+wkLj15OluNVyHNjFH7rSN6/DobNxukG7qoOX0NLGE3WSQtnZ69owEnQxMu47sNMoIVARl/i6R5yX2Np6r/ZmsQKftQ+x08Zbtuz3jJsDEZ9X448xjnzIB7syEGYtbcs/J5/jvgCXc1MTWadh7Zr76iLTBTeu2J0Vnc5cyKNsPDvPDY9OcubBPFmr7LS+5oRI0ThbG8iPefSFxafcZwBCPeQ8VjNCq89aCmMfFdjbH+9f1n7VJMpknXeAh4ec3msaB/ccBN23abgCFxcu2j+lUzGKgRVhEp8UHTW1xD8Hf19oTD4ajK1rw9/lcezzPPfsdE+KuwM+KobCe4PeIbQzgsBwE74l+kqFvIuMiJNWdn4iNLx0O2j/qzaCSSQQ2PDmkYF73i4t4M5pAx5qpfaKm2jQ2DLwksH+EdRb8BNE2J4fkADP6PDhmIe4H7VdGZkVlhRzAEChNBECA9qb1k40bFKVBVstiRRwDQIMFeWyrJtqR6wGIg320JspdX7h2254QMZC+supNgX6CdxqzeZ5cF8ErV9Bpx9uaaPkltqkOb0Uz0Vb2FNgH+CiQoMxufMzI3Hwz9H3Vwkd/rLLY1727fM/ce65PVmMaPFsWzDgTcwMqLCdk74L1J54nckGhObeCEBZfM//gFQYZ+8k8Qykb7MatnVv36vrc0OPIIWn7bC+jfcznvsWo+B2imK2v/En3wO8GVPhxdRjRtAcqOt3+nyZQoQwC17YnwDJc6B1WVHCGM6pamxNsErA8LVDRvnmdgQouKRu+9EMDFUUmMJggcJJGrUBFqn8kMMK2imyrltMqFZIIOdFXypAdMkZFkpRHq+AwAMAqDy0wxUJplSRI+q4sLfM7rJ7MZMggwGIyPjntFjgExSonoElcBSuMUWELkm2QDaTA9ZEkR1IFC6kZVVughfYYqGEsDAt8bHH2N+tK+awpsJPLsxoD5804HXAudB41E9+1vmAA5iQRAMJAFx2eHGgjFuOe3m6aZQE4AqBBWSej6UZw3xq0WyLFgl8szrn8uuTW1+kzgHYh6Yz7ANuCgEMsJj09fTShXl1eke07dsrg0KBa7NbrMjQ0IpOTkw4A0b5HEo1VMg4ssOBGqafGqGhIHb4ZRWVUhJsKHbMGRiFI+81bb5FRsf/AIZmZng5MxS0Jw2NdsOlXAKF/AqBCGqTMQo99oH+wCaiA7AcYFdt37uB5rK9xfppxe/IXwTUJYtZV+klicvH8Nceo+PeybfukRJwUFu7FkvVoD94baNySzcBgsyGfffyp1EplAhX9I+pREWh/ujGL8WNVLqj6ffP130gqkZBXXn6JQAWYDag21/GNIEd9FDBuATBEGjV5/vnjDtBQQMfHkK9dvUpGBYEK86hw+rZoPxJ3586dk5MnTzqgwpnrOaDigw8+kGcPPyvjo/ASUHm28fHxJqkkC6BbV41Om07btNrxPlDQ7lytGyn/vJukQ3Tz0UEWqrWtzRvLiKS6MtLT3UV/mWq5KNevXpL333tXdu3cKQcO7ZFIrCrprm5JJ0ekXod5LtaPiv6xCRtrCtkU4Sbdv47NOX4/2L+DTYCrJGyXm7BAuHWT7N9b5w1zq/TTsjx8eJvST2srBckXAVTkZH7fAWk0eqRUFAIVxfICfWxmZw5JPDrM+f5Xr/6zHDqym0BFuZKQSCwuCzeuyvUrX8vMTK9MTQxKbq0uH3zwuZx85bCMTcxIQzISjfZKpR6XRgQBPAAK67tmNoqOl+aq0DDpoYwKBTigjb8sp99/TeZmpmTXzr1y7/6yXL+1IIVcRVZXHkh29Y48d2xejhw+Jr/85RsSi3fL9PQs2RQAZtHd8DDA/LuytCSxRFr6BmBqnpBsPk8D6kq1IJfPfypLDxZk545Z2bd/n5RLdbl3f0Vu3rwjK6sPCDLv2bNfhkemRaJpKdcAnCcllkhJFPM+WGWFojPx1E0zJRiS2ADr/GxyDEg066Y9ElDLTbbONkeYywFIY36nrGIiwQQyN+KlKqUdAVRQ+imV5jy8srJEwB+eDJB+6unuYzJgPb8mWLZ6+3okR6CiJJlMjyRSKbL4IP0EoAIeHQBXAHYu3FmQsZEx6R/o57Os0CgySjk+SKlhjcJ10d67i3cIwOM+cW+aiHA0eiTxS0XJrq5KIhmTggMqKHkAP6lKlTGBARUYBwAqjFFhG0/MxziGXhYxABoRuXfvHuWZwI4AUKGsCfB43EY8AmkiZVQAqEK7Hjx4yH6kF0UKMm/6Jqr84zp/5gMV6HcaeEeiBCpwv2xDQgF/3fhGpFhWiQBlVDzkz1SmCtWauq7780OQrPWSbJ3mVwMqAFTh2rhPH8iwJI9dg0nAGPo6L7ncuiTBovSkn7iZdvOoASc2PnEO36PCkjDoM0gHoj9YsOGKNigdCTZGCqD3oPyX/0eBm63PVg907IGnxJ62evLPrwcCIMkDWiwx+aRb/uZU/gaCRkunbQ26P79RtHVH/9o98L/8Xw6QcnLJACmYT2FOSA3Oa7WKGnPbx+2XFBDS2AXxKj05nI+IgZQaFxlzhrs9FmNqPlC97dTnMWRUaCyEPYVKzVpxKy7PHJRjhylwqo2ymAkFkRrj6N4ORtjYV2thlQJZPN4VV5KZYaAKFSnUK7MBKWd6fKoR+hZQ8a89Mreu9wfvgS2gormLA21NP6P/RNGLTmb6cf9uV9HxRwQqiMX+qwEVBckj4d6GUdE1ONYke2STulYIAqiggqGCBfBSKOQD6SdUJxqtFb83TUxsotnzDhww0AHXR5IIi5IBFZGoSghMTM0oUCGgxcIvQVF5Ayt8RoVt5C05bpXsSPI+KVBBcyZqK8ZoHoxFBdeyikImkJ0vACoWYGi6vLwsiYiaaLICxIyX3EizvsDvUjDoZJWKoveghw7095NdAHYDEjrruVxAP0T1BM8JiiYS4y5RgCpTVN+jL7Cgr6+vyXo2S38KJFXKeRi1ooq3LNWGVjlgzKOSA1rSO3buYrIOpwUIgOp9JHTSaSR64vRfGJsYlcGBvqCSAtdWKq4qaOqrA5PomuQLYOmEjAomPjwTNyTE3nrzTRkdm5ADBw/JDKSf0ipJ4oNMmwEVFep8N1gRk88Xpb8PJuAwe67Ia6++yiTNT37yvGzftTMwSmd7nXSUJfsMBOF1UVEC8CBaxVOXyxduyLtvnZZ//J//vcxumxQhUBFKP1kQg6pjxDdV0EcNqPhEPSpOvPCC9I8OaOUqAiGnzapAB4AKZ+4mSXn9tTcJVPz0p6ckDdNz+nSY2ZoyKqKROJOc3507y0Q6wBgkwnBtSlG5wA3HXoP00/0H8tyRowGjwpK8AVBx9qycPHVKgQrSg0NGBYAKyEaNj41x9KLteCcBViD5aBXCfNds5+jGufVTEH8+YaVoawKuU8UX+36zqtYWoKJz0r6FfSZCBhMqyumPjn6tluXa5Svy1ltvyMFndsn+QzvYVz09YxKPAiBDtVJFGhHHCmDjlNHlCo+C98b6o7UKzb9vv63cMrtErgFq+JH1C+TdOn1a7zn8vwdUIFgvrcqjh7cpU0SgorRMRsX8voMiDSS4G3L2qzNSKC3Ith2zMj11UOLRIfoG/PLX/yzPPjevQEUZ811MHt69Ixe+OyOTk12yfdu45LMNee+9M/LSy4dkanpOJNojtXpaqvUEAUGtSgtBHnhU6HBxFUltPCp0HGO0AyBSRtLKygP55NO3ZW52WmZndsj1G4uyeP+hlEs1WVt5KLn1u3L8+f1y5NAx+dUv35CuniEZH5skEwCST+hfMMpw7tW1ZYnF09LbP0rPibXssuTWluTm9Yty+8ZX0t+XkRdfOinZ9bxcuwpD6SUBQW9u5zbZvXuPJJLdUqnCgyIthZIa8sWh/0/GH2QE87K2CkmqAudXAAXJrh7OZz5QQQZTBXMFvCTgNQQfnoquQUhsx6LS3d0bMCo0AR8lEwLzbrlYCRgVBlTgPglUNCpqil2oSG/PANcHABXxeER6e3skm8ux7VhfkqkuSj9BFpCMCgAV5ZJcv3GDskdgKYKVh+0fAA2smwQVEmkyKpTBEJN7dzsDFWBlFgt5WV9bI0hfzOekuzulxpm1OvvB2A3GqCBzxEk/2Vpvvglqug3d6qjcvXuX7cSzRjs1gY/X1OIXlX7C5ljBioTcv/+gCaiwtR9r6vo6PCAUqEC/4dz4Du8TjIpsls8RTAlf/ghjFRteDG/IRcIDAysojsOzBKMPG2x/3rM52+YIfx6wGMrfUKMYA/2Cc5rXiRZAaLxkxxKscEAFmJuIX5o8KiixEGti6eE7YZFKY1OgolX6Cf8nWJGMbAEVf/Cd4p/JBbZyxn8mD/KHvw0fwGg9e+vvnhyo2BpwP/yT2jrjX2IP/MP/oXkGxBjMEjhWi/peqrck2LL0YITJNlQyWIhnptTYL2t85sc3zSyt0HfG4iLEKOZ9AmlOek3wE/q66d4BUmfOnNspZ5CF4Uzf9SuhdD2lxSoVMk0QV9FXDrkh7NNrWjCrLHBliLhL8i8tjNScFdki9N9UuaotoOIv8e34M7/nLaCi+QE3U1u9rL5LnG6gJAQRjA9S4JytMkqPH0h/aEbFvx5QUXKMihyTzK1m2j3Dk6x0bGIZOAojgApN8upEXasAqAg9KrD4YLGxhSYAKtLpoFLPEgD424AKLFw0085kxAcqlPqHpG+oR9jKqLBKU1vg8HszAUOSAUkV1ZdUCQb8MQDBP1dQyQ/R7sCsuqIyQqQWVgOgojvTzUUITIb7d+9RTxvJ/q6e7iBB4FdJMhkFA25HGbTfoV0joyMyNDpEfW4YkRqIA0YFGQ0RyGUoMIGkDBJCWDhxv6AWrueyrGhcW11lFS6YFahshARIGVrf5YpKNJUqNN3esWs3ZX1gbAV5DSzySNigIhbyJ1hQk+m47Ni5Q3p7e9X8zuk5wsgU0JFJgKH/wIqhj4Sr3kdCzRIqBlYBqIA5OqSf4JnhA1cGWGA5NxDKwCFcFwFCuZBjQFCiwXlF+nr7A6Di9ddeY4Xq8ePHZefuXaxewMF8bp70k73hAUDSAlTcuHpH3vj1m/K//ce/ldm5cRFKP+m9oMLXkj5KGxUpoerDyUH99sxnZFS8+MIJ6RsZIIXWWC8WuIRABYCwuLzx+luSjCfkr352SlJplQajhqhjVHCsorK6XJZvv/mGQMULL7ygWqIuuWVABa5x9coVuXf3nhx/7pj0ditbx8Y03odbt27J2bNn5dSpU4GZtgEVpXxBPvzwQ7IxxhyjQsdXjYk+S0LZc20FGDpV/LabVf2Eeuv3NgUYNgEqzEx7s+9bW5qSgqisScakr7dP4qicgfYuDeeiBIdOn/6lHDm2X+b37ZJGPSk93ZMSj3d5bBYrw9H1xICK1nY8KVBBfV831/kU6KAi2gMqOgMTrb2+EahYenRbhgaGZHU5T4+KUhWMCgUqCoW6fPPlp2RU7Nw9J1OTByUmg5xrfvkv/1mOPr9f5mb2S6UGGaeo5NaW5Zsv35Ohwajs2jWjjIr3z8jLPzsaABVgX3QCKgDyNAMV7RkV1OltlB1QEZN7927Jt+fOkFExNDgm164vyPLaOhkDj+7fkXo9KydOPCMH9x+m9NPg0ATZY2AbqHdDVBKJFAG/1fyaRAFU9A1TWmB99aHcvPqdXDj3hSRiOfnpT1+RYqUqn3/xjTx4uC4D/WMyv+cZGZ2dk57+QSmXG5RUwvsE4+VYPCLpZFLqtYqsrz+S5aX7lEscHoQ81rBEE92ykqs688xoIDWE9QBzNYEKJ/lkbDAC6JQJDIEKS4rjWMx3Jv0EM22AxwDB8Y4tLz+SulQliQ1XsSo93f0BowL1B719vbK6lpUi/X96Jd0FA/AqgQowHDLpBNeTGzduCGSPDKhAeFWhFEidifKuZIZrFK6LufPu4kIHRgUiMLDTwE7EmidSLualF8xCmmg22A+ICcwPAeNdGRVRyhwZUKEMDseoiMPwEkDFPVlYAFDRx/mLHiCQ3QNO5li1ADUCoCKekPsPmoEKt9XlfWezax2BCgQ2YFTgGq1ABcZYoVgOZB8gI47xAAAgAElEQVSaPCriWFtQ8BECFT6w4K9X7UALW5M3Ayr8uc6ACvQfmJs+UMF7dRKavpwgruEDaT6jAv3fJP0UxxqmsZKt3/guPCrAqPjn/9urpHx8uL11xF9iD2zljf8Sn/rvfc+PAzF0Lg8dJ1qzCr93A7ZOsNUDf+E98A//p0o2VyB5xdgAyX2ABmDna14BsQ7jNsdkwJ7X97VUM3kUMqnMV5NauzN511hIFwozL+ce3fm8qCfFRnk0/Z76bJqRu5qVGwtefWWtwMOkMvF7FLqY0T3OUYNGszFPnXy3+chowZqCNWwj8xEqA8WCmS3pp7/wN+XP8Pa3gIqWkMIqdV1+KDDE9SavJrDCD3y9WU/lJ9pQMVo0KP2r/zkAFfQTMOmnAhgVACrwd05yjmHROzrFxLPpRlrVuybZHfXOY1QEHhVJSCiEjApNMpe4gTfzZJvEqVFYrwVABSqFIYeEBAncPUNGBRL1uvCRXeHMhpE8x8JBBgQrE8PqfMomodxV9PpjY2NMZJgPBZkITgrIKt7td7hXJGdYnVpGEr8SeF8oul4HfE4KIBJH/H61Ru3phw8fSiKVZHLFpDwCpkckqjqZkNRB0sTT28e9Do4MyOjYCBdQ0+YE+MEKR3opKP3QpClYSUvdxzoTY7lsTpaXlrTNBU1a8VmDVUFfj4YUIO2RA1ABRsWgxCG3USjwd6lk2ulmwx+jJKVqUUZHRyh/45u84d4xBugT7wAftBOAF3VInf64mn4pCwTP4K033pCR8Qk5cOCQbNu2jdeyRAuSbxwPNC+FpJFWVah0Bsy0CwQqEL8USyUCK/CoQKoLFcnNQMVOSpEYUIFxg7EMQMYqPHSsqEcFEId6FOMoKjevL8rrv3pN/vd//HuZnZukVn3EA61ovBYYi8eoPQ4gCPf4xWef0Uz7pRMvSu9QP5kuaIPpXQambhGnfykJB1TE5a9+9ookU6jARsW5VmPgmSjQIFIpV+Wbr7+i9NOJEycco0L7Secknccg/XRv8a4cO6ZABYM9N17BzoGZ+jkPqED7+H3IY+UL8sGHH8qzhw7JxJjKPZkh+KdnPqWkFZKT1DN1fjCbLbebARd+8uxxgEdTMt7zv2m9Nim3DoR8XBhgQTKOwxIAwA7vczqZZnU0zBrjkImpVuSLL96Xr77+RJ4/cYSyQRFJS3f3EKV9NMQNgQoFQZUW3PrxgYpNQR0PqCAjB347AMNqCPLBYQ4FsAx0tWs1XbdpHWv2qKiWVmR5aUEGBwZlZbkghdKSlKt5md97UBrSI4V8Tb7+8mMple7K7r07ZGJiv0QdUPGrX/1nOfb8ftk2u19qDZhpx6SUy8qXn5+Wvt6azO/ZJrm1qnzw4Rl55WfPyeQ0pNi6pVyGjnCcxzeaGBW2Dod96Us/BUwK92zrjomBqvnbt67K1WtnZXZmStLJHrl5a1FWspBsysvN61dkeDAmJ08dkf3zh+TNN9+X4bEZJq3TqS4CFEikJ5IpKVUqki0XyaSgsXqjJvduXZavPntPItV1ee74frJu3vsQ4E1UZqZ2y9zcfslk+iXRNyTxNO6vRrYa2AnFUlai0RoT74X1NYlFGtLT2yWjw0PSlc5IpVSX1VxVinXIPOl8YJ4IqNrHJgivLeZyvGu2BhnIDWkmJOfxc/MKAOsK70AhX+S8Dw8OAhXpNIfH0tJDaTSq9McoFivS291Hvx+A3ApU9MnKapZAMIGKTIaMChiMA6gIPCpu3qSEHOaC/oEB1eF1Bo0A73F/mswGkBCTxTu3ObcBdAB4QeknJsUVqMjlslLM5yUaBdBTkL6+HknAq6dSZz/40k94h5RRAaCiyzGY1GAbrAgFCRKc1xcX7xJQGRgclEEHtLIjogpiqzQTPCpUOguSUQZU4Dz4uW1E8RwMqEAc4Ztp4/+4n9XVNYJAxmow2UTcZdEBFTgn4gQ8U5ppA6iIqIeYzYn+O8332avWU8ksBQFsPsE6hmePPgiu7TbKVvBg62zAqECBRQ7eIMqo4PPQhVsNUt3H2uRLP1EuKqnMEgMjfOknsFSsqMRkE+KpKM20d47u/+N6VHRYGDqR/yiMGOw3noi2HR7/uEXo9/n9E7IVg0t0aLqtF8Gvg0rWzqy9ds1+kuKADd/rAEgEbWr9/dN6VHjG2P61LSnFYikXX25m7Mzvtu1vVwTCeDg04rb9Tbt++v/Ze9Muua7rSvDEnBmR85yJzAQyMQ8cRA0kCIKU7HJVrdXfu7uqJUuusleX/0n5J3Qvd1V3ly1pVbddZVGkRFIWJXGeRxAgiXnIETlnxjz02vvc896NyHgJgKIl0Y3g4gIQw3v33XffveeeffbeXrRw13c/6lZb1bJ/j9lFEV5dQVWyu56ge02+xNMb0MO0CG0GP1CvBsw7lEtx/kScK7zG2phyTWJca/OXNkE16fd6McHnjG7Na4BzcvtB2PZQOp/qRzq8NcnpX58/fpv+7h+xpbE85B7xJseEZ/bN5KtTE/CNvP3qcTMrtnUnYHM7T8agOdYWr//00pwkjff3wOjb5XZNFqe1s3SvoYbTLDS0cziFAN076a/wd5o42x7NXadp+XNtQgGQx6q3ogIrZrNCO+xLtPpe9xV4BRX5nH/t3unJ+b2kSkBjr4wXz2Om0K463p5vLWDCPswx1L31jefC2muV7q7/pKF7cBQKGjMea7cm3UN/Ba2HU1a6FpmGLAK8pXs+oWw1YhLEDVjz9etY81UaSSWMkORXM2qTFNIiM63YZ+zvPHXwHaotYL+I+8Z+iDFvYQWaOuD1OaMHCu+n9gUT9SyGUaa29TvlllCYkEyS1YrfoCgPbbR/83l2HjC45h/9dVh88N3/VeeE0GMyqWxSJ4OssWxZ+wB7Y+ZvhPKioeKBjgOLb/y9kl6DXgeuAf9WL5MUxy1zOAEjohWoMCaGqE8big2dn5A9dwZ6aFGqFmeywMUVUNrnuO+6N1YZU5qJw5CdJt06b3JMOgNuk3SnvBXi3/tARdu5+v6bX+EeUKDCf+haLsatHkFg4Ob2MCcfhgz+YhPIHwXHbu0kLxyINNNurWNoz1LYHY+Ex44O/9t/EgQS3se2SLftpyagwq7R6da1GReWYG03ZHZ5SDT1y+72tr8C/93Wb/zTSz/dDVDRNTTO5LIBFVgsLHHsm2kzSV+r0qMCCe8YpRA6QlNILCQl1dHOZLOiy5LTMcSS2RACFUiwQ1YECf4sNACpHx2XyWmVXKkjMe4ABFa2M3GHxEaZSUYDKVTzWY24sGghCYBq/FagwqqTcUzKIznzbTuOgQwGePgIu3k1mBkmrgdBA2STbt9elqX5OS5WMBalvAgXVV2Yk0ldvHxQJUxENKSrKyeDg4NMYvgLNRP4WAgTicDMUmUV1JgUfb+zvSWrt1fUOB0ARzyu7IMyGBUKVhQKJVZRzs4eZAInnUlJqaLXb9WgpieJ3+C+gSWCa7UxgLblch30U2DStFGnfEepWNCKBvpaKKhiclWlYkVeAFAxPConTz0o0/v3S2e2U0MObPS42YtLnBqWYXWpMVkArJUKWyKNqpQqJQY42c4cwgEmCAFUYOw88sgjcujwIR1nAaPCAR1OJ9yea2UFaeIHAkoIL65evirPPfOs/OC735XZg7MiMGx1sju4x8jIGfiWTiQIiBTRf/WavPP2O1IvV+TM6dPS04/qcwdqYD7mBkWlmuALkkAfxRPy/PPPS2c6I0+efVIlRJCYJlOpzCBWA3aY6dbk/ffelVijSiNsSMfAWBpJca0ewXwWkytXLsnS4qI88vDD0t2Vc1UpdZp+A9C5ef2GnD93ThkV/QNa5YErx3NQLMmrr7wqD5w8pdJP9DlWHc4XXnhB/viP/limJielhn5wSfAAaGphOlg4aX1tgaCNIciqBTNxi4nqXks1A26XVOMGwTtOa9LeP37rMZsZFRgrkK3JSq4zK3FSTML2FQtlef211+Xm/Ofy4NcmZXS0WzKJfsl1TEodiY5gc4P5TDXpY7wvSve1l7WvXVLH2F3B5paJVEDp2ITo//A04aYTD4lL2rQeS7eHbV7Y7KNN9FWpSL20JttrC9LXNyjLmwUpFZY5Z8wefkAaiS4ypD5+/3UpFW/L8eNHZGDkkDSkj3P0z5/+W/n6I8dk6sBxqdQz9OuoVary1hu/kq5cTY4dmZDiFsbSa/Lo2a/J2P5TUqp2SbyegoYRW9hIpaRaK4car4Hmq25AwUIIpOUcaBmMJZrTxZlovvT5J3L9xgWZnNwnqUROrl29KYVyRZZWt+XSxXOyfyIjTz3xiBw69JD86qUPZGh0gusL5upUEmbA2OAkKXe0WcIcmJSerg4p7azLh2+/KivzV+XIoWkZnx6Sl155VWqNDpmaPCbj+45KKgUwMiHpbJdkOpG8LkkhvyGNepEm37VqUTozacllOwkCgIVTr8E8GvOtyHa+LMlMLmBUGDOis1PNFtEPmIMJOLv53ICKXFeO5smYU7DeIsmOxDPGD9ZTABAA/QGcgAqPcWhm2vCowHoBIAOyedvbO3rdPX00D8caAb8KSFehDTgn1oFkOiO1SlluXLkut27elMGRYekd6KXUYa2imzqw5AACUfqpIyPxRlxuL89JB8zD3Xpi1fYaTzSkCAmizQ1J0QS7ItkeGJFrAYBJz5H5kExzE7y2Bj8L9YbAU4FN+uam+jMAvKCxYiIEKiBxhzUsBB50bdL1WEEYBSqSBCqQ8Mf3rVjAYgQAFbg3WAtxLQBrKOcIBkytxnUZx0E7TH5JAV0AFSUOX7SBxQzO24LsA043mvTcK+Frm3QDKpjrcAkI3E+0G2uzeVRokiNM7tjx8WfAgsjng+/jeWJ7vUSO+TLh+xg3kLsjWyYFoEKNy5PJNN/b2VJGiXqQaNGIARVgZ8JMe2bo2O8ZqLjDnmLX1IlEbFOW8847yTtlX+98hDt/417PEbHJ+rKAiqgGazOj16S2S5UV8DTt26Iz2pHPTARQgXNaUt0KYZiYJSCIT11G12uct4prZYNLTFqSz4AK/sQznm29Pk1J3tsL+Ulrlf/LQIfdjmjNAngQpPMsraf3gSk017+WaKfsiXfJ/Kv1nYstNbEfRDJaqERZOQUSuEdz8W67q2PRjetbJukZM90JqEDco3MiAV1EQ0ZXbXOS4BJang0t+HFyfy7WxFdafbD8+TS8Un8QNI/BqHjTbxrjXcbmaiyMP0vlijN21j0KC2PYv/rv4Jl0hZesTQmACT+eDDM4wTkdYGDxua0BZoxMZnzE84h2QgaH0s1M0taZsGYy2wBbL+4nCO6S5HYeK2CyQivsAzWeg2SyGpgjHmHC3gHaWiiHPZGy83AqAzyQ8OaLYJjzA3ASQljjDfCxCvwY9mRuP8+1CKbJxVJQLMZzuiQ0jo01j2uvuz8c08770mqisE/TJLrzMxBNdLNZHP5IzON/lYFl3OCS9YgNsPkqlot8rxMxCwogGc9xJmI/4KV5BT0uixXpDanQAl7sCyTCsVdHdT8ABLbX+Zo2hOxQxCYGlsLcW1kJ2G9q3KPG7Vq4pGbSuq/Q5wySwlUWaikDoM4+NgYEfTvd6dj38Zj8zf8ejvj/8d/BMFyNsyEnrQULOu4h48nYD/eI/RljzIV9KQpWMUGg7+x5xVFtfjbAMsz9qXw2XlTccMwK/In4B3GtPlM+uKbfV/UI9UzjNTuwgX1MKSeNDRXwQQFRivdG26OyVXUUErkxw/tVqfCeAISA7JTGWAA4FAjDfk3Nwl2R732gwp8m7//9n0MP/NV/+JMwugnWqehkNzaOwatpbW0NkZiJciGNzj7N6KX7N7/j/xZZD/td82dBjNAwnTdiluE5mo6zV8I+4s65ypVdn+4hCdK+bMOiujZ94l+adyINtEIg5t4CzqhrbT6KBhFtkZXQQNyr4kXoif+1W3QS1KSlq1gJ2Ad1StFg8kXiHhtnNdOG9FPeMSryyqgo5CU3OLbLo8KACi1egI+DMxg2oKJYkEQ6wwpOBjquwqZagmkogIpOqbHbgaRXtSfrwg1+FFAxtX9WYokYk7IIGLAQ4LcMYJGQx2INNgUTv7ooop1YWMrlkqD6Fn8CqEACwaSfsJDYooRj+FUIrB5wskqtQIX/bxzPAjMcD4kT+FWkE9BOX6eZZ7aziwmheBzBCNB5JDajgAqtqsRxoasNySUmV1BNgeDCARVIRFkVqCZ9YrynkKACUIEFvOoSXFiU86UyK2v5950CE1Ozs4ekr79PMp1pBkUmz4VEhwUl+I2vTa3BpWpwj4yOSH9/r1ZVBUBVngGHbWIsjMZYBFDx/HPPEag49cBDIVBhWvwu6GQy1TMWDRgVpYKUizsEKsqVkpMZAVCRkkqpJj/72c8C6aeDkH5yvg0IvNAeJF4RwFqSWwMcrcLh447qDAAVV67Iz55+Rv7se38qB2YOSCMNU1QNipCMxZ/4N1lCCHjBFqlWCFS89eab0qjU5PHTp6V/YCDwN0HMpywJrWxRjxc13QJQkU13yJNPPqkVqgiE4ClS07GL8ZZMpKVQqMp777wt8VhNnjhzVhLYTDDYdIEnJ6eYXLl8kdrsX3/ka9JD6Sc9J7yf6VFx/TrNtM8+7qSfUFmDNkFDH0DFqwpUgFGhj6dWHT733PPy6De/KadOnqK2kYEw4ZzTPCO3zmLNmy/Ebf/0QIWd06qF/Bbu2mTGdRNBlhQqDC07wE17TDY38vLGmy/J2sYVeejhGRkcGJF0ok8y2X4ybiiGBp8FIEKc2XRT3QpUcKy1qcLzQUnFSZTyrFCacOPAgB/VXyxh1Ku5W6CCo4PgCdgMZQUqVuelt39QljfgL7MilUJRDh59WOrxrJRKBfnw3Vclv70ox44eltF9x6Ue75N6tSLP/eRv5dFvnpTx6aMEKmBqjYfnrTd+LYn4phw9MkH7iddeVqBicN9xKdd6pFYCRUCZXoKkd0M1XHVjYo+i26g3dB5xV9m0hOu6ogDjhfPvy9LSVdm3b5/E6xm5evWGFCpVuT6/ItevfyZH93fJ2TNfk9nZB+U3r34so+P7pDOLZC58EBSooFxSqSz5Cp7thnSkRS5d+FCuXjwnEyO9cuzIQXnvwidSqcZkZua4dHT2SyLZLfFkl5TKdenoTElHBn5Fm7KzsyGNallSqZj09/UycYzxUasrQJHPo7pMPYB28iVJEtR3m3S35pgHAu6tMSmMWRECFVnZ3NgiUAFAHNeCeR0vsCPL1TLXHcj7ZDo72F9ra6uUPcLmEcmB3p5ezglb21vc0CtQsUmGJfwqUOVmiTis32BDYC2/fuWazM/NyeDosPT09TQBFVgbOtKdlC9UpkFcbi/eUqACxt8p7W9NtscklmhICWzOrU3JABhpVCXX3SVxePBUKpxnlJ2YdibZdVlbg6dGkgkPq1g1I2kACQS3k4mQUdHXR+BBK+PwE40RLJ7BRtQHKsBU8YEK9B3aDh8ogiHOowJsDQMc0I9M4KfTjpWoEo8WH4BRgdcuoIJM0BCoaPdM27zlz2fWfgNcERO0AyqswALHsDnbwCeCC2BUOGkwK/Lw9wC2mTdAB2sSQCgAFRh3mmxK8drz21uRQEWqI0FGxczwMXrC4H6StQo50XhSx0KwZ9ArDtoRlex2QLo/r99TTB6d+/aj/uaF7bf5172CC1Hnaq42C7+15/HbX2xkkj+yI60yV7cpoV+gFaaEifCgYe32ZrHm6nv7riXJ2116VILV3y/5pIvI28skfPtPNT5zlf8eABBZyxfBXog6d/tEu8ae2qEtHY8El/t01041+gLbg0N7ATd7ACjo06C/1I82GlCNHINWac7eDWKXpvsQtE9jbKbvfVBlr2dvD2aDX5TiHyKq+6K+31oYY3O13dO2j0xEfxgoYb1hoFFzxNgyDWEfiMQxC8RURoZJbM+LyNYbP16w67G9FMAIAxDtmmyd99/nmkGUpH3HaxGVpZDcc+M8kdrNK/QGIIsd7AFI4GR4YBShGUsR6w0TzW6viXgXIBWq8iGRiySx7TlQ9AXAQIEQxzx0xzdGhlbGg5EMj0stfkTMhL5QdgO8sABYJMgcwAv7ABRzGkDgnky3L9WdDX4fAAQslqjy+DyWY0zgWsjKqFT5p+UbFAxRtjohIBfLKqijbAQcB4luZT6oh1kgUcTktzIoVJVC24TjkP1BMABAAQycFbQM9kDcAIexgPpxakGKjROfzcKvo4jInkWs0ZRGUmUIjNcf/nWYE/s3f64JfYJbrsgFAAUKSyBJzT8B1Dkwx+4fx6FjoKD9lo/AdSujQ3MguE4W0Ljj81yKvnqFtDFVVHD7I8VH9TlRsED7g+d0xRwKiNloRmxoMRnOp0UzuG7cyw4ocziWCd43DwrcrxAIDDZo4fxt6Va09T5Q8dtEUvd/+4fYA3/1l3+yu1l7VPLTcLR11QwWm5aEebAJuAegIkiU7E6oNwMVTeFnm6712Rd3ucXYC6i4542AO2dwak326atN0Ih3zTDnC1TGhB0QDdC0D6D1+1q14/cp6201278LqDDZGK3UY5V9AFTAT0ClepqBCkg/5QlUZAdGuZD71e22sU8kHE0zpj4PPqMikVGgouoqQpFoQ9KcFZC5nNhywOoBzcBzk9seqEjI9AHIDsWlSvQ6zqpLVme0ABW28FgiR8GHMpO9+BNVlUiiGCBhQIXPqPCTqUhA4FgEPBDAuEDYQA18hupNo77it/gNgIrerhwT2Z9e+JQB0ODQcFA1sRdQEVb96EKPZAlkSsiuYNW7VhwgKYFzhVWbkKgqUcZhdWVVK0IciwVB2U4BwFSRAcL21o5sbm7JwYOHpK+vXzpyGQYACAwQLJqcgwI9Ws1rBsomQ4UR2NXdJeMT46zap/TU9rYUiwAqQuknHan6jKMqHUn5oaFheeDBrwVAhcpIIWGl1TE+UGHjDX2BYxfBqJCaVHlflbESAhXPsv2PPvYYfTVY9OaMQSkXVSgow8a9LHizPb8+RQ25fu2aPPsPT8u/+/4PZGp6SupJrTLlxgDjwFF9STdFgIpqYlT41Kqsuoe/weOPPSYDQ0OuUqROMANxNBKSmv9W6jzaB/Amm+mQp558in2PBGZdagRjanXV9gSjolCoyLvvvC2JWJ1ARTKdVkYFKKgumU6g4tJFmZufk298/RHp7erm7xn4uoAXQAU9Kh4/I4MDg/ps6UWR+fTKyy/LA6ec9JOGv7w3z/38OUpCHT92XHp7uqVSqqjupvVnK7uh/VZZR0TLHO4nxu60/u7FqLDA1I4RVK+0SZQ0gQWcVus0Ge7t7mHg2ZzwaCC/Lhvr6/LWW7+RncKcPPy1E9Lf2yeJBEyZu5msQ2wMXwEd81pJ1voKNt5tNtb2GfoVYxGbEGyWWJHT0IBYPU5CqnXrhrCdkiHXDm44MN3GpR6rSKO0Jlsrc9I7oEBFubgm5XxBDh9/RKrSIZVyST589xXZ3pyXw4cPyvj0SWnEHKPiJ38jjz/2kIzuOyTVBqrak5KQuLz7zktSLi3LkcPjkkl0yKsvvybfPP2gDIwfk2IlK7euzUl5Z4sgnqTSrMbHg4qNFv43eTqtrgKY13CGzKEhMO8xgQqdNz54/03Z3FyQiX3jUi8n5erV67JdKMnFq3Oyujovx2d75Mkzj8jU9HF57c0LMj45LRmwKVKOTeEBFYViVeKNiiwtXpeL59+Xvp60HDsyK6vrq7Jd7ZCxsSnp7h2S7a2ixOBdk8hIvlCUpBSlUQMAE5dMKqOeCs7gulyrS7mKDSTo4TUpVcA4S9GDCcAC1krb0MF3BvfbJApxfTZnGS3eByo21pVRAb8NJI4hPYQXig2wZoHFYUAFxgnWJurvJlDRV6YfEd4nUJFMSndvr2xsb5GZAWZfZ0dnsLkmMN6RkWqxLNeuXKW83ODYsPT09pCtBUYFXvSoyGRl03lGAKhYnr/O/sA6rDJVLjHNeb9Bf6sCgApqGFcl19MlcVSmQXah6sy0U5CMwjNWl/X1TSYYLMGO8/pABcH7JPxLlujJgzU0AP2dHGErUEFAPpGU2ysrAaPCWJWIcdD/kDyCLBeYIug/M9MGeIHPzbvBwH5jFOBcBlTgmPCowPnwO2UeWqwWPV/48wjXNbfRNoAzilFhQAWrRl3VpFYRJigdhjajHfSmcMf1z2XzJGOvFKprAWwZUJFz7IkEj1PY2WZM4gM0ZqZt0k9fNlDB+cALp8N5+y5QiLv4SmSW7k4LVbvP73l/EnGSLxGoiLqMaFAgWF35l2D9aSikHnSpf61ti8gsJesVLLi/ct1uaRg/su3ZrvvmkqQt7+8FVLS9PYgCmgoowm/5ScumZ3GvRHSbk7QHhqKBCshyhmCQd8CwVqFNjBEh2xXRIdq37TvP2w1rcUCQt25/sCjgC8Ue9tJ4z+nPG2hhIydMIISjyetjl2fdfc06GNsO50igIur7d3pOveeP86OL8+4VqGguCtW2c55udyAmV5WVHQImWrzH5LiTyvEZDVq0Fyalg99RjibU1w+eaFcqb+2yuT+KxMJkuPPtQ5KeBW70cIweG5SWQqGCfReJYsoXO4laJ4vcJAdFlkSFLHSL6VVDTIcIkvNYdwDcIClucVQgC4U11kkn6TXVGYeYjBOuH/EgiisVsEFyXCU3ddrRG8KCL5fYtilNpVh1L4e4ysAYxO5kz7vvGzCFdmpeBbLAxujXiQ33l/kUN9UZq8SX88Jn6D+TrcbvkDynd5lrFHM2jr2CfkYRHdthcr1u72HjQY2hFQAKHyP/7+GAxLvKYnGM8UZDfvSflBGC1//87xWoYL+xiFGBJvStJf8h56nAC8aCAkmmKYb+NeYrcy6BKbWysGzfbjJeLjMWXHsAuLh7p3umRuBHoWwSBfuU6aHXiXGrRY3Yj6gkFt93Uk06HrRQVtukclPKylEwCb/FPee+LcQp3C46fCa4p74PVLSdq++/+RXugS8XqNCpN3gFnIG6ss8AACAASURBVM//HwMVTV1i4MmXBVTsBnPcNO6NyDAcbL/EG1DRsitjQkwZFX6Vi1JNNcloCD0qckGHI6Oi7DMqFJgIzbT135B+Mkkkv9pXK+x18sf6jwVXgYoiQY54KqWMikqVkzyqkyEpwsrD7i5WX+JqSAN00k+oBFxdXZGGq56ENAdKPxH8TO2fIciBZDCqMNVks6YLHyodQXN0/hSW2MafBig0AFRUy6pLjnZ5SLsFHfZdQ/XRPgMBwuOoDiQSQKxyTyZdBXzCUTRDoGKgt4cb988+/YwVpUPDIwyEmGxKgK2BRI2OM1a5BBrUnuSMW+myYFf09UlntkNSGVBZk6yGVSmGdCBfgQpoJKUAVCA4qJXLbJ8BFQBOAFSgCnd9fUNmZg5KLyp+u7PsZxyzE9WwmUxQbWJVLaweaTT4HQuEATCgT4cHB7VaFiydQl6rfOJaDa7JIK20CxkVI3IKQAU8KnLwItGEowa6iKpDo3NL9ODc8KgoFbdB3GSSCO/Ry6QBHVFlVEB7HbJI+2f2U8qIQZ2rbuHvSyq/EQSgDvhjtYZ7kq5dvSo/f/oZ+f53vydT09PSSDk5DAJuFVa0o72scsEzhuDZgRWvv/aa1OhR8Zj0Dw4SqGAgWa2StQBGRfic4vlRRgWkn7791Lc1KUsz7bpUqkXKbLCJdWiQA6h4RxJgVDxxVgENt2lk1ZMged2Qi59/LvPzc/Ktb35TeiD9ZEkwekTX5OY1ZVSceey0DA4OaXAV14AQjIrXHKNifGxcE1uMDGPy/M+fkwcfeECmJ6dkbFTZFgb6WdLP36TieFGJAh8Ovtdl2VJ5Zlrmn6RdciUKBGluK2dKBqEAKqgh6jUeG5taDb4VIstLi/LGW7+WhmzKI48ck1znkCTiGenu6WPVPICAhmDTAEC1OfHon9Pm1Nbr50aKsCSSNXGJw8+hjiryZenuzpKRVW+gMrzttrit5RLOgeNCMUrHOYCKddlavSV9A8MEKor5Fc4Zh44+IpVGRqqVknz0/muytT4nR44elrHJ4wQqANY999O/lTOnAVQclnI9Q6ACAOMn596WtbUrcuzIPunN9clrr74hDz18TAYnjsvtjbp89N7HUi/tSF9fr9STKTlxCsbd2JxB4qgic3PznK8AxGbSWv126NChJpYnExwEbjRZ++abAEfWKf1UyjcIVCytrMnFa/NSr+3I4f05+fYT35CJiSPy1nsXZXRiigCzSgCobI2B1fntHdlYXaZ5djpZkxMnDktnrlO2C0VJ5SYlFu+QXFcXAQE8c1W2uyy5dE26OjP0bMB9r1ZhEF2kr0wjAeO8DNezYgngLzY0WNuS6nnQ2eHo54mAxaemfep7Qx1d5wOk7Dn9P5vr5FyOfgNQAUYFKt3x3Z1CnmyEHKSfCib9JLK+pt4I+B8Vg9mOLM+BtR+byZ6+XjIqAFSAUdGRwfqh1XwExgFUlMpy7dJVWViYlyEyKnqZWAEVHnNVFmyVZIbJbCTAUTm4snCDMQPW/HRG6fHUXSajQqSwvSOl/I500LepLrmenEDCweIPAD8AYlixxmdBgQp6NDF5IQQXcD4wKji/x2OytLRMeSYUKQCoMEZFPJYMWI0qawVZKZUsWlxaIsvAvm99j7WjUMjz+Jin8W9jVACcQT+hDfgM7TVASUF+ABW69uDf8KgwiSiVLWiWfQqTMWFCyWJGm89szvUZFQAeAJJY7BI13xgwhu/jWhEnUILEk+Dz5/QASEvCK6umgEy6g9JP9AOJKehRzKv0lV27rd+498mMMioODB39UhkVnNvuAxU6PPZMsEasxhFM9F3+BHdaqL0FPziTtScKqGj1QLCa1nsAKvTpuUegIqKvuPK29KE1/fcFVFAyhLGA99oDpOClmVzOne6Z+3wvUCrYmQYgRST844ZgVJJaq7JVVllPHJXQ1iLB0Iur+YjRFf5RlxsFVJiW/F12U/Mz5i7iywQq+AhFsF5sDmbc6Io1FLCOCbwdDZBWqT2nv+8Vw9i6oYl4Za23iz0teW1MOt0rtZfzRrKWc735CTivA7uOdsc3RojJKWFMYE3Evtrazv0VkvlVSB0J4xDEMXgfrE71NdACrACoAHMB+y1jSzk5MmOR0OPN5L/i6reAOMfWKsgU2fqMe6BFepqA172sKxJyoAQ/jycYN2mBDQqdsCdDzIZ9n0oK6e8VYLHqe3pRcBMU5zEMoFBgo8EkOtoX+GE4KWsrnOCjwbnTZMUUxML1o9iC8sEOQArlsnQeYTtcUp2+kygAdT6Sdr+UocGZxP3ps6HC/BiZ0PCoiAIqIDfsJL5svFFOLJ7UMVNTRoyxEyjJhZyR8/Gk2TWBBl0Y2GWOeaF9YDRsSIYpSxf5BxYEkqnSYFyHflVlAtwvZbbwOXKFG+gHjGVIqKIYE+dF3kXZO+o1gb5FfATmMcYmGEG4H+gD5HPYbsfe0U7zZ2ztd3+evQ9U3NOse//LX4UeuHegwiIZb4FpWu1bkhz8TKtqm1H+COmnfzaMipYJhd3SCuI0j5B7Z1S0BgR2fP8eNCPWukDs/lwLUXYnqNRMN6TJBkCFM8eClAwWBZUtgmdBkYbElH6CoWIg/RQyKnpHp7gZx0JjKDXGhm5EdeFVoEIZFdVyiZITkkhIprOTwRNZEwANimUm2LMEKrSKwD5DggvVkKsrkCxSmQcCFQgCEgnZN3WAFYykMGKhuANQ4VeU+IyKgYEBJjaMfmmBgyWdjT1gSQLzf8D76Af7HvrDgAokJczI1CoBwAwZ7O/jNSlQEaPckVb/x2Qnv0XE3mSjtPpQU7e6GXIMA29zh8U119UpPf090tPby6BNpRhADdVKRyTi8T6ACoBE9WpVgZl6XXZgruoMqNfXNmR1dU1mZmalp7dPevq6CQQhOWiyFhbo+lW8uD4AFRbYYWHG7yDlAaosEpi4f9lshyRTaratJmBa/V0uqeH10MionDql0k/QWeecgypfaHUjKHFa5wYiGagAaatyaUcAPCGYCIGKhJSd9BOAijNnzsj+A/sJHuCFvkOsDRkrsErwsmPak83HCsF7oyEAKp5/5mfy3X/zbx1QofeHcmWQfnLJZwMqwFRAUgyP5Zuvvy7lfFFOP3aa/h8A15gUrFRJRa2g6pjNMs3QmLzw/AvSkU4TqEASDwlM6IpWqir9xG/XoXFekXfeBqMiBCrwTGhli8oT4Z+fffqpLC7Oy+lHH3VAhasEiqt5/K0bNwlUnH70MRkaHFIwk9deJ1DxxutvyKkTJwRABYMr53NsQMXE+IT09fRQmswYV5bU8mfKVqDCT5rxHnzBhZdswYhX6zmiQAr2aVOVHlqrVT6QfurMdOwCKkgZxlReS8jC/C157fVfSCpTkke/8S0m3hLJjHRme6XWAJCACi6VQ2oCUvxztjAq/I1jI6bVpvC7wP/YYnz4wduyb3JYBgf6RWKYS9r3YDuPCg3oMUxVSxdARa2wIoXNJekfGJbFtR0p5FcoxzVz8CGpNuC3UJaPP3hdttZvyYkTx2R4/KjUY31SKRflF8/8WE4/9qCMTx6WYj1NOSkwKq5c/liuXftQjh6ZlLHhcXn3zXfl8JH9Mjx5Um4u7Mj773wgO+u3pa+vW0anp+XgoSMBUAEz4AsXPuXmEY0FuL1vclyOHj3qVRDqs0PKPSsME/LqK78UkbxMTu2TzdWSXLt6XS5fvyk3F1alMxuTg/s65TtPflNGRmflvY+uycjYBAFOVvXHIFujPj+YX25duyKXPjsn9fK2HD06IxMT+6RUa0ip2pBYGnJPCiDADwF9CqC1r7eXnhaqhBmTbQAUFXgGwR8pLqlMVuIGVBTLrNTD2MA5KdWTBVChOsWWSMe8beuugYEGGGhyIgQqsJkFUIHNH/oOQw4FA9h40aOikFcz7YbI+joYFbqhw/XC4we6yvgdNnpdvT2ysbVBpmVPT7caM1YrlIDChpwFCKWKXLt8VaWfxmCmHXpU4NFEW5LxFGMBrCcAMNaWbjJmwDVgzTQvDm6iIcuXz0ulUJAUkh5SlyyACrfpw28IVIDRkchwPYNHBfoL/kr0U2iokbWuXwq0Y94CowJgAtb+JqAiriaRjCdwXZC1IsMmIQuLi1znAD6grfierX0GVOD+YD0FCILfYRxgU7uxvsHfACwwnwYmK2Jg9IVABeUh02llMihMoXOt938rEMHItCU+twQI/gR4YECFFTD406QVaOA9q9QEk6YADxMn/WTzpcVQVhFpchwADo1RAR8SzHta/Rj3gIp0oN9tiScAFalMglKT+wePfLlAhU8ybioM3zuhqgvr3SxCd/WluznQHYCEuzuEttsT3m5adPdq6z8NUBFUjipJNHjdsdewxnE9DL9pxQF8Nlu6g99qs/RHARX6/h63OKqaXl0cwutwzfPNj/3PfQnL5t9FJezbvb+39NMuICGQpFcj69YX4sd2ryiwpfX4QTe35iut4jo6BGuKq5r7Q4EKvCilGiRbvW8FsR11XSLlufYG5Nr0RwQl4J6BCg9E0FSB7oO/CKOitZUGUESBN0jAEqh3yXYtgmmwlIUMVBfTGpvNNPXtPOp9oHsAeyp8MNrWQ/vT1gusYyywavOyanKTX6QXguuXtj9w48kKKFWqGYU9ChAGCWTmFpTFbodD0Q6L4BQ14DXAfxExiu+pxH7wZVsdOEZWuZPIIugDOamiypCib6xwiFX2brzoYXSPxTHrciwai6nZNPbBlGliArvsPCPqgQQT4hhIDmNvR8aG2xPiyLifOBZyMbheSGHhXpIhgaIAeM24wk5fEgttVS8HlbwyT0kkzW1/bvtn9lEqpcAO5YuUOWnJf5yP7A9XwIn+VT9Bu4N6/SHmrDkK+wI+/VtP+slnVGgBBv7XfAdzLAAKuA/Wokz8G2wZ85nwxw3AAQI5zufEbxHaQA8P7BXKWtRj145j23hSiSm9H/g7Yjuwe2lCXoPEso4plaB1wATjUC3sM/DEcjS8JhQrJhRkYh7LMWFMRsyNWrtE12wtQNPnFFuAsW/dcY1s+xDdf/N+D/yB9sAXBypakt3Bk/HPE6hoTVTZ7YyKq6w7mgI4PxHWFhQIjxYV+IXDyELl1inJjrE72dR+8rIEdhugwkxVPaBCFxZdbDCBs5oA1ZmOUVEmUFF0HhXwqSjsYlT0jU0zsUudQ8/cWIEKlStg4gsLXL3mARVxSXeEQAXR6GKJCwOACiRFcTVYtMG2QPPh53AnoIL1A3cAKhgEu+DHQBmTfhodHeVnFsBZAmIvoIKVHg6owPf1mM2MCtvkE71PpQhQ9Pd085o+/+wzVtgOD4+w0hQMBGwiVlZuM7GA4yOpYYwFamd7QEUYeODCGpLuTDHpgkSJD1QALCD45BgVqFxFVhVJFKyW+UKJiRVU367cXqP0hAEVfQM99A8ho4IVqaiSRHBa9eilmtxAX1gCBtXEODZM1JEU29rYpFzMxMSYDA8PSDqjrBFjVBTyJWemPSInTj5IMAHSJAyDWoAK3Me9gAqADgZUwGC4Uq7LM88+wwCEQIVjVOA4BCpiwsQczd7bGDf7QAWkn+BR8YPvfk8mJ6ekTkaFAhUA3xDcqOlcyKhQW4KYvPHaayFQMdDPa2O1NmS0qug/iCzhudE4jR4Vzz0vnRllVOwFVJRKVXnn7bdopn327JOSBFXZmWlzlnESOgZUPP4YgIouDYywQREFKtsBFTXKCyij4s033pCTx08GrIlWoGJ8dIz9jHGI8d66IfKDSX8u+22ACh9waL9l0rN+UaCCv42paRx9KrLOp0K3SSqvFctLAyZz1Yw0qkmZX7guv3npp9LbnZKzZ5/QZH2yQ1Id3XCiIauC8kReTNEERrQkSsLPAA5p9U2M3g84TlWef+GnMjM7JmMjI9LVPfEFgApI7OTl1vy8LC7PSapRkKmxXhkZHZOljaKUi+uUMpuaOSU1waaiKOc+eF02N27JqVMnZXD0kDTi/XzeAVScefxhGR6blbJkpA5GhcRkcf6ynDv3ihycGZODBw7Jxx+ck6mpMRkYPyqXr6/LhXPnZWd9WfYfmJKZo0ekM9sNhJAVUEg0X758RZaXb8vg4IAsLc7Lo49+iyyF5uo/XddwTzAuXn35HyWZLMvk1KTM31yVy5evyueXr8pWoSbd3SmZHk3KH3/7URkYnJYPzt2Q8X1gVGSV1RADUwASACW5cuWKXPzsA6kUNuXIzJQcPXJIGrGUFKpJeleg6gvgDdYzsA0GBvqlu6tLk9hljMq45ItlJ/GTlCI2X8mUZFIdQQUZNo2QijKKOTyFKL/kNlHmi+QzKsgYdAwuSyC3AhVYW7DBhv8QXvlSgewFABVIrtNMu96QjY11tgVjulAsSC4L2b6GMioSCUourW+ts5Kv15lJGyiPjTMks2plABVXZH5uPgAqTPrJGBWpRJryU6hQwzq/vniDQAXWEDD20OecU1FVFwMoVZbizjaln0BbynaDUaHVdaj+wxqZSQPgyHCTuLYOoCLB+dKS9ZAzxFpsHhU+UGFm2gT2wfBzBpqtQAX61YAKnjODJDzWImUTQvoJxzevK4AguFdkJIjGMeZR4QMV6BeTfjJGRQBUKGUuSIJYwsRPIgVx7B5Ahck4GaOiFaS141rcg/7Db8heApPPZC48WSkcQ/WyVY5BNbQrZMsAqMD9xb00RgU8KnAsSxgYUIHfmUfF9MDhewcqbHffuj/jutvyZpBcvYs0wF185S7RjLvbOe7JeLi7Q7iFLpDKaPrVF2FURJw2usre7zRd3VzOyS3CYQQQ5PnancMVV/kf+UCFrrzhS8+6u1X6nd1V9ncEKiK7+04Gz80/jAIqog6/p0eFZQ/96/akn4LErfu8HaCjj0pUlBRxV1sBiTZlcs2FHa7P21xk1COlIGyz9wdlWILkdngwxtoEWzRJGowFd1PbXsUez3IUoyKS0RHl5eFVRRujV4EKPXnbPMNdPvMGUke1yWdUIHHL70NWB4V7qMJ3yVKd97HWuqS+i4v9qn5LCvt7ITs/q/5R0e72YHsBFZQodawHxDRsC6rZIxg96AplQOpemmw8xxawpLBej5MGUi1V7jsRJyF/UaV0ZkwT3PR+UFaAMiLMNN0BIM7vQY3YHXCJ9wD6wEwZbXfvk7ns/CLQNq2Wd2CqkxyyGUgLQUPQDfkVtAVqCYgv7HzKCFF2CI/nzJe5rmJ/7fqayXQW4Oiza4CP7p2daoUrrDAgiUUeNDLXduA3YFPgc2XyC4EUSBKjT3FN2P/jPRQFIveCdqMvCHS4YtamuCGYVluUHgIACcxVkf/imWn/W+dREcwQDQmKXRBna1wULtroFwOMyPZB3OdMt21GwBihP4fLzen4UuCN+3HE8ix6UZCKDDQHLAXXQzN27XfOKgYyOu9T9JuBOuqRoqoNuJ96n9QLRMenCpijOWDTKEOpwaJNAB/4+27ATsdmcE33gYrIFfj+B1/RHvjiQIV/wW5y2LWgW0nSV59R8UWBCg0yLMzw/D3aAhXNAdXeQ8pm9JZOj/QXscqa1qPahqAVYEJbQx5wGJC5Sg8XRBGooEeFJlvgZ9AMVORlGybaeZhpA7jIiwEVJkFhiWOaTiZ1LBGowMSPavEypJ92pBFPaIICaLWj2ylQAUZFtzQg0+QBFSgHR4XhHYEKJ03ABQPSRhUYian0E6h7vIduk41FSwEF6Ogj4V6W8XEk92BOqhUltmG3oA7JGQ3QdJFDpQYCDgMqcP0+UIFz+PIQmvSAnMeW9PV0kdnw+ecXmRgCUAGZBIAlyRRouWUmNZaXl9luSC4hgEhAu5wsBF0EjYLJwAfmg3GlhSJBNjIySskKBCxYICuVEqsj0Y9c6B2ogyAkXywFHhXLSyty+/btAKgYGOojnRaglDEqLFFGPXwHdtm1G4ujjP6PxXjOQmFH1ldXWWnc2ZGRmdlpGR8fcUCFVvAiifaLF34hg8PDcuLEA7J//37KhgReEmBUIICB94irYjXQiUFECVIqeTIqENjgfqhHCIKKujzz06eZTFGg4oDqnjqpDUSAZJw4RoUF4n7FDiWcGpCOuSrP/MPT8u+//wMZ37dPYjDT9oAKY1SwKtXU4aBNKkKgopQvyuNgVACocPegApCCQA/GowbULAwSkeecRwWBCkiZIGhEzTsYFfWKo8uj4rsmb7/9pki9Ik+efVJSNCPGOLYKGA08dzEqnHcNwIgooIKhG2i6pbK8AaDi2HEBc4JUZM4vofQT3k/EYpTAAasCz79tavwg1yBam8m+KFDRCiyZR0W7efe3ASr0ZjYIwvR0ddMLR19qkF2PbUqjUZJGtUMatS5uEufnP5fnfvYjGZsYkae+/R2aLSfSOcl0AIBLaTLdqxilLq07Zmv7mxkVSm0HUIH/4fsyN39J3nzr1wRFBvpmXKLKrQd8iLTH26UoFLTGXF2SldU1efvdNyW/MS9PfOshGZ+YlOXNkpQLa5Qi2zd1QurxTj5vxqh46KEHpH/4oDTifVLK5+UXz/6YBtX9IwekGuuURizJ/tjaWJD33v2V7J8elhPHjsu5jy7I2OiQ9I7MyoXPF+TyZ59LZ0roeTEwNiYSR2JagYqlpdsyPz9PoGJoaFBuLy/KE0+cYWU7Nz3Bht+ACp3DX/7NLySdrtH4/tJnN+TipSty5doNKTeSMjzUJaN9dQIVPX0T8tH5W7Jv8gCBCurxx+KysbFFkOLatStSrq7J+FCfnPnWNyXX2SUb22VZ3ijJTqku6WRV+vu6ZWxsXHIm9bOxIZub25Lo7Jds1yDX0GKpIrFEkubceJaRfMcGEgAHNkJYI1nN1RAp7OxIjkCFyh/g+cc1mbEkrhtzFmn9kA10wC/+Ddbh5sYmQQWw9QC6oOAAz0u+XOQaAEAF7AjM69g0b2yuk+2AOYOsAQA2ca3Gx7qS687J+taalMoV6e/rc0aQKsnA9uE45YpcB6Nifo7ST93wqAAQWlHt7FwuS+aDmTRjk76+eD0wvURS3wADAhVxzDslehzlKFVYppk26JqsePM9KmDuDYaGB1SgT/DsAOjCsQ2oQJvAqMCYwjwFvyeVikKSJ4ynfEYF2rPYxKhQIMSAinxe5azQ38aoAJiBeAcvMFZM0slAJ6y/OAZlHCAjkEww3mkCKtCDTkbBJDfaAuptgAqLy+B3sr0dSj+1mx9ZtOK0qNE+Ayqw/jO95cVP9ntWbToNcN2klz2gAmAFDFGVUbGztcnrMjaqST8RqMjEyaj4wkBFFP3hPlAR3urfAVBhyRZLiGrc3UoWCfc7UXsy+13TODWmQMR1MB5tlxB2329NFLfGIHvv1cKVOUiE72E+bceKBCqiJLXor9S6CXdwSzugApEA2MltEvH0tOPi2HJl7b7cppAjjM3ctUck++0afTwjCgxpBUj9+M+SrMHcYmwELxEciruH3NCmpN9e9ySKJRPBqIgam1Hvm/mxjl2deH5XQIWeMzRWZqIVawYS2ya5ZM8BEuEuCR5I52hrVeoH/hBNngQOaHG/U7lCle1hspbFDe1e9jQ6r0pjAETKyYXnYbxLzzRtv0kU4bpwXvWc0MIw7gNdYhnrDWILyiah8h3JYjIQVNKHyXm3JyEA4EAR9p/t4+o1Hh/FJ8o00TgL75mso4Jlui7zFVDHNO7EscnIQf84c3OMWEodkQWg8kt4QJFLQOyHa4E6BG6TVuJrIR8S31bwZeA+8hTcIzqJJEvgI35AX4CBDCUFSGJqMYuBGhqHWVyEPSJiHMoh1WvOiFp3CVqEWmdBBsET+mOEwJsbMrtgS9urkJ2biMn//b+FE8f/8uchm4tJfDIPtECUMY0zErdHFfcLuSj0GS4YLAkwTJDbwHsoqIEkAu4HC2TdM4DEAfqCuSSAE07pQMcRZFnV3NyeG3zPnhOMDxYKOvYM2Rb0TYvzfOgT7DtMqsuec7ChEfuZb5wBQNbXVuBJMNrmNG/cYBK3ueU+oyJiSrn/9le3B74QUMHkk1UjhCEcsb49qg/CXrIkCB/14G0GIkGVh38gL9HPJzvUovSpYs13wTfJVMmbdkFCUwLMLYZRy2Zza9tG0d5P29VA+O+1+fwOi7DOjHaK5lKVEN2NOodKyGiFUFTb2rVJzxP2XdiP5lFBoIKMCkg/lSiFA8knM8/G4m8gBd6H9BOSGSEdE6pO0AJURJ7dQAAEi12ZVQPYrGLBNJNOLP4AKAwhB6MCCxvBASziNFNKyubGhiwvLrKyFCbNuS5UJWvZ+f6Zg+pRQfMjBQOQLMF58TKvCw3ItB+wwKESUFkBGmxNTEzwT6tQ9SsXkZRTZFxBAq3YUI10/N4ksPC5skw0yLDqRQbgLrDBdwf7B5gguXLpEq9hZHSUC9/Q0BBBAQsSkDxHYgTVoEh+AXDAcShRRVMmJ4vEKlAdy/qealiOjIxIb28PAw0keNA2JEEANFmyAMcqFEp8D58vAahYWpbZ2UPS298vwyMDkunsCGQjslnVb0ffIe1pGuAwwEIfaUWuSLWBGv06aZvra2uyvbklq7dX2H/dXVk5evQwzbrxb4Il+bwz0x6SQ0eOEqgYHBrisZjQcEAF+tLGnP5Wgw2VftqkfBLOiXGGpBGSJHjv2WeeZaLq9OnTMjM7q48PghFSexuyubUhG6trrChPJ5KS7ejk/UhB3sOdB+eGUewzT/9U/vRP/5TyVAIzbQv8qlrha4wKVKEoE1nnrldffZVB1uOnT9MwGIEuk5IuQYTnibqe9DHAoRP01kAF/1NPPhlWrQoMeMvKVgKAUhce9523wKioy1NPPeVowggqHSgJH5BGVT69cEGWF+blzGOPUb4Fm1xIUNEIrlaX61evyoXzF+Sxbz0qg4ODyp6J6ecAKl577TU5eQzST2OqAUsabV1++eKLcuzYMZmanNTEaiopPd09TLRizOuGxpnPuf6ImsujNrM2a/o05Dt9d6/P9wIudrUN48Ul+UEFUwAAIABJREFUSlBNjvFhEimQO9F7jbHpDMy5ya7J3M1FefonP5RTp6bkG984IdV6QlKZYYklBkFOdsbPmC8o0uUuEX0a0qnxZnPVH+Y2fFcZFdVaSeKJsvzshb+T6clJmZl4gOAmE/11mFljw1CRWLwojbpWzO9+YVdYpfTe5vaGXPjoTZke62Pifmkd/jaLBKCm9j8olZoyKs5//IZsbdySkydPSf/IQalLTiqFLXnxuR/LU08+Kt2DB6RUhycA5qW6FPLr8tKvnpMD0xNy8vghWViYk3g6JT1D++VTgAjnLkh/T06OnzwpXX0jTt4vRZmkmzfmZGlxQTa21iWX6+CG5aGHHuQzbpscJgUY1oBGX5VErCQv/vIZGRjoldHxaXnv/fM0igcI3NXbJyNDXdLfUZGnznxLsv0jcuHygoyOzUquMyNSK8vN69fk6tVLsrS8wmr5vu6UPPzwQ3Jg+gCl1lbWtiSeSsvQ0IgMjY6QUVAq12Rp8bYUCtgIpelFkesZlK6eHicLtcW5DBtJst6SSPKrvADeA6sKf8e8hnZ2dymrAd+1BIF5KVVr5SYJKNXh1fk0l+2RtbV1fk4JIRo2F7nR3CmVuVkHmFjc2VEvCgBJWxvqgSMNAhiQrYIsATwtsGZiTK1vrvM6+vv6AwYinmt4eXRk1Ivh6tUrsjQ/L8PDQ9Lr5ByLDYCwwr7tSGVke3uT3kUoYlhdmGNxA+Y+ABmopLTKSq6pACpcZT+eOZpRw6gTMgjVqmSz8KhAAhzSjQAl0Mdx6ehIq5loAwbbKrsE6SfEFKiyAzsChtdgMhpQoXGSalsDSMI4o4QR5a2S9N4AcNPX28dzMJxzQAPiG5WEUr+p69evB4AD+n1jQ4EKfCdkVGD9ikl+p6iM0GSSjEbcY7IPeE9DcD6o4mx5gG2NsWSfxsqIWQBk4vgFep50dWclndY12s/b2XHtT/Q7rgdrkslXWoJDY3wsPWFCS8eAgqYARVB4gf8xlpOJlKxvrLNggQkGB2z5QEUa0k99vTLVfyiaUeHYpHbpYbzcZjrTK2wrD2O7nra/ikrmt5syXSe2q+DWiuo2P2IIelcbrLB5d1l1HdULTe9HHuve2nR3jAr/Etof3wpvNElq32/eF2k3h8l4jad3vxBv8nn096MR3c3tyR73Ibo3Ij6J6FfGCPqwBK3as6dd0UDz1XlXy9yvd4XcrjvmgXsumaBuC3i4nfY9AhVBW7yGB6bZbe4Ffa7qmhC921ckKOCiFa2I1twEJVi4Bw4T24yRAvaC9Yea1urXdvd6kBSMyCugUpryMa5a3fZckbNNi858cE3GDHH3zsazz/RpTWbaOSx56uc+mtrt5qBAus/F1gZURLdV1xSLycP+d14JjrmA41jsGXU/UWBFqUznp4Rn2goYbX+GddnWdDumMSN471CARikg3UNibbdrVhkeraYPwBG7Z46FgWMgeQ9GJvIYhj3ZPGXeJ5Q3gpelY1EEvhUx9YO0dqMgCZ+hgEMZDWHiGsfE2heMC5fAV6kmBSKoVJDPM96wvT/6IJzhwvFoDAxjBaAdzCEApLB8havEZyFmC/CqcW84f2KNRR7DPBJwDSpj5uSQbDxjbsI1u3wFfkP2p8OXLK7GGMHf0XeWbMd7AWO+of2J+BJ9a7kWfBe5pB/9Z3jm6eu7f+FklniNocm73Wv0OfzUrCAUbTdmickrcaziGpzJN8zAteBD7yFAH8R4Zm4OsEbzFcqwQIxroLbKS2kM1iz15AAxsHgJYilTQp8TL18aMe8TEKNXheYAzGib4wvnTMRZmBjkrHgv4ipDhd/cZ1Tc7dJx/3tflR64N6BCdcU16+KH7Pp3XdPvJsD43QAVtqj7dLA9E0y/d6Ci/ahpanNTAOcvWPZb6/820k93BCr887vjmPxTMKn+9kBF/8R+Vsvbwo6zBhtPVFxwJ6CmRLUqgIoyN/hYlNWPAcll1YC0agFIS8SIgitQAdpoOpmiVjeSVKjKNaCCmT0BUDEraZh66j/VHAm+GZjsXWUC/vSTpKwYAVBRUfkitNGACtP8xv2yIBELON63ZIBuyuOSTGngpAlmpR4qeKN0SiQkzOAKn1mFAhKd0PC+evkyfzMyNsbvQi4HoIAl4y0xALACclCgYwLkwblU+9nJIgUsC2c87RLCCBSQhBkdHabJLgIJsCXMbJvyGOk0ZSfwHhJli4vLsrS4FJhp75+ZpoQGkmYm/WS0V7I43CayVgXIowErRrTa/aqvARIe66trsnJ7RYOBSllGRoZphAvZDbQDQNjzP/+59A8Ny5GjR2V8YoKyLsrQCc3Fcb69gAropcLUGvOFSrggIKjKMz99pgmoMH0lVrsI/DV2ZPX2bXnzrbdY5TzQPyCzBw8yOYfkLTWIGw25fvWa/NQBFZPT0xLbA6iAsaifQAJQgSAKrA4wKqwS1a7HpNQ0SR1rAiq+/dRT6v9Co/q6lKoVBSrcXFIsO6CiXpcnCWpAz7QFqJCqfHr+gizPz8uZ0wpUQFoFQIX1642r1+T8J+cJVACoYaUONWK1X19//XU5cfQ4gQo+IwiQ4yIvvvgi7+fU1FRAzYaXAxL6lpTzN1j+xiuY9drIbrWbTXWz0eyXFLVW/1MAFWAsQRaHwTKHBTbO2odWYazzB7R00/L5hQ/kpZeekZMnDsnxkydE4llJdwCk62QSUcEsbDSs2gh0qTsAFXj2KP2EpCOetbLML16W9957W77+ICSRhuh9UK93ijTSEotXRQhUaFDe7hVrgNkDkCkmK4tXpLq9JuP7pmVhLS+Fwrx0pJIyOfWgVBoAn4py4eM3ZHP9pjzw4IPSNzQrdUhC5TflxecVqOgdmpVSHYBOVZaX56Va2paPPniLQMXXHjouG+urUqpVJTc4Jec+vizXL12WscFBOX7ipGT7h6RK2npcCvmqXLt2XW7evE7JuK2tdZmdOSAHDx7k3GHjwTZrdVwj9bh25Jf/+IyMjA7L0MiEvPzKO/LJJ+elVqvIwNCwjA33SHeqKGdPf0MS2R65Orchw8OTUisX5db1K3Lr+lUmyOOpJGWnZg5MUpJuaGhMOrM5GRgYkoHBYSZWt4ol2dzaodfO+uaOZDq6JRaHt09Jenp66R2E9Q5rINqM+VbnNgW8DaiAni6Syxi3kAns7obhvW7AjFGBzSQ2xPCPoM9SHZV6yvjTZHdKsp2QF9zg+mTygdg443ndKha4CYe3Q3Enr2sKgIrNDVanIfxjMUJPL9dHsDyw5mHdhkcF3kOi3jaw3LQCqOjIBUDF8sKCDA8PSm9XN+UcS1IlwwusCJhiQwaoA+aStYqsLC0ECSHf7JnrG0EAGFVrwtyACoAGlCuoVZxBN6SHwAZpyNr6JvsVQAU3+w1lVBhQgUQI1ikYY0OeyRgV5gGizyEKEiD9hapEsDzUO2N+/hbXKvwG983mFzAiEKeYdwX6/caNGwFQgWd03QEVdj8UVEK8EyegZf+Gmba2tUPPEXfJOQfSt4t//XnO/u4DFYV8kUAFvKzaARWW7GgFKkz6Ce3Ed2yM6Zy1G6jAOWHabkCFGtKnZG19jWssQByrCm1iVKTjBCr2ZFREARXBxqV1VtsNVIQzXyTycG/bvr2Ahy8LqNAg697aFfXtPziggk+5a214jQo469uamNK/Uwk+wiz6XoGK9jCWO2dE/0Vx2iMT7X717F3cQUvCNX/V7c1dwZN2RNhn1boyMdUnw74LNsVu8WEFaNpLP0VdQ9CW1iHoDGtbnyR8TauGdf62117Hj+w/G69OCpUJxYABYYMi7B+tcP9ygAommOsqbYx4Gm1kUrfNcx1Ca34nWfLYjV8bt06Cxr9mf59gCdxg7Lt1kHGOV3CnvgiOtWEAlwEV9n5EtOcX4vljTeNZ3fviT2MumMRj07h07BUr4rMENxPVdWVo43hafKUJYe69HaPBAG8CF1BBYPEd9tVJFkpyL8kiKlT7qx8DWfVuPjSgAG0FoKQsAx3zKC5rzbnw6XDAS5jcD9kPJoelnhQGtCFXAKlkZSHY70yCiqwltw5aISNNlp08FZpKTwkAP97c2wT0OmNvu04WpeD7TuHB2CIKAsSY/Na9R3iNliswcIFFg2SdmhekMmAATFAKzBU5ElQikwKAhcptA1yw59ZYJtZemnk7kIZAkzNTV5AJ909jUPQT9o5gpfzwP2kxIV7f/XMFTTTuUUaI5lxiPBb9JmrKPMHYthiLEks2bpy/pHp0aHIfMSuNq+kLosU++vzq/eEYcabsvBYH8PJzl0exNQd/Ejh0QA7lyryphuC6e75MAaF1ajfwyQplwmIqbY8BPnbfAK4ZOMPp/T5QcRer5f2vfKV64N6BiiDqc8GfBTg2HUWZbDctaV5E54X/XzKjIjyjq1DyJ/uWigquX79noEKNq9u8moHYIIT0FyxdYq0v/fDPC/Y4ybacYw+pKL3B+v1w4d4LqKjQzyBkVBSUWbGzHUo/FfIyuG+G/zZTT57GbbxRAUEDK+oXg7lQllq1wiQNrq+zQys8DagwcABABZJCBjAYUIFE99LiIg2gfaACt3/6wKx0gIYHaRZKMsGMCZUQWtluzIyQDaGIP9qFZA1ACPRLFKMC30WFPpPJoMVikYrDNDxBoAK/Rz9Y0IS/Y1FCVYP5OdhnRudEYmjBMSoQOIBRge8CqEBinLrPDviAPwT+DtmG24vLNMRWOQVhEsSCN1vw7E+7H2g/EtL9/b1M3sAoG7rkSB6orAWooRXHqCjJwvyiLC4syoGZWRqhHj5ySJLplCB5gjYa+MIgJamBAIPaOioQVM9Sa8NrApN2JLdx3wlUrKxIqVCUQn6HAQiACCTD8SeSMj979lnpHRiQY8dPkA3S091N+SaTA7F+VKkyTer6jIpScZPBSrWsASsALAMqWhkVkH5SRoVWXeUL25Lf3iHTZXR4hGMQ1wuQAkGvBSY3rl2Xn/7kafne974nk9NTBNYCRgUCmio8KpS66wMVaCuAikKxSFbHwNAgx1MaVcBuM8TEW7ksNZpahEBFNxgVBlRQsgqMCq3WsJkA/37nTUg/eUAF6bwho6IoNfns/HlZmpuTJx4/vQuowH0kUHH+vDz2TWVUYHxpLUqDzxWAiuNHjsnE+LhWqFBuISYv/kqBikkwKty8jO8vzM3LzMwMAam9GBU+8NAOxPBnVHs2bIz/LhZrreDT2Rnspu5clwNL8LbpJSuI5m/0uJGpN+STjz+QD95/W44ePySzh2fIHEul+yWexFzoKnqCKkhUj8KfJ5z3mxgVMZwP/4MxoXJwlSpkfary8ssvSq4zIUePH5Rstk+k0SXS6KAsXCxe5nMaBVQgGq9Td74qWys3pVrYkNGxfTJ3G6a6c5LtTMvk1CmpNnKkYxOo2LglDz30kPQMHpBaHUDFhrz43I/kqacek77hQ1JqdEp+Z1suXrwgnem4XL30iYwM9xOogKfHGhLWPWPy/vufy+r8ghyY2icHDx+RRGcP6fsAHgv5ily8eFlu3bop/f09ki9sydcf+RoT7WFS1tGmWXGpesLF/Iq89OvnZHxiXAaGxuW//8PzlG7L5jpkYt+kTIz2SbK6RqCiKCmZW96UVDwjczeuyebabamBXVgqy4GDhwWeOwODg5yXRkbGpDPXTRCqUCzJ8u0VKVQb9JxIJTOyuZ2XVBqG3AAqiqzWBzsByXYDKgBKqgwONu/YBKuRX7lUccyAGud8yDPZPId5H+MAf2plFowVUT0IDWSVYFKgIinZzq4AqIAEockOYmxu0DfIMSq2IS+V4zG2NjaAj3F45IsF6QZz0XlU4LiY+9c21plUwDVZEoPAfQKyCCGj4vbikoyMDArmLgzjYkyfixwq7dMpygBlIN9QrcjK8oKkUyrDgHtqbD+bExAnYF1tAiqwsa7XOA/CoBvzaMyx+VZX17k+mzxAW6AimaK0IgyvAbogrrCiAmUraWIChQ8EKuiB4QMVPaE5I4suHFCRy1IeDmshgQr4YsADRGoE+5GoB1Bh16b3LC5FmKsz2RiX1bVVrnkEKpK6Plk1ny/JYfOeJmc8SVIXi6mMB0w3Ud2JgoENyXWBUeE0ub0w0uYXW88Rl2w7jwq0wyp+W4EKH9gAqINzggEKoAKSV3gG0IftgAqLFxEL3BWjoo20lfVB+/z77lg8KjwP15B7BAR+V0DF3hd690vg7xWouMu+bfM1lTps2g3uuuZWoCLY1TZvd4PffZlARRSQxFjIKwgMLiHqPnigjH+1GlO1bCJ1V+cKTTQhaQU1ftV1K5CA+fBuX27nGMSZTceyJrUezFV4+8yPIJG/hz9GuzYFCeUWOMuHtppgrqCy3M7Y9GnTKSxOjYo3mah0Wv1IorKS3qRp2jE0GJCG8i0+Y0JvlQ/EqYSOJVHxMdYf2wv7cY21L2Tw6n0nd8gBC3p4PX5Y1Om3pbl3rV9397n+xuZ7S+xb7I5r2PV4ujjVjmnt1UI/NSI2mWBDHJV9p+x3rDX4jSaiG654rsTkOeVlndyyFQ7aWgX5VZOGAvvcPE20ELE15xGCZn4sbf4d5oWhbNY4cxP8ezxBhob2dahhh+9zP+rkg3Hf2FYH8LC4juCJxmXaNisE9sYBTaw1iY5jkUmC/5z8FgAHjRE1J4e24/s6PsIxHppq62f4Db7L4kHH8NDx5kAEA7ycbKh5WlgRIoEp17827gxQQo7FYk6VsFQQQe+/AgZoHeOpuMj/5Uk/fffPlTGgahSQ2FIvEesjyMvi3oFJgfNp8QhAL2UcKGigZupWpGSgCH1NncQXj+fAL/hkGVDAvEXKgTJg8TolAZzDB+fwYDE/5QpileVj/ipOucKpCbSdt1gkqLJaGlNBslULbcw7RVlQqtABcIXPLu9L/T5QcbcL1P3vfXV64AsBFYz6dBEPE+RtgArrhl2rkwsA+P59oCLspohg3HVRU41Li3YrKuv84HT3311ozUp2L2SMBCrcEexW3RWjwoCK0p7ST0OTClQgseonDrFAILlOGltN6YLQPgdggCQNmgCgAguvD1Qg4Ojq6ZZEShPd+D4WHlS343eLCwtMaiDpks11ScMFkPsPzEq2Kyf1hC7uDG7AlECAgAQe0HqaiZlsU0hNDBLDtZrs27eP12GovS1aWCwtGWSBoNIeIdmh1QcGVKC38XetwAklHizAwnEQkGRSaSbEwajAv8GoMKACjApLFqAvtXpW+xFxifUF+p1ASApsA5hfaUUCNwcuGDENTvwQFFQklwDOaLWK6orj+JYIKhZLsrCwJIvzC4J+7evvlUMAKlJJSkbhfFbxijZmsxkyBAgI1TSYIFCBYCVWD4AKVKDCTBv+GDvbO7KzvaV6mI4pAW+O6elp+c2vf025qRMnT8nwyIjqeXd00FTbql2tksWCTR+oKBbWSfnF/WeiP53hRqNSrsmzzz7LBN/jjz9O6ScFKmIcp4jjSqWCFHYAyO1Ib3cPx4wrdWfylhuBel1uXb8hP/mHnxComNoPRoUG2ax6QWCEgMqNGWOc2KbjlVdeYV+ffvxxAhUYT5Qqc8lt3GeyKlqACngiPHn2rEpwGKOCgbECFThOqVKW995+h+Dg2bNnJZPu0MCKxTcM9VnVDEbF4twtefLMGemG9BMhJZ2zKP107ZpcAKPi0cdkcGCA00zNVZ9U4VHx5pty7PARelTYJhZbCUg/HT16lICfvYr5gpz76GN5+OGHybTYiwlhfaQJvNB/5U6rsP0u6ntNVVUtX2r9rf9d/zOTVjCgAvRyjBFN2uGgzjPCsaZs7qBOcwPzGMakyPvvvSeXL5+XE6cOyP7ZUYmBWZHuEYlnJBaD0ZpWISJRGqvHJY4o372ar0NBsJBRYYnHuszPXZWPP3lFjh2fJciQjPdJow5mEeZHJIuje7RRhUh+CrbqsrVyQyrb6zI6MUmgYmvzqvR0Z2Vi30mpklFRkvMfvS6bmzflaw8/It0D+6XW6JTSzrr88uc/kj/6zuPSMzQr5UYntfk//+wTGezvlls3LkkmJfLIQ8eZMF2FHGDHgLz79nmp5Aty/NCs7JuelkosQ+kdsKF2tkvy2WcXySrr6clJV3enPPjAqYB55veNFhaiyqoqq7dvyhuv/5rssFz3gPzX/+dpVtAPDvXJ9IEDsm+sXypbc5R+unV7Qy5dvyWVfEmq5aL093ZJRzojHZ090jswLIPDMCnvU5ZWHLq5Fdnc3JF8AZJ6JUl25iRFYDQhG1uoHO/k9+AL0UegokfykE/cAUgLT5lSwKhQySZlWQCoAGiBZwXFAZRnc/OED1RoxZlK63FDyg2xMjMw53V19RBcxnEw7+OcqPgnIFEqcWNE6aftPFlPAVCBtEBczbS7cgqSwEwb4wcsotWNNX4Xsm4GmLAyPp6SdFrZM9euXqF84PDwgPRwrVagAoMvB+A5lZKdzU0tKqhVZPX2IoEKvAA6KMtEARy8sLHDumfnA2BCjWewInEdWYAMClTg/kPyChvgTBoSUlpNt76xwTWwI9OhQEgyTXYh5JnAjjAwR8FwfUgoW+QMz6OACq4LlIxUQB5tw3nwbxwbbYbudL1WlY1NyE8pUGHxiAEVpaJKUKKfba31pZ9sTrE//afYfmfvGQjSLP1UpLxhN6WfwI5wiRa3trUeH+0z6ScfqMD72nZNiPmxisYbYFTANBtAhcpEAqiA9FOxmOd9MUZFCFQgzkky3tjXOxst/fQ7ASoiV5I7LUV39/lewEbkEVqSrb8Nu+IPEaiIWJN2F3FFQuwuPnOMRA8Y0AIT7djWhP3vBKiw83pJzj3hGqfN3zwUNCnZ9tYFezsne+XOE3XNjC4C5ubdDtlooS8/a+0DSZbEDeIXnSgjT9jePUu/3myq3bxpViBIcxj6aIUJap0XVZO+3etOQAX2AEyGuuSxJkRVlqf1kIzDmwzg3Tn9UzcBFdpWq8bXPaMmVK1y34+J2Q+OSWLehDoHq0eSXnooHWoAxl7xr61dfDYC82BNJBt7E79nctdJQbWuO2wXq/ZDgERBiRA0MeYH+o1J7BiK7OAxgUQ6AAGNW+wV7ok00W4yTVyjXBEYvou1nHtqGixrIhvnIkjne4S4ddWu14pZDYQh89nJOOo6aH3pFQDQ6089J3Q/xaMF98qkqeiJyXhI9waIDdmXDlhqggi9scr+d8VQ3HM5o22cBTGI3odQDkv/rRJCFuOotJTOE4hBUMimfpSaLCeAg4JLp8hAMAaFoZ4ctsqn6XcBVJhEtsUr5sFofan7ChRDaE7K9uNoC3MvMZEf/ufQw+R7f6GsJMpvwzPEgXOIkcolzSVxLDgGlYJcKkcGwAiFLPgOGcnwCXWKHABqcA+UoQHZqwzbhHMpUBF6Y+Bew0QcEuUGLOnqoHfVQA1TAkBhZyaddfOQMtX07u8xn7FIEIwkZUfr/dTpCeNC74WOBmWrAmZ3Yw9FqvcZFXe3ON3/1lenB74coEKv1y0vu8O63yNQEQYc4T2JTCr9vhkVUZOXC6aCKwgCTIYJAVykn/shdXN4zYDOSe4E3/vSgQp4VLQDKmCojeRMQQb3Qacbmtq6uNiLchapVABUsPKzBkZFlRtYrPVIeGOipkeFk3DAQtTV2y2JNAxUEfzUmHCG9BMSNvNz89R8x0IFo1AAFYjPpvfP0FzTgApWvtTqTMaj4gKLMeJHS9rbRhvtxTnRfvxvkjWKcoeV0VhkWq/RdAWTyZjAQMnACfQDzoeADMGJJfUtQav6i0leE7Sxr125wnaNjo+zT8AuACiAYAG/wWc4BvoQ/6Nvcf2ozES1JvoT10PGgdPTtiSFn2i1oJUgEu6N05Nm5W02y3uKhR9JtWWY1s7NE6joH+iXg4dnA6AC3/XlrHp6upjEYmBZDYEKxl+JUC4I/QO2AoAKGLxub8FLQitI8Ryjr8bGxuTzzz6jmfYDDz4sI6MjDMLwOaRTTHoC57cAU4M4rcQFCyi/vcYqBgYFgor1DIMe86jAtT/xxBOy/8AB56MSkzikm+K4x0WyVZBIZLW80XERZHg6vLdu3JT/9nd/Lz/4wQ9kanpKxDEqNBipSq0CjVVl2sRQxe4lV15++WUmFh973DEqHB3Vkj0GVIhgc9SgtvHzzz9P8+azTzzhNMu14gJST+hm1R5Vj4r333tXgYonAFQgUAVQ4Sp5UCEiNfn0k/OyeOuWPHX2CSZBawiOzFC7VpOb12/IJ+c+oeG3ARXATZhszBfkTR+ocLJPCA5V+umwTEyMB14p+P5HH3woJ06ckMOHDyvYxgSg1Tp+OWtsE6jw2yRxvObs2uC5OFaD+rj09/a5ZwnvYE52YI9nSMsNTR3+HAiIM5Lfycv7770hSwsX5YEHZ2V4fEwSSUhjdUsy1SUYtuqdshuo8HsKycB6o0KjafhUKEtCQY1SaVs+/vA3UosV5cTJk5LtGFZWBWnjGjz7r6Z5AiCfY0MtXP9UYpUdmd4/K3OrYERdlv6+LhkdOy41yTExfu6DV2Rj7YZ8/evfIFAB6afC1hqBij/5F2clN7BfyvVOuX17WS5f+lTGRwdlZfmWbKwtyqPfeIjSPFvFvBTrnfLuuxekI56QB44dlYGRUanAbFzwXNZkfW1bPv30U246oNc/MzMtk5P7gk1j6ygCiwi+SNeunJfz595zQMWQ/PBH/42srtGxQZk5eFDGhrtlY/GS/Ml3npCPL12TK9dvSW8uK/29PTI6OCSdnQBFBqSrd1AynV1SqqI98N4BeF2Tza28VKp1rmOZjqwk4JOQSss6jZuz7PMdABXdXdLb0805lkBFHDq6uoFlNTkT6pC/yxOoQBIZzwqOa9JPmLus2i0001YQ3dYxm9dxT7u6uglUYAwiCW+JZ8wXW8Ui+xIAcGF7R7KZTq638IJi/SIkDEvKqMALczx+DxBhZW2F5wMLwTaZBBViSTIqsJmGRwUYFQZUABQu1FGVKNIND4ckfKdpZLTmAAAgAElEQVTWyaiA9NPa6jI3dGgr1jcF0RUAtjXCPCYUIMcaIFLB5tUBFWAGonofbYPMk0o2odpPWX8bm7gnYDdo8jyRTHEsAEwA6AJGBe6Dnk/nVNUVDhkVaBekn3AfwXTB2mOxAhgVWOfQNhh2499Yo3GvIJ0IuUMABVirbQ3FbxWQSYgBFegDk1kkQOCkCS354xdQ2LVxnnHJGH/9N6AC0+7OtnpUAKhIeYwKS4pZQsr+tPGCMaheT/oycEGrPrUKlgk8F1P40k+QRDOgYnNzQwoeUGFxmIIWcckYUNHzZQIVKqnX9LJ/7pktbrcu3fMP2i9uXwZQoYP0iy2ef8hARQuSoMnuoMJL/7YX0I6qDB2kTbz03ydQ0XqTgmR6O1kwfDkSqNh9u/WZ1+2iJXEtsnL5+4gx0p5R4UvT+D/UmvbmV+QOlRl75ynifuIDCFGDdi+gIkwM668NBOGpXOLbzCg04atFRT6A6//d2nAnoIKygUj2Yj+XSqv8qZkct8BeetnYNJgcbsuVavZbh6ex3/hPBYxtDx2CzAY+hHsI+47O9xZHuwp2F8O3xq1RQIWtrf55bR3xjdANNLBEt/V/Ux+6wUG5HZp4q1mwXZcNdcvjUO0APo9uf2fTmfa1Jq+NMUIZZVfMFSTLyVwIR6QVfnA9dnK05u9g1+/ff/PDYB+4wygzPLwPlJ0yvwBn1hwcw12j9R2Bq1iMwAkS+2iPeUQgPsOer6Mzo/51/jPhLpxeC2DVg0UAn00wGUyyKJCWwjqrLAW/+t/ugxa7QeUgxSJN9Y9QRpDFKXi+AVwYQIC+JksB1f80ydZnRtkubhw78IR9pRVkAdvBGA1+vgqhE75rZuGxREL+y1+Hz0IIVOh5MQYgOY08B02oObEoQGSxDv1A4zDR1nyRmsRr3gDPJu4nxojKcCFGx/U7A3CydBS8QkyJohcAiohJ8X32AYo8wWgBq4cG6iF7BefFOWgHyTGbDMAw3nfHamqd11Aka+CIjX+/yLIZqHDnQ/RthvP3gYovFt/c/9Ufbg/81V/+izaNs0y4Pvj+i8h/EMA3K1mG03+bZBI+DIBH//gaHHKddj/TKdkPb6wN9rsvZqbdulDy6tzkxs9+K6CiJVLe85Z73w1X4sg42k8INZEhXLBivJbddT97ARXevd3lK+K3Lwzw9G93kn6KACog/1TIK1AxeUCKBZhM68JnAQEWEkgFMbFc0wR7o17xgIoGta4NqDBE3ICKJL0XNNlsQAUSAPNztxg0hkCFVmBMOaCihgJ5VjJA0LlBoALsCgAuWDQM6TfpJiaWazUCC1ggp6emg0DUAiwNFjQZZEGcjjeVfkokFKgIvAUc0m9ABdpq8hj4nVEoEdDM3bwpVz2gAkkJMAvAqMD3LCDGAk5TJspJpVkFjwUQ4M3Kyqqsrq6waqMTlZupNM/XNNZce20oW7DHSs8MWBbdgawXgIrFhSUCFZB+ghTV/tn9BCpMfxvtsWob6F0jaaOalbg+rUDiWMBtcHJBuH+QfEJiCKba0EKHxj3615LXOOby0pKM75uUBx96iJX5uBYk9JAsssAHnhuQ07D74QMVxfw624Bxg0oMABW+9BPOAbbB9IH9DEwwcahuKhL9BSm1ASqQtPOcAwRAxd//v38nf/ZnfxYAFdxc4P5WazSHxSSgwatuMjgvSUNefull3sfHTPqpBaiw+y4xVJIjEd2Qf/zFP0pXZ5bST0zgpbT6woAKMxpDEPfeu+9KrF6XJ86cYUWJAiC6P8J1AKi4cO4TWbh1U779xFnp6Q2BCgsKIW0F6afT3/IYFUxeCu/hW2+9JUcPgVExrtelBjAEKgBGmPQTrhvf/+C99ykJdfzYMfZ5a6LNxmXrhupewId7+e4XWcWD7YWTfkJg29fTq8ZzpKWH66k/pjlG62Wpo8K/gQBbZHtjVT5673XZWJuXUw8fluHRcalVOyTTMSCNRJr92SBQEaP8U7uXJi3DUal7CkWTAObOz12Uzy5+JAcPz8jI8H5JJXtZba6mvNE9ACN2SJ1B+una5x9KslGUmdnDMr+yLWtrV6Wvp0vGxo5LPdHDSriPP3hVNtduyCPf+IZ09U1JvZGV/OaK/Oq5H8u//FdPSa5vWoq1DllcnJcb16/I9L4x2dpckutXP5dvPvKA9PZ2y/rOttzeqsnFz29Jb2dOHjh+RLp7+6Ucg8k8KtLKcnt5XT7++BPp6c7J1s6mHD48K9NTk7qSuUR08xgAs21bPj3/vizMXZXp6RlJd/TKD3/036VYLMj4xJAcOnpEcpmYrMx9Kv/Dv/yOXF9ak5WNTRno65Gh/j4Z6OuXjo5ukXiH1GNp2dopy04eMgVJyXV10zQbjAqAgVhDwLKxBDiS4jQzj8UIPsCTCP8bUIE52DayBlSgag7a/qgMBFChAHopkH7CPNcMVOgmydYmAqNOehHzBOZpzLcYj0z+o0KejMYGGRXYUOP9PBgVmY4QqOD4i3FTiAQ+XlvbCojj+ytrq7s8KrCxBqMCYA3mvStXLsvqMhgVKv2EfoCZNubF7q6sZBIp2Xbsgnq1LKury9xEom1gf6j0U+j/QKDBeUxgjoV8EddlJ99IRgVltFRyCd4eAB2igAqsJWCtAMgBmIBz6lptlX8uoRSLM0EF6ScAUOhXGMAbUKFsCIsjQqACgIgBFWqKjXbtAVTE4B+lEpT4H+0HOKBABWI1PLehobYlTCwpxEjbPdi2vutTDgNSyGvVZXsLINmWdHVlKVlpcaYBFTYvB8mBRILtuFugQosgwJBBQYp6VPjSTxsw025hVLDy1AMq+vv7ZLz7wJfIqPhnAlR4CbWmPdUXASv+UIEKwyO8BD6TkS3vc/vppEVaVzIk+9yi0LzjdWte6+7ud8qosN2wq8a2mLH1GvQ5bikmsL1dMA6ajccDxmeTT4VKj7R77QLv3Jes6GVXm9oYj7fbKQfvMeYMDc91fsKbukdrH9OEFc+77qs/Zj1ZKcaf7hpt2PgJ+GigwkAAGy4tfgYuYmeVvJPIMa15O2e7amqt93cgUCDzYykTAyqU8U5pZLzl2P44rskEWbvDRL/+JgQqgmGuLXV5F//7flzdDqywZGxYPBT6L1jFt/kE4AT+PlbPGY4tVOzbcbjqOMknK4ph1T8St65Qibsh7K2d54Tp/BuTAfs97PsULFC+NxO75pvBAgHESCoPhb+TBZJMsepeE+0Kffn7dusTlU7SY6L/A5+BYAA7SS0U7jgQIvA7IGihLB99TgHSK2NBxx7GfdhWJLcRk1js5j+RAWjh5K3QVvWOSKhktWPLhLGQygSZAbiaSWtsoGNKny2VQEq4pDv82pStAZDCWLlmDE8nSTIRVOqS99H8p+gxoiwJk4tDEahJSNk4wJ5bizdTBGXwG9wDemIkE/I3/0f4zH/vLwD2qYk2cicoqAN7F2xdKmxAKokMnXC84z30DZ5Bi3Oxl0ef4xhm4K3FnQpGYOxYLGOgjcZqVYIUvB53vzB+KW1c88AgsGQxlpyHGKYZky8jZuPAj7aTmSsbMwN5vRYFZawo0fJRfuFYvaFMLaiK3GdURPXs/fe/sj3wH//DH+/R9t0hhaKjLT9pSnS3M3E2lALTv/d5kwpRCD5wIfNP0xRs49ytCfiwPUGsGiRquFS1ucaINgXf3At4CD8LFl0vSNaqhz2yOnczWoKfu47wA04XDLU/TAuos+tLre2KrG8JKIrNwUUYmOHa6YkAql4V5pwVKdKjIopR0QxUGJXQ3+CmaJgIZgOqBABUAMyoMtmNYQGPBgMq8KeBHV29PZLMpNjtpPqVypTfUKBijtJPBlQIFxf1qICERZUa7ApU4PdlLHrQfi4WWZluVQVc0N2ijo0NEgpIIgCowGJlCWJbUBShD5MI6EetHoyTLorf+kCFeVRg025AhfW9BZKo2L9544ZccdJPYxMTDCCQnMe1GN0S58aCzKoMUFzTKSZVcBws6mgjkiZrq6uU2sCYha+DLYL+sMFnmsTQgBSBCRI5YE3U6hVW+iKptjC/RF+BAwdmKU80MTnGJBCuC8kv/I/EC14dnR1SLhZdJK7BGbQcKTQEDc8YgqAaKyZQTb6+tkZ5JQAVoFMyMU96qFZmgnGxb2pKHn74EYIAYM4Q5EAlhQs80D9oAwNiF0DjesiIyG+oRwWNzyFBlmGfoEr52Z/9nNrhMLIGowJ9GUg/AagoFijNAl14VMsbowJJOxasuzqPW9dvyt+TUfF9md4/jfJ6jjsEmAgENZBT346A+eSqi15+6SVeJ6Sf+gcH+B2rXrHxptcFfUyVLPvFCy9IVy4n337q2xoANgEVeHa1ryHB9eH77+HBkTOPn3F0Yf5TZxoHVJw/d04WbtyUp86eZaJYCac4lW6wYBZ+4fwFmmkbo6KKz8A6KZYcUHE4kH7ihi0eC4AKYybhWAAqPvrwI5memqLxMTwvyLAKgvpwhNomzN6xjZT/7ERNuf8UQEXrMY2WbfA9pJ8wDnWT0AxU2FzItqPix91TbkRqddlZW5V333xdNgu35Gtff1iGhvZLqYwEeD/HGsEK7oGi0gH4XGneBHWp7+WSjxg7+W05d/5tqdXLcvz4g5LNDUo8jgqjZqBC95rehhNSQtg4Jxty/eI5SdTzMn3gkCyugA11Rfp6u2V84oTUYt1SKZcJVGysg1Hxdcn2TkpDcrK9viy/fuG/yr/6109Jrnda8pW03Lp1Qxbmb8rBmUmynj7/9GN55OETlI4r12py6eaarK7kZbivX44dOiiZzpyUJcWxDfB0Yf62nD//qQwO9stOflNmZw/IATx7toENBrkb6yKycntRPj3/gezsrMrkPshSpeXHP36a8/bU9KiM75uQRjUvmdiOHD+0XxqprOT6+6SvJ0cPEjAESqWGlCtxKVbjki9WBYpykDdSoALr2TaBUawhnRlUfWFNSLJ6P5fDs9VQKbmePsoLkVkGc24fqIDfEYH9FOdJ0N8R62BNwdpiHhUGVGCTCJo8NmOc65zBINe5hNL18QKLAtJGLABwXh44N16bjvXX1d1NRkUnZOIco0KHkQIV5lEBoAJrCo6zur7G78Jo29ZuAgue9NPly5dk/fYKGRVd2SxHWAmbMLQLHg6JJOX/AO7UqmVZW79NpiHmIBzXNJmtLhrj24AKbIQBVABsQOKjUq1xfkyl4aOQYH/4jAq0kUCHx6hQTewE+wfMRqypCsAbA8OYXwoOZTygAowKZbp0OckKPT7XOLdGglGB4oFr164FgEO5UpLNzfVAPtHiEZN+gkeFJVUQJwGoUOknrbaMAir4BLuKSGM5cK1inIMEAhIGNQIVYE7muiB9pSAQnn8rLPCBCnuuAFQgvrgbRoUaw8PgvNwEVCQTAJBQ6LAh+cJOk/STghSqvw1GhQIVM5QtRMxhBQqIKZAIaU0O2hztz9VRa4S93zSjtgvv/VJ02164aRLTsW0J/L+3P2eEVM+uAq7w102ysN5BoyQmor4f2Qd7ABsurcefNq867fdQ7ZKfe/d9m7p8r/9/262WNtwxi7yKdUuY81YG53OJaquCb22430/m/+K+E7Wj9KvQ/cNF9lO7sceD7wYq9BlvbmTzvVcZGH1u9bkOV8LddyWKvaDHiGpYuysPTc79caPzmMUnbc7fKsWD7zcxTLQNFoO3G1cqB6XgrfUxYzN4CHqecvwtmsn0AUx6Ia2kpszWTt/TIRz9nmm7a5tfZNOuTfQE4vlD8EDlV/F+OzDEEv7Wt25cev3DVnvjkUlwaPyDcegKFfxCTf++42joJySLsZfg9aI9qC5ngl/32SpB5edDXN0p15WwNjXwaAwkTtXcG/serJ1opoIU2geUwWXlur7P++MUD9D+oLA1MD1WwMGQF7uPYE2iWM4q/pVlqBI92NvTs8BJQXNPBW8IJy9EtlFN+1UT1soAbJ7lHKPASe+EzwDao3KsKUiiemOO+xVnBJ11SXbkOhBb0BPCsd0po4RYpVyRTKcWLOC+afJfnx/6LQbeEQp64AXQBbGhMi2Uect4r+E8EG3/68AG62syE9z1UpYJxXtgeoCV4GSfkVcAK5qgkTF9HFNE8wNaROC3zf6+O3mIOCLJ46GvUahh+1nEaD/+P5Wpitf/9H0tqOH5IZPlfCfwnu354skY4ykrujQpZfPtaPXRUCDGe7nr4b4IygrwygCbhPe+LmB5mGm3iiI7tgjBCmWhIOYycAGHMz8N/RPMXQWSEPPbftbAFZXPcs9bo+6uA3ku9Tqxecv8UJiDc3sYBUDuSz+1m1/vv/cV74H/+Jd/tPsKIpMcuom5N6ACgUS75LjpRYaLnC14FlxHB71fBlDRSmG1NJJ1x90CFf8fe+/ZJdl1XQnuMBmREeltZZk0ZWEIgEYkq4ACQAAi2RI1Us+s+TBamhFJtVbP9D/R/IT5oJnpbq2WIeVGFGikbhEADQhDolAFoLzPLF/pMyPDz9r73PPei8iIRJUcB7MqsHIhKyPivfvuu+/ec88+e+9k99l3jBnyrwRUPLA5dreB2h2oUKDjcEUU8DwIULGV8KhgNd46NkKihawKmmknE/RJoCLXyySw0ZgVGNXMVFsa2c2GNr5M6HBjz02pySU1JP3Uk7dEC5PNTEqwopGV7jcWFlCvxh4VWoAB7J2exeDwEKqBzqeKBFakygwrre+oaoUJZcUnRjl17dLSZhmVeg179u0z4KFStWQzWSKBFiiD46gaxJ4fJoxlpl2toEQzbVZmNBqSOFIg2JNFsa+ozbYHAp6gokk1JXYuX7io93dP7UG+UMCevXtQ6Ke5rgUiLtXEfmYfccPPpArPT1NmqzKwwPX+3XvyvSDQYmCCsQ5cksH1LbUoh2onLsg9+R70MLBoNgQm0Ez7xvwNzM7uxxiNridHQeCJQEl/vwEVDDL4ooQF5ZI82eHBkAMh3BBxGFD+hEAA5TvIdNmgSecGk3zGqODmgQm/O3duY/eevfj0Zz4tHwleK6+dpp4KYoKnRP/gYKTLSfCBJxFAVF5TRbIYFemMKjqt8qaG7373ewJmCFTMHdgfUT0ZxKeyafVnmSDKyrKq5ZV8ZtVTeLQoxMTdDitw//rP/wq/941vYHpmL9K5jII63hN5mbh0mMzcmcQmkEE5sxTeeOMNBfXPHj+GsclRozkTgNFYsw2EnlfKmtTqGsOUfhoZHMLLL70cADarbmHiq5miBJBtqLbKNZw68b4S45SJMl1TAyr0bLJ9zQbOfPQhbs7P46UXXgSlu+qooxY8LHjfyKg4c+YMjh07hvHRUaNvpxnoNtSed95+G48dPoK9eyi9Axk58tl67bXXIkaFzwUcs6dOnZKs2r49ezE+OqYqYQ+W28GJllm4beP6ccWj0Zr2j5yy2yuvvJLOE50tK0qzKdBrZJgG4ZroWtYKP5b6jpqwrmnrAWy9rnH2xo/+HlvlFbz8qy+JNt5sZFDsHUYqVZCsXQvzMRTksdpewa6NFP3E/ch5nVVWady6cR6XL3+Iudl92LNnTn4Y2Z4+1JvlKBnRClQwQKbOKzc0Ncxf+wj1+gZmZx7HvXtl3L17DmNjg9g7/TS2qjRzruLMqbeweP8Kjh49hvzAbjRSfVhduoM3/uu38N/9+q+iOLAP61tpXLxyEUuLd3D44Czu376DMx99gM9+7jF893t/jaNHj2NzixVdBUyOT2H/3EFkegqoIaNxubS0guvX5nH39l30ZGmQnMb+A9Nin6kHbDceNri8DbYRuHb9Cq5ePY9arYTp6RmUNpv49rf/GrsmxzE9vQtjY6Po78tjuD+PyYlBjIyPoVDMobK1gjt3lpHpGUSudwR19KLSzKBcpV4yNx15eTdwU7a+vqFNJMdzb56yT8bSMqCCIBaBlk0MDY1geHhE86vAAs7v8isiQEG/o6x+p/E2E9wpcENZErOlr4/rgQHtbibNZ0hzDTdflAxoNlWRn01nkQHB+hTIdqOnB+dYbqQ51/P4nKvWShsg+MgEP4EUjj0l85eXLPBJp3RNDooTqGAbyFwwoKIhc3DKLRGwEm2+mZZUFosJLl08j+XFu5gYH0F/H2WDmihzjms00UegIpvTmtlfLKgo4v7SPfTkzNtoiMUK8tkwE04ygbhGrK2u6zy+DhGQqdKjolbT/TCZP1sLKZ3ETT3BDzeJpEeFfKNYJKE5F7h79w5u376jBDn7qF1uihtJ9nlPNqfEOfvg5s0bAqbYTk8Wad3ftBiJ12dABaWfzKNC96tGT5NlMQ24jrpMhhcVbJXKATwwRoV5XRijwjbNxlpNJss6Jej9bzZ/caPO/6ewukLZzvWIUeFVfp5UU4zC0CBssPl9Z1SwHUlQwFkbDlR5nGGSZDTtNkYFf9h3TGK4R4XJnFkSJPl/JjdGRoYwNTC7I1CRvOaHASg67gg6rBU76U53ir67bxF2WIg+bjFrO9G/PFDh3IKQIG45/ycHqNB66d3OZmt5jFkZ0Xsf0//J/k5KT2lf2OW2dh03XVgN3T7vKVOdK3kfdpBsVLIzJD0NoHSVoc6N7QZUWNyyfZS3ai7E7+ujHb4QMzw6PWAhkEnEd4whBZz6oRO/WP369pcVApkMJ1+MT82A1yT7onaFY6loisCGKvlN7tXZGN3AJA2duGrS5t+kHFl7swJrxI9n+6Kk+XEr6JD8+scBf9H7vGwxAbhfCMAI9fnDvG3HjPvdyLYGAHBNjQCTkJSOri/R5y3yoIn7K+PhUGQUgzGeL/GcgoFmjCN5bAESCQUHySkxoc9CwyBrxCbaftf25aqg137azJHtmTDZLQc/HGiS/KQS88Y2cGSFx+A6TdCCyX4VJFZsT22v9vyTAkk7lw1srZ3uecG4g8+BKvlZGFe1JDv3aZJj4nZRAIrtAwkoeTxie4i6Sm0Z07n3gbMPvD22jgb2Qpi3KKPNIjQDPAwU0vobxkAEMuhvlB8ObBHJcbJ4jvtrk0KSvBRlkkIfiMGj+xOPF7PhsDFr0lwOfpo/i8Ug23OBcY7DCkh4//06/+gP477+3X+PCKDw58/HlO+1lP/g92W0bVJMKmogo4L9HuaKiNXQDOM68UApByEmg/ny8fvOPqZqB58H94hwLzQ3VneJJj+cP1tuAM44MTY0jxlEHlOFR878beQJ4kCRyXDpvKFY1AtGDOALLCuCJ4+knzrO+4/++Anuge6Mis4J7JYcUBQc2GdjDL2tQ7YRGgIo0IZOx0BFTLVIwBiJg/6ygQpvSrLSIU5M/qsyKj6BQMXE9MEWbwZPlinx0kuZEUsg8e916no7UEEl80JBi7uh5pbsqNVopt2PrIAKQ7/JqGBgUN4MQEWlKi1pVrRKrwcp7Nk3g+HREVTSlpRXgoPGwawwZdVMMI+yAN5+7HNpjXUDKqryiejpNdOlJuU3KBgfggsDUqzK0o+R6WEQZhIeqpINhkkEKvhixb68I6QpGUIRVaqWMTI2jIWr13Hp/EUlbaYCULF3eh+KA61ABa+fVY2e3GVVK1/8W7IikUFPabOEO3fuCLBgIpUa5FFgxjx/UPzlrVE9TmCW1LOmi8l45eaNW7hxfR7T07OY3LULw6PUz7dKDlbpJitP+XsLUMEkZwhmKIvlyQ9KhbH9THzIuHt9HaWNjSD9RNMtmkhXcPPmLbFKnvnMMzhw8KDazwCN37VEtGmnU/rJgwC2gYs/E1/VrVWxJxrVuqommEhT4Fip4dVXv6v74YwK0Ss5FhioZbNKDFY2S1hbXjIzbTJ0ZLjdREoVXwwgM7h+7Tr+n7/4K/y7r38d+wRU0IzbJEBcL94Cb5q5M6Djewxk0wIq+Jnnnj+GsfERJRlJV46AClXvkMHRVEUQGQwEKihD86svv2JUZZBCXUO5yqRj3QyzGwRjGnj/xPtINWqSfqIMip69BFBBC+YzZFQsLOClF17AwGA/ak1CFQzQLQilmTb9AI4dParzMnhKAhVvv/U2jlDiaa8BFU6h5bVR4onST55MI/hz8tRJzM3OYe+ePchlspicmIxYFTstuckk1Mdt4pLP5YN8ttN5PxaoCIkPrVoEItMZSaNJW1/iYK3Bu8zRwvxnX4krl3RfWPm9vITv/+A7yGSr+MpXXkQ23YNsuoj+4jjqjXQwcQ+QhINYSsSrNC26DA/G7Q/cpPdgq3QfZz58C9meOvbPHcbg8C400as7Hb+SiQnCakCDXjjpCq5f+wi1xiZmZ57A/XtV3Ll9BmPjMVDB9vP4BCqOHX0Wub4p1FDEyrIBFb/1tS+jv38vVjdTuHD5PNbX7+PxI4fw4cnTuHTxHJ47/gzmF86rrXfvLmNsfC8OHXocu6ZmkMkW5ZVRJVCxuIwT772PYm8vlpcWMTExgsNHDMSMNsCSAjHJP15eeauECxfPYeHGZaTSNczMzKBUquKtN3+Oxw4fxujoIEZGBjE2OoSRoQEUi5Ra21SC/dKlj1AsjuHQ459DtncU9VQelVoa5WpNz1iOQEV/v+Z9JvndV4ZzkoAKMhYSQIUl/Efk6cB1gt/h2Ob3OG9x8yn/CQH3ZZvrkFGRABPNxaIliTnfJc20xUxq1lFrGAtmq1JBT7oHmUZKgE6hL4f79yj91AxARUbJdB5rtbQhgJFzp4oF8lYBR2Ye5zx+xqWfOG7pUcFXsdiPpeVljWUyH/g9rjm8bjJQBFRUK7q/y0t3MT46LDCIXj1UsuNcQTNt0v3pX0OghPPYveV7OganS0pkZcP6zDUaaZMuomwV+4DXTTCAzx/ZOGSBGlBhlft8n+btXP9kZBikO7j28N8EKqjjTF8XrpW3b9/GyMiIYhJnclhy3+IJ8wYxSUX+uwWoCGsdP+uyXsViodWjIvhiEKig/BHXIDfTVhzCOIZAMwGqUFVJ7yl+LpZ+MgNM//H5rtM85vGNzTlMFnE+IOiw3iL9lJSrcADENtpWpZwEKtoZFd5uByr4Hd4bA9KqkZk2gQoyKiYRZZkAACAASURBVPheEqhwkMKLKPj/3t4emWlP9c91BSrsuuOr/jigolOatmXX8QioCJ1pgPfDvR7u890YB1Fs3DGn3SXR3g1oSPgmc+qwov6EfFSSAKA1tFNtcNgDR+8nR0y8hrf3VVd2S5e2OoO1/TiWkm0w/Ewu09HvUWuSD0LwhEjOC61FCNvP0uled/OoUOV7hy9E+dy29wSEdLnuTuNAMZsKPnwYOrrQfUS2Az2KrzyB6syn6DAB/nGJHCZqBVpY5XjXgpnw/UgMwo2Uuwx9bXkT+03fC3WOSdvjxc7X2v5dVqzHALFVa/Pu+DXEn7fjO1ChorvAqLfKbnsx+evzvydPky1J3kauj2KNhw8k+81ljT2JGyEGqva3+cUT3ZH/nzwSuBONDYyT1ek8ja6VkjwJPp1UE7hWBTAkmczmPZX8E/2vgrQw4wiXFOo2ogygiFlfNiRdwskMnh2g13Ej4KBqv8sDzgySPUluHl7GJNV1kE0hiaSEwXKosNc9DOuuMyQZy0iZICS13dzak+TMtUhu2C8qKjizoje1KbSLeQ2PIy12DEWOYh20jkVL2BMiDNX9LJwjyBN8wzoBFSbnZMUllnQPzJ9Mq/TTb3+zGvlwSGpJbDFTBfD4h99lwaWv7yaHZewW/90koNzwu7VgOfnMSNEDUDzI/TaLZjMqtHRmQ5h2tF+zH7/Pfn4HMPQ8hfe9y5P329ofQNdov2bgk6a28J6P8Wi+88lV4KGN9EdARfe5/9E7n9AeaAUqulXXJ+GCDpGHKjU78yBspm3vnI8BKpyr2i6nFB3mlwBUqOKmPeR6BFR0ln7amVExOXNIm3NVdobNrQIfJl4INijBa4GbsxSYLGAQzmpBARBbZD0QNa9J5qNvoA/ZfNB9rtVUwU1GBZMaYlSUKy1ABReAyak9qvwnUOE6i1xiHahQ4BgFaXbvfaPNBY2SC1vVCsYmxtFHc2EubDVjVNDdlnU+TK57MOSLV6YnDf4QZGGyR4t6vS5GBV8EKniNTOZ4AoB/J1AxOj4SARW5TA67d+9Bb7EPBCoGBvv0rHkiy4EKtoHtZpKG7dY55ZVhfiD0C+EixyDITULX19cxOTkZ/BgsMPFKlEyoFpJeo6o2GQRksLayhutXr2N8fEJAxcjokCpSGCxSvoRJOjIT+KJfBgECM7Kir4hVrCjRkTWzKraZbeVYYQKG10U2BSVHvDpjq0xWypaMTdkXDlQwGalETrhnzFIsrS5rXHhQMzg0pCQTk5PlzRXUKmZozQ0Iq2wjoOJvX0VvoRCZabcAFZmMGBWVzU0BFWRU0AxcQAVZEZo2qHlpjIoIqJjei3Teqls8+ajgUonIKtNdYeIkCJTGj370owioIFjF546+IqI011wuKiWaOvUxyQz5wQ9+gKH+QXzly18OiSBIv3WrWgJSfG4YGJPZ08DJEyeBejUwKrYDFWJUBKDi5RcJVAx0BirOnMHRDkAFxzoZFYcOHoqACt9AEKg4cOCAksI+H7AS6NQHpzC9bxq7p6Z0PRNj4xpDMrnviJjbArHTe502fg4g7gRUtB+z/bPJfyeDZq/e8w07ZxHOMfRLYfV0Z6DCQNrk3OjH17NCUKqRweLiPXzr2/8RuyaG8PIrL4hinsvm0ZMbRgNkBIVXkLVQ1ZeozkmgIhmos4qHdfUl3L55AZcvn8H+A3OY2j3NcB3NFCvc4+8mr1lVhw5UXP8QtXrJgIq7Fdy6dRoTkyPYs/dTMsgmhf3ch+9g8f5VPHvsGLLFXag2C1heui2g4t9+7csYGJjG0noD5y6e4YyMmem9+MkbP8X9+3ewf/8EnnxiFqfPXMHly9dx5MjTOHzkSQwOThijopnC+lYJa6sb+OlP3sTMvn24cYMA6h48+eRjqtSONtGhypGAIv9IGbwLF89gaekWevtS2DU1iXyugI31CiYnJjAyPCQZK8rNrK8uorS5hoWFebz55o+wa3IXnnrmCxgc3gtk+tBIE6hoolTmelQXS4vjl+sB51cHKpQobwMqNN8TqBgYFqOCIIXP2z6/c83iJkqGyuWq5klOADw2E/xMfPMx4bzOtYQJASawHaio1huoUMKQ7EMmhQNQ0VvsweL9RQEVNMHm3E5pP77WKLuHVqCCxyVQocRBOiWgxD0qIqCi0IellRXN25TH47xPoIJm0dlMD3rz9FMq49KFs1ghUDE2jP5iXqBvrWEbVwIVlHPk+kzD73JlC4uri1bZ12hikCbVKUpJBQZdmsUDNazThJwbczFECsikCFRQjisGKhy8dqBCAEobUEF/LLJXCAYRpLh161YAKiiJZAkEARXB6JpAMpMeDlTcunVToAIZFb42MdPC9Zf3jG0jO4Cf4VrBtYk/TJ6wXW6mHSXrucY0yAgsRW3lcfgdrv1WpbkdqOg2R2otCvOnMyoIXq4sr7UwKjjekvORJ6vigpPuHhU7ARWNhkl85vPmURFLP61is7QejONbGRXsi95CWkDFrr4DktrqJP1kCg2JfcwO64dPm+1z/L8eUNFtM7lDgv8hmRYPvV3tenxjzD8cgfxfHqjo2oM7ABXua6Fx4ibzES02gP6+pD58B7bI8CS//rBARbfkdZJRkVj6O7Y0kiFLVKzHMkDdpMd4qM5m2l1ZIUoXbIcqBA50bJkDOh2RwCALFVBHv5eqkk58PqQoOsZ6gXXsc5azJFg9z8Mxro7Gcjik+0d4URHXIpfleRCggpfp4M/2RK11ggqiFfOZZj8TqTpPSEDbMbo/Nw/yHtdxxh58JWX7uhX2iHURGAo6f1sy1mVulAR2aaaIVaBvRHfYZCZN7kYJ5nBdXq3uaxIT0L7uqppcpsNuBJ2K5HHNU4Byi7GCAP/WOsenUWswYW/7dm8O7xnbo0IhqTDFiW4lj0FfjazGrYAOXUbMotmJUWGftPyW+bbQX4BFEMbg5HFNkpkFlvQtY84ilgByVgPjBib42U+KXYLRtsk32V6dCXl5Zun74XOh/QJ9WIhSrUb+lg6sKUrxokCCbTSGJtuCZs+SSTTpLfOwsHvooJYbSGsmaJFoC8XKQQJOz3cTimuVF5HHTFJaLpqhokIs9pFyHtz3M2bLZluknwhU8Lp03YEFonZwPxTiFl6XTK/VRywqsYI8A3voF2pxACVQTUq4dcz4I+YyZ9ZXxtbRuNF9sFjP92IOLvkzagUf8ZhyWTzzw7B+iucBY2/wvBEzIszJbJsXq7oklwOGNn9Z2/V9eZXzWHgEVDz02vzoC/+f7wEDKrYn4K3h2wMM/eVhqviDbnZrRzwgUGGzj321hUr5SwIqxG9PXkk3oKJj1z3cWIjO8zEeFQ9zLzq2oBs45d0eAvQoSPqnSz9NzR1R0oWTr5Jx7FRR7NIw6SeVW+u96lYlwagw+QcHKlIpo/cxHugbLCJDKZ1QLUG9blaaUut+YX5eQAWTq8W+fjSDQTbNaMcnJ1ANHhXOqGA1OhcEJt6SKLkHVx5IlbcqKFUrGB4ZweDIsC3sDC7JqEgAFbxOZyewfZR+yuQSQEXw1dhYY4IprcWdC5RXI3owLCPyidFtQEWhr1/+DAND/UpQSYc0sALo0cAEFvuMshF8j0kv9ptJU1BP3WSHPGhkEERmBTW4CTRwUefnpKGaYFSQmVLPWBBI2RQGVvdu31V17OjYiAyXMz2mm8nErGSlgvQT74W00UMySOcPoAWvwfud40QSTiGxRzbFFuWytFBbkErpi8tXrmJ8fBxPPfM0Dhw8oPNZkGda1gySVtdp7LsYPQXUWSfTg9UqldKqqK7UA6X0k4AK+ZVUxahgAPX888/j4KFDxqRwRkUmbfrwAahgEk4lbRmGq1YN1ATBmEyQfvpL/P43vo5903uR6sKoUHDeYEDK8J+V1hn8+Mc/joCK0fFh0VsJVDDCIQsk2qiQqcOqp0YT3//e91HsLeCrX/mKJSppMFzewlZ5E80AVPDYBCpOvU+gwqWfmMjlOHLpJ0h+5ayknxbw8osv6t5W6R/DahIl55qSJKOZNhkVlGpShR+T5NT3rVTw9ttv4+D+A9i3d58lAkLv8NpmZ2f145szAionT50So4Lm29LqbQK7d+/eJqXmAWIU+nZIQvkG5mGACv+sB4PJTVDXDWpohM8VnYAKXjur5Pk8KiHYNoc7QOH/t6A/waqoN9Gs5/Q83r5zHa/+7bcxtXsEX/ji0yj0sgp5CD09o8aQICzCIFY6/8FUt+kU9rYFQfJNfMa5iVrDu+/+FINDRRw4sB99fUOoNQbCMW1BjvfNvJOsMqwhm9rC/Pxp1GpbAiru3S3jxs3T2DU1iqndT6KGPm0Yzn74NpbuX8WxZ48hU5gUULG0eAs/ElDxFQwOzODeSgVnz3+EgYEe9BXyePftX2B9dRl79g5ifGIAP3z9p5jedwAHDjyBuf1HUOxjAtyAirVSCYv3l/Duu7/A+MgItrY2sXtqAk88+Zg8EQTYiKseJB2C6fCN69dxbf4S6vUS+gayGBoewOjIKEaGJ1Es0FiaJtfruHDhHC5dPI3HHzuCt372Y80Xn/nsMUxM0m+jF5ncIBrpHMo1M8wubxEkoHSPMSp8PpMsHzX624AKjjW+N9A/1AJUsOdjRgWBCmNNcA7n53ldBPXpJUDzY74XV6zbRlAbNDRQIfOQYEWthhwZFUiLkdBbzAl44JijXwYZJ5Sq4mt9i0AF/x4zKni8xcX7mr85n29sbsijgud2oKLQW8Ti0rLGDYEX2zjWTBYJaTEuapUyLp4/i+VlY1QM9BGoYPLIkjaF3ry8Kbg+DwwMSsJucXXJ5B7qdXks9cj4PXgqkVFRbwjkVkUnzbSL1ifccMqjon8gAhJM+mlJYDrXvRioWNZnCFYT5CID5PbtW7h16zYoxVgUo8I3rxZPsS8IVOj/ApPScKBicNC8oDSvwBgobGOhkNf9IVAxPz+v9Z+FGUxqLLUBFX5fOYkSRHLJAa7tzjq1DXZc7efzic9n7eGg5rdI4sOkn/izsrwuoIL+Hj098aY9Oe86sOrtehDpJ5M2sCSCGVyaRwjZjCb9lFe/d/Ko4HcE2GRSAipGRgYwWTz8CKh4uF3Gg396pyRpygoy/uVeH+NR0enEXdrTNaHLPGa4xo5AhQ32B7tEq9sL29b4Ow/dR12ZBZ3a0SrB1amhmpkCMyT2S4kTsEmgotuFdoUX2o0wwgHsPA8DVMTJ0Y63NRQUBH1lW7+Thw9do1vQof+8pNJ70IFZr5JWsi8Rw3kbxPQISUGxmJlol8Ftt4HWuQdVWNT2VsiGBBDGE5wGWthcHcaSj6kO15W8Vk+itreADAgW/jGZ6wlfKzILSea26+a9diaiji+5LGMHcM13KSj1hdayNOqSDGxtL//lAISvU55Y53uM7VXwaK7DxlQh6BD8KqJkLN8PMlVsN9dcB5wskVzX2kEAgDGW/AXIMK9WIhYxz6+1Wsl4S2h7Ql4eEZQskj8YpaWNDblJ9YZsrG7Q3q8uL5XAzdQXUWJez1wsvWgyPcETJ/Q9k+9xsUNgAZBREdZkL9yjbKgS7ZRKDECGch6BBSGGtFQl6qjWq5LmVByj5Dh9P61f3TPCzbbVB/K/8PWdwIqBFearYFLLKrpgcZ6KDF36KU7Ka58igMYYFVaYaCzgzk9KbPZOCWc3tGZbWazwR38Y9/b//PsmTcUiNvl0hQNKiolJe0lmUVY7vlfKvYhZY0ARAUm2370nDLgzoCO5n1EcQ2NyxonVwGAOviLMHzngoNkt8W8D5AwM8bnB9m42Xv09L0q0q7OcmiS+QnGl+YGG/ZpiJLbZpJ94bv7fJT2b6QAAqj8eMSq6rV2P/v4J7oH//T98eQegolOQYUmJ1pcttTbnttMnHt6joh3lNOHMZEXULwuoSF510IRLzr6hWSb99E8cFP8/Bip2zR42X4AABHiQxQnYGRWUZ2Aio0rpJMo3rK1qAS4UrVqQVYjpTI99plpH/1AfeghyBAotpZ+4mBOouH7tGmpMbgwOgMlpVhSze8momJicRI0kDq8mpGyITElZYE4EPshCJarzbRFqoLxVRbVhslPDY6O2QBNgIaLPBYufqZR1PCYs9DRxUaGZdmBUSIYpGHeTUSFjSYIDeUtaRJTCVBor62vYtWtCCeGLZ88jl+mR9FOhrw/7Zui3Yckh05U0VoaSZGSX5LNmgCyTWZpMGxjDwI2Ai3TPg2Ynk2l8b3FxUcn1ja1NFBjwBBZGLh2YK6wHp65rJq0qce5V6lUm/4B8b6+SfMaOaIpRwaRLEqgw3VCrtOGXeH4LiK2Shm2gPBQDEyZg2GYacPPHki5QEMH7T8mhsbEJHH7sMGbnZjA1tTsKDBRoBT32e/fuhiS8VSPQYFv1WLWSaMaS72I8XKtjZXVNprc/++mbYt4899xzmNu/X74bumYGahlKrZj00+bKspnIcuMepJ9MOpISPxmZoP/Vt/8Sv/e7/wsOHNzPovhgGGdyZZ5IkvSTRjuDRso7QUAF/y6PiomRCKhgwElwxasBadDtZp3f++530V/swysvvxKScVmxcrYqm6g3K8HXIoOtcj14VFTxpRdflPQTg79aLVDFWUnSbODs6Y8ijwpKP1FKq0F5J1XpN3FjfkFAxdEvfhGT4xM2tmplSQaJUfHOO9g/O4dpSjzVG6pW4tz+05/+FPv375f0k2uBstr5w48+1OfJ7OFz5ZtrjiMCTHwlK8OiZyUK9kxf159hr0T2RKYHjT5TJxN5/A7vSVJqJAlUdE14dNogs7rGiYicT5BSdfTwcPAzSZTw2T7cxrZvwpIghf0ONGusFjIAYv7aBbz++g8wPTOOZz59BD25PuTyo8j1FAEQzOI93kQuZ7qnSHEuCpvTlk1vCikOSspRpaq4ceMKLl44jSNH9ovNguw46q7pGtYnyXtpc0+vFHr0bOLOnYvkkmF632O4c2sL1+c/xN7pXZiYPIJmekD9evrUz7CydB1Hjx1FtmCMivv3bwio+B9/69dRKOzG3aUtnD5zClNTIyhtrOH0h2dw7/YtHDwyhVy+gV/84kMcPvIUZmcPY2b2EAqFYTRTPRGj4vRHZ7GxvilW3eBgH3bvnsDMzD4lmk1ai2AgDRjZkXUZ9t65eRPVSgmDw3kMDvViZHQYuZ4CGrWMpKQoQ0Og4saNa1hZvodqeRONRhVPPfM5zB54CvUGk9IFpLJFAXgV+sXUqyhv1jT/McHPeSwJVJCh5R4SnJs5//I+c5PV3z8kqSRnlsXVgNwwpsUa5DxZKgXpp1QGy0vL6MllBOrz/iQZFWaESPPlhiSpyJSSVnIqqx/OV8X+fGBUNDA4OKwNIDfurExb29rQ2snrkEdF8LxYXlqy6stmU0AFGRV8dvg7/0aZRno9sP30Z2E7DKgwaTuCQNXqFi6dP4uVlfsYGxnEQPBcItjDYxTo2UD/pDolIIsgCL+8vmrSDLU6hgYGJEPoVfugdBGgdcw2eQQq+rQWc8PPzSsZI854EDNkaVHnYLt8nadvRT5PhiOZE5TayssTiXKDZO6RBeHHcOknXjuTGwRieK38940bNNMuw4EK2xwzkULJo1UxKrjm875fu3Y9YlCQUcF28T32u4McXiVKRoUngAh4cPwYW5Jxjm1oXX4yOZdErI4wAfK9GMRgjE/Pkh4sL69hfX0VAwM0Hre13+cnxVtt7C8el33mySJLlJCVad+1qkCvSDQ9av4kGRXuUcENOvtmY3M9+LHE99eKEFIoFDMYFlBxBPke3rvtZtoee/lcn5zLu0Xq7XN8S0jfIevygGns6HRicT30q/N3uiWQH7Zav2tzdmqrihHiV9RP7U2NssMPe93/fEBF13vdCUXYloSO9Z/sCrZfR7K/o17x5HmXPWG3WKLb+Ogae4T70A0Q8eO13EqSssJ1tjwT3UCSLh3YrXDDk/DtX2OXdLsOS3Rufynxq0S1+bf5HTC5qHjL3QI4dairJEjP80eARFtbXDrL724yyWx9ZO+YBF6cmG9p8bb+s7N1Z2B4cZb1GD/n87x9Jx5rybm3IxjjwENbG5y1npR7sk5MHDt5nlB57zJJ3n4HgbywT39nwZKOk+xV65Fklbon73UPW2SnLBnrwEh0/cFDJBzJ7r97IQXDZp7XTYoF/YfrF6AS9hj8mxkkG6PZPTPE8AixtpnJGzjD/YeDJnY8ejj4vW5FxmImUwx/SXoy5AlsrFhFvt9LsY/lo2CySNy0+WfUnuCz4TJUDMyMocFXkAlirk2pJovB+X1eo8VbttdLsijkcRD6QJJJAeDg1bhBtPnVeBxg18B/Mwfj1yF5IYIPjJ/Dk+R9LtlagRvGGuFLspphH9apKJrtTfpfeKEl2/LH/1dcVPU7v0c/Sh7bEvZipHDMMP7jflVgCgEBk+5yDxLzlbE8hElqVZXvMDaLTRCtj0qY3W2SCgCl9buNIzuPgLsgP2Z5C9tvas+YYETx+iUpRvlR+fgZcOKFKh4LyVeFHmjR/s+eCSsKCx4k8nlpe64SbFEBNo88KjquH4/++AnugSRQEQdZSSpl0g7LqzY6ARX2IG8jeipRlwjo9JCF8KVlYYuBCFU6dpB9ihfltoiv5Z/+FMd/9KCm9TZ1BlvsHB0iyjChdZJ/ClNY2yiIrzo6WvsMs23cdIpk2xgV/h3/6McxKpLVxR2Dz+Q5t5/fryLZ9/67G/1wYSJ6zwWAiXlKM1D+gQlcJlgovcCEBX/n3136SfTCoO9niyApeTklepm8FwhB1kWtropDmWkHoIIGV5R+YtJLQMVgfzDTNkbBjkCFgtwUyKigRFGVUj3Bo4ILjAy2yHII0lTaYAfKXkQ5lJ55VdIZlJ0apnkwk+dEulkJwQoCmghXacQVqIruc5FNiWnASn75R8isdFOSRkyCM5HiRprJqmr24+TUJOavXsOFM+cSQEU/ZubmMDhsZtnGljB9bAcqKFUyRHkqJuQ2TXbLkxKU0WJfCwDa2ooMtfk++/3q9atYXVnVU0FmRW/Q3WbymolqvqT9KTNe28xRd52mrPmCGXMzwZJkVAwODRotlQFhCIYEVOhoDAQsScyxxIDLGTg0RyejwgJgCwx4/z/44ANMTEzi0JFDZuQ9MaEkklgj9MlgYJBJg+auXvUgI/MgO5VN1SLN1UymB5SUunrlqoCKs6fPYHRsTIyKuQMHxDBhcKTEHO/dVgm10hY211Yx0NePhoAK29DYTBoDFX/xZ3+O3//GN7B//yyaWRjYAQIuRtG13yuC0qgR7kAFpZ/YJ88dP4bRFqCiEZm+a+bKpmSQyzH16quvoq9QlEeFSYGwMqaGzfIGqrWyVaGkGNDSTPskGjUCFS8oqehAhQVmTVSb9QioePnFL4lRsVkuibNuHhwNLBCo+OgjARVMbPNZqTaq2hbKTPudd8SomJ2esWejblJXvLaDBw+KUeH3hvPIifffx+zMDKZ2TRnJqlaPdOEJbOwEFsRVWLaB8n97QN0pUdWaqLONdJy4a91YPzBQoXUjBipscwclVEdHWVneupP247pPBf/tc4BP/fpMM416heaOPaiVy7hw4UO8d+LH2H9gCkeePIieXBE9WWr29wNNAzxr9bKBL6FSuX3TrKY2wkY5RaCmjHff/jGK+TSOHD6Anr5xKPkbCgd8k8J7T5P79ZVlGUrn8mVkMnXs23sEt2+WcOXaKcwdmMbE5GHU0K9n/vQHP8Pq8gKOHTuKdH4CVRRw/+4C3nztL/E//OavoVCYwvytVZw+fRIzM5O4dfMG7t+9h+uXL2NyqoiZuSmUq6yST2Nqaga798yiUBxCAz1iCG1UtvDaD98QkHv7xg2MjY3g8OH9GB0Z0vJuxUesGOP6UcLm+hrK5RLymSwGB4oYHutHhusC0rh08TquXL6l5Dar3mnyvLBwFQvzV9CsV/D0M0/hyOOfQrU5iGaKfhN9SGfo6QGBFNyktAMVzmrjfOvANO8N/04QjvfYGRVDwaOCoHYrUEH5vpzmLQcquA1fWlpSYr2vz6rpOI+69JPLDvD6y9WqeTWwUi7dg5wDFX05LC4u6VwCKlJprK+ZL9BqaR1NAryBUSHAgd4OS4HZAERAhbMrkkAFfx8dHhWDJAlUkIUnRsWFM1hbXRJQ0d9Htgg9dyyBQEZFIV/QPaOBNftjaY3sEduoDvYPmHcHr1nyTza3MsmvNYAeFTQHl18Fr9uO4xKIDlSokjLfE202mXQnGMHkOTeSlCQiUEFGBdcYSrglpZ98Q08QSUnzILFIjwqy7whUyNcpJHgMqFiTpwiBHyb4r169pt/JjuCcTUYF7yHBriR4yn6h9KFvxHkc3ptOQEWcTGit5kyGofG8aHEw18LlpTWsbxAAMUaFnSueD5MMML92ByqcTWIbbfuugxX8m8lhmDwWPSrIqCAgRCCK7BWOvdW1VZRKLOIwQIPfd6YkwRgCFSOjgxjvPSgPkxaggmOaMco/Qvqp47bOJo5OOequxUndcvyWOO6UtO+0Dwit6e7I/M+yC+3kAxCdspNcFtcnzXRh9xiarv91xSO6vbETCNP2XvuW8gGvvivekrLiAO3lQjza8lyE96LT7pjIt0Re9LJQsHuHdO2Ozgl7O1KnMRjt1uz8ifO2tCfRdp0hvvC4zQ8JVIjZG43nmAXQabjuBFJYA0IyOiREo+to6ce4f60vtndi9IlQ0R6NR6k8xNet9iQ8KghUtB/NE7w2PvxZJHAS+2m2DMFO7VHOt/PN5v0xk173g/CTdE/+dwV6ut07JfnNENyTpioK5X8hkevJecWdysO0Dlt93z0KE03k5wXohHFuOZfYPJnnMRYFGRlk7lpcLoZkuRyS+kziWrGDErpuwCx2hclhyaCaCf+66fnb8LUksfbfYZ2xJDyLMGyPwcIDggJaO+RjYEl0Vvy7NwXXDgIbdm5b43guO4uBAFzTXWLK+ihI92gOTN5bi6N9T8eiBWMCWOLZQUPGCN0xyAAAIABJREFUwpaoNlN3roN2bcHriqbbLCLMMa61AkQm2Q3IofqESWRT34r3VL6DYa/rSfMoKR5ADf07FHmZT4JV+3Ofp/0e2TICVghQxEoHvDy7Xph8Va2qXIn9TmDHt/IuZ9TGBA/3SsUk8iyhkkMAWMQUsPhAgEtgW/7Jf4zZEf/T11nwyZxAWfkNL0KzIh9nixvDgfdGjJsA7rDv2Mku3+Z7H8UuLCkK7B3Gdxp/LFJtk/rWsQLDhf0sDpFii6Ay4uPWfSXC/OXLiRmW2/PNc6iglMxdP2YAMfgMOePJ9p8ub2Zt4znZ37zfbD85NMn97COg4gGDgUcf++T0QGegIjnlJoEKLT1dGBV+zTate2CkIELRSjJws0ncgov479HCEyb8xDu2IEUVLm2BfDhcS68r4eJRRYyyx595GKAizMAdfCqS4E7y/ElwpqW1bQt/60jptEHpBlSEvvulAhVmDCWggosWgYpqDFRsBH8BJtg3NwlWGFBBM20maHwx8kWDE3BvMR9qyW1yZrW4AxUMFIqSfsqDQAUXFQYflOzpGwweFaKZ1iUP0Y1R4cm2SUo/7ZqU9JNrPTKISQIVXlWtsRmqAZUEkYZ4RcnWYl8fhkZH7FbWyaigKTMXbtOI5KIXJTwDA4GMijoTWGQ2pFKq/KWsEdvMRdwYFb2hYscCnhJBnt27cP3KVZw/fTYCKor9A5jdvx+Dw0NaBBmEWYKesk4VVCpl9OTSAiq42JaCb4Zv+KkVzh+v5nQtbL5PWYrFpUUBBkuLS1hfW0e+xxgfDJ5qKTfe4vOcRkpeeAwMs8jlyQ4x0IWyHOwn96ggUKH7G+i3bFdWMiB8GRU4CVS4pwlBCvaTPEVSIeFUreO9905gYnICRx47gt5CUYm6sdFRAVGSlQhRlFeccMyxqplamNTFrpXXlBjh2KKsCBOADCpc+ol98qUvfUmMCl63aMIEKiT9VEKFoNzKilVD05siKy0BJdpkNo2sGBXf/pNv4d//u9/D7OwM0MNKFkuk8J55kt6BCgJxBCq4X3j99TcUUBKoGElIPyngFxvDguRmmom9OnoyWXznO9+RufcrL71sFaus2slQt5WA4mYI4jPY2qrh5Pvvoymg4kVdOxN5pOJKK7fRRKVRa2FUkL2zVSmbxFWa1bANmYWfIaPi6FFMjI3puzWY+RrHzztvv4MD+/djbmY2bEaoi5rBa6+9JjPt6elp9QHHHQPLkycJVMwKdGIVFH0qKEfGPn7yySe7V+QlAAZtoNr+Ha1UbYkX/1yy4jfaCLUt6TsBFS0fDUlxZ1RwfLuEGrXqe3tz26Sf2sGKJFBh7/GaODc2kevpR3WLc+AWzp47gdNn3sXsoUkcODyHTHoA/YVdSIPeEmRVlKwKvlBUAjSZbLQ1u4kUxxMZB7AKsOX7t/HOW2/gVz79FIZ2TSGjCnj7tPeNPre4gtOnTmHx3jyefmYWfX057Nv3GG7fKuHi5RM4TFbGxBGUG5ZoPvPh21hbXsDRY8eQyo3JTPvunet460d/g3/7G19Bb+8Urs7fx0enT2Bq16CMiPPpPM6e/hC5fAWf+/ynMDq+F/ML9zAzexgTE3vlo1FvZlAqV7GysYEf/vA1zM7sx9rysqrBn3rqcRSKZG2RLVSVHFSZUkb1MnqyaQwO9GFkcAjZdArLq/clA5RJ53Hi5x/h5s1l7JuextBwH3K5NM6d+wh3bi7g8ScO4emnP4WNUgO5gb1iU+TyTIbnVOFVrVf0s7VZVZLcGRUOVEiWrzcfdIurEVDBvu0EVHgywyr4Oc8mgYqyNtSL9++hUOxV4jsJVPDZMqCC8nbAVsWACraTQEWW0n5NoG8gHwEVw0Nc11JYXVnTc7SyuQ5SzQf6+9VWB4FXl5dN9xhNrfFkgfCVZFSsrK7qGGOjYyYfQUZFkAYo9PahWtnCxQtkwaxEQAXXAnpU8FUs9KLQW0C9UhUTjucno4LnbWdUcO1wqQ7KUjlQYYbYVuHHzR6BCq/oF+DiZtpB+snAC/pD5JU8N8YGTdxppn1HoJIzKiw5E9Ia9NvSehIDFUlGBY/jySCXAuvra2VUeLEC530CFTxWJOsUEv7sFwIV7YwKXhOTLTRNd0ZFcl7baf6yODwAFekeeVSsbRAAKaCnh7G0GzyGNSfMsR7H8fsOVHDdVNIoSDwl2SDaZAc5CXlZVSuRRwWBK65DjK9XVlf0rDKeSYI0DkoV+3owOjqM0fxMACqCVCXX6AcAKromDzsl5m3Seyh84eGBinh+bVt2tsvu+ge6ggLbjrDjH0wOr8uupGN/hIRmskTNt17qq06n+yUCFV2keigRk3y178S2bbO6gVXtlxuSg9oPdpMJ6rTtU991ASoSiXevbtZp3YvK1Qf8MQ7xT0vTQkJZQ7nT+R8WqNBjYWCPtkq+r287jveynb77OIiMYVsAl85D14EKj988Lokkjfw8hpCE4pq4WjoCWTpsqb0LDYzb/opzEi21lV2vreu8q6S4sbkdhI0r8O288Xd93u3cH93ZLeZ/5/JH0vKXsbOBBy7vY4nU7RJV6t9wShMBDu1S4p0FSwZMuLGztTkGcpT0D2uLKtI1xC2xzvWZYIlhTsHQOeyz/XqMfW+JaMXRkikylo36KjwvPvb0tyBfFYMfVrih5H5iMMp7wVUTWGQWkvLRNTYtH8EiBgc8DFwwI+g43+MHdTkfA91U9d9oGHOWQIBAHXte5GcglocVrLlfJN9jwppHNKnK2FxbQBMZHgIWbNw4WCSj6CxluJoBkLI9lRghwT+Bn1eeI9xG7iO591URBwvlWEihQoLAQiFzgQyiZiPIR1lBpAE6lj/xl9b7UHTnABLfSxMMURtsjPNYLG5U2wQOGdOV+RX/3B//31bQwddvf4NATVbsXgE6YuU4q95YK5WK7Sn9udWeOjApeAyOzeQzyL4n6KEioc2NINPJvrXY1PZesQeGwCfJWwU/iJAX4jmi2Syw3g1oI/Mj9sFg0YmNc9tbS5I09JXAFYJNZIUE5kc8/ghM2T7b5LGMTaJnksBF8HJRjPeIUdF5Ynz0109uD8Rm2gFgCNWSUQwRgtMYeGhHjrV0JDpgO1Dhj3CM+lnS12bXVpkkLTyJ6DYJVvxTgApb4JLtfFigorXy1YCWuHKkNdprM/fqzNHoMGgeDqgI4cq2vo8WDJfh6rbhsmU/Ue2z/fw7Myo+Hqggq8KMQGOgImJUBNTcFw55VORZJWBotRLZVTM8olEzQZFCsSjdRVbZy6SqWpO5Ev0ZmEAWlCagomJGzuUKrl29iupWqUX6iYsFGRW7pnahwqQ3gx5VEJqOpypAJH/DhdN0ObXYJmiETCRRoz+XL2BklJrwtjGTZ4BkUJjsZVKY7I/wfQZZaQYgRkulhBU35NQA31hjErFXusus7pD0U42BJOWoWJlbwcjEiDEqTp9FNt2DPXv3gh4Vc/sPYIBSMmnrN7EyQhUJq9Oz2ZQScWxgRX1WiStNtioCIHjtpa2Szk2ZLN4XAhiUO5GpZ6Uqbe7Fe/cla9HbV0CapqOq5jDNSFZkq/Il3EsGclxYKf1E3wjqefO4A0ODoWrfgi8GrNIrV1LDDLC4aHNBZuKL7eCxDKiglwcrY8ykbHNzC++fPImx8Qk89sQTqkTl+xwnM7Oz0iXn8ehhEicZKK1SxsrSEu7eu4v1VV5TTt8d6GcCmUmZnICK7/zNdyRl9dJLLwmooFSLxkGPjQuaulK2i1XZTESqYiYwdPREaU5L4/rVeXzrz76F3/vmNzE3N4tUj8myKDFfqUQVIgT9eAwCMUoKNYE3CFQ0Gnj2OUo/jSq4IbtFgZT0Kk0eQSI87MtsFn/7t3+rxOuXXnzJAl7X1W02dO00gieoVKVHxcn3xah4/vjzos5Kn1RTpNGkK6jh3JnTkn760vMvmEdFrQorwLekNiXJzpw5g2ePHpOuv8ZiygJdSni9+847ODC3HzPTM7oPvqF57fXXxKjg3/lM8DmUmfapU2JZTE5MWuDZaOLylcsKIJ/59DNWDeUgRGLPa5V9Nt/73OJA4U4JuiSgkZyck8eIA8cHzwy1wfRWQUN5tHwOI0MDer7bN9kOsHT6v7WBerMMdrOmXkQpn/IGTp58FxcvncBjj+3H3NxBpFM9GBgYAtL9qNcLqJQ5N/AnSCcIWDQtekvG8H4ZU0iSTs063nn7TdSqJXzmVx5DnvNTivNsAWhSA5ibJDKjMli8cxMn3nsD+2fH0TdQxMzMk7hzt4Tz53+Oxx47gPHJg6jUC9qonT/zCyzeuYpnnzuOdH4UtVQOd25fx9tvfA+/9Rv/BrnCGC5fvonLF84gm9vE6updzO47jDd/8jZqzXUcPfo09h88iPurFQyNTGOwbxKpRg61ZhPLlGa6eR8XL1xEPp9FXy+B0l48+cQh1OsVlDapub+mMdjb24PhEVbF05i+hpXlZTDpfunKZWSzeUzv248TvziDcqmJPdP7kOtN4/7dm7gxfw5jY0U8d/w4Uul+3LyzgeHJOX0nlysIvCPAJ9C8WhaYSaCCYC3nUYL2XLukhdyb0w/XMYKnTH5ziGhdGxgScCrD5Y0NPQN8Nq1iPqX1UmbXmyXQl4lg8b379yT7xEp/zk+cY1xaymn4ZH1R8klgCquz0j26/1zr+gdyuHvvnp79wYEhsUpW19YUla2yDQD6+/q1sZNWcrWqeZRjiu9xDSFQwXHO6xGnrCenhDPXCko/qSCAFWU0xAyyTtUKmUHnBB6NjAyKEaIEQ80KTXhNnJcpB0mwcn1tDSsbtm6J/UHpJybotUYTqLAx7kAF7wXBBpOXMKYLvTEkt5i1issVMRfM3Nwr3yS7lMsr9uDnGOtRQpBABa+T986AAc6xFvvR54ibTR6LVZhkuDmjgpJvAivplcEYgAzUzY1wfTGjIsmqdFYHixfI6NO0G+I6amjzmh185xqk9oTqTQcqWuPfUHSUYEb4HGmf45rCeCcrjwrKnfX3F5DJ2vqenFsFuIRqVp93Ce5wTXOfLa09XjGpGChUxoZ132QwKmJu8h7zJ9eT1xhk/EG2kwMVDlZYQi+Nvv68zLRHc9MJoMKk0RgjWMVia/yf7ItOa0J7X7UE68nEZ8sbnTPOnfOxxrZ82BcLER70pfn8wT8e4ldnzcdnsTqzrtl0q6SP9omtrdteUd+9Ua0CUi0r8PYLSVxXt5Z17Kcu/dGeiP5nASqSB/EkeadG7QhUdGhw+FPLuPVjBABCUEECqIhZkK39qvjiYYCKbuMp7Oe94jou4GtlOzwYUBGS8pEBrwGD3ceH7R+iV+hrVeGHgshkEtFYwAmgIsSWDvq0SG5FVfudgYoYnA1n98+HRHz77d4p/myPOeMEaaucth+j27G6n8P2xub9EJLJgYmQTOEkZYscnIhi4E7338cjgYoEy0DXkygSSjLv+BXu77SOBY1+xh5UIIgBjZjVrLVYsQ8Z+JacZjvF4miTHoyAigC22DrrFfsybAt7DwNnOLa4jpihtFXzu4yPivkoQx2SzTyvs16UtJZZd/sDZBE/p0WuWYzjfD1hAr5Wr6InJJkNh7Ne4Dnt+JaA5/rJa2Tifau6pfjD2RRcg2OZID+fJdDFWJFPRRUZGkqHKnzGh3yPIISn39z0WVK8lKGS8beBWX4NzsJxtgvjJrFNmnXti1mEZsCBjS/FmKEAMVYzMbaNpLgC2CSGQ5CDZP9wv03lhAj0aDTxx/8xBip+5xvWLvU/71fNcgvsJwN8CH7Y2PCx53teA5dsHfNH38A404zjd1VQmmaBiUlkcf+TnFf8ubF+ifeYHgvxs8y7MN7yGF0+KCpOC74jdZN048ufRWfo8G8qWhSjJYAQYWh5/OSADgEP3xv2KAav6DxStngEVDxoiPToc5+UHviD/+2VEGP6ZOtPRiK7LjAhGQm1r1YPBlT4Jsb6JiRnokm6PTCNg2OHPv5RQEU4VxRIR9fxkEDFtg3CTkCF5/5DPyWC/J2D6ocEKrQ+td0LjzotQxqufqezbr93baFsmPP9PPEkrYq4NkbFVmVLVE4ml41BQaBi3X4PjAp6VHiFvE+2PImo/T1GGVVwESrueR6aMzYbKRk1M5nsRswm/VRVYt2AClsAmNgXnbFaxbWrV1ApbURABauFGfiMT05havcUqqoocSDCkhi+0NZrZoTt7ycTnuVqRUEGpXJGKf2kLrLK7yYXkobJ+RDQcBqrVTWSlmgLLWWYuCk3oGJT0lbMr7Byg7RYskWymbQYIkq+D/ZiQR4V55BNZbFn7z70FvuUtBsYHtT5GQwwqGACRYkyGXVB0g2W+KmpcoHXwmQvgxQm2tk2JpbYb66TTpCJSQcmz8RwKJdx88YNaW0zUVVgQqy3EKrE00rIUNdaAVHWdkpWBZDVMWh4zQqGoZFhk21iMBYWblXVhPueXJiZxKFkBo+zVdrAJoEKBatG/1xfLympPTI6hseefEpgj9M/h4cH0UdZkXodk7snzSzMyk+QThOI2cTCwjxu37wujwuOK+55qLFOyRX2/9/8zXeUcHnllZcFCBGoYANois4YlUHC+vqaADlKc/AalJRxyR8BFSlcvzaPb3/7L/D1r39dngz072Byz4GKmFFRtY0UjxOAxB/96A0BX889+xzGJsciQ10P0n3DRNaEBdfpCKh46UsEKph4sydbsk685+UtUW/JwDh10qSfjh8/jiy9X6IqHaNQl1M1XDh7Frfm5/Hi8efld1JjZbrMiG1OIGOEMlnHvnhUzwPbX0sbUMFg9t133sX+uTnMTE9H0xbb+trrr+PggQOYmZmJqNIGVHwg8IIG2n59ly5d0rT2xKeeEFvEJiezjfYXK17aXw8CVDzMmt2+Gfy4xFfy2P5ZPiMTI8NiH3UCKnxj5+dKVsr578n5U4nKtVWcPPEzXLl4Gp/7zKcxM7cHzXQNhb5dAMZRp1l2aitaN0z+2IAKM95u7TszI17Fa//wX/GFLx4EjdyLhRHUa0WkUBSojDQlpbLINKqYv34C9eqqQMeZuadw+94mzp15F088fgBjE/tRaxa0Ibhw5gRu37yM48+9gEzvKOqZLO7cuoZ3f/zf8Fu/8etI5fpx/vw1LN1ZQDN1H5XqGg7OfQrf/dsfYqu2imePPY3Dh+ZQyQ6gp3cXcukRpGsZmbcvl9bw05/+AqPDQ5i/fgW7p0YxvW8SI0N92FhbQSpFCaBejI2NBamdMhZuzOPmzZuqYl1aWcL9e/ewby/H5AGc+MVppNO9mJyawNLaPSxcOY+BQgNHjz2N6dn9uLeYxvUbGxidmlZCnkltJnjN8I7MiC1sbjERTUYFzbSrqoLnM8b5Ntfbo6p8zq0u/cTxws0VpYXsOzWTP6yzsi8AFVmaKvK5ZpXZhryGeA/v3bsnxkGhNwYq3ERba6KeW84Bpg2s9SHDDS1kAF0YyOLunTtKtvcX+/V/rk8ca2sblMsD+vr71HbO/dwoEuAhcMJnMwIqMhmBCfxeLp9TwpnrEo3kBUKLFZlGutlEMU+gxoAKbuRHhofECjH5ASsQIIuDkoKcSwj48NhrmxvGHGg0MTQ4GBl623pt2s1kSZgHQkMMCkkL1CpKitAsnJWEvH728cqKMRf4TPpzagbbuQBUZDVnklFx9+49ge8ms0jgiIAJNAbZZ2Qf9dIYmj4iSMlMm6A61yQrfjDmmN93MhbYnywsoPQT1xwHgsj649rCtvFvyViaa5YB/I1oDXLghLGE4jSvcGyZ5EwuwecXS1pYbES/CAEVqSxWVsxMu3/ApJ8sLx2AzjY2Bc/F7zNm4HU5UOHtdbBCUiOhXWJnUse5Wo4YFQZU9Kq1DlSwn9VvoZLWmDAZ9PXnMDQ8iNHcjFioTHgQABPrMfRzlLgN178jEPFxC0G3ZG2Xv3cHKsLi9XHnS7z/MECF+ry7etCDnzVKfnf+itdeb0vutxSw+Xc9cf0wCEp3cMPX/+0t63Yzul1Da0c9EFDxoD0YZ8kf9BtBHqbz+HDZp0j+KTTWE3DOhoqAikTXtzYggFIdtofdyA5JBkHLsULmM2J4eCY0iZQlDrrT3fc5yZ9RzU87ABV23Qk5uzaj4sg43BuckH7yc8Q+HRYaxbtd+5IpSWx/JWOyFjCvC3um5fMdjhclPRMsmE7AQ3Lebj9MV6DCE/ehvxjXRwlRm6C1L2o5dgsA5n3TxihLdBbnAk/0q9+Cn0g0xEIhGt9Tol0V8CxasAp2T4rbPadcqXksOTDhPg2SgArGzRFwEylxWByi6wg+GyZla+wHxh58Q+z6UPihvbZYFk0VH3rxA4/BIjzFIV75HooErDhAUElLHibKA0RSvpQMtT0yYw7tRRLrkPtRWL7GmA+Uhqbfo/krpFBrmnm5/MTo0ZBgU9its+JAvrif56EIoogZEUAhY9Lauitz7gyPU4sK2wzkMKDG2aHeVhu3gSUS7imBCvWvGTFGz4zFV8byV0zha32QlmI7LQ9h5+F1GehgAIeYuQ32exp/9H/GIB2BCrtWi3V4DKlmBOkw/p3jw+IXY+VIqUHHtXvvwIhgT92olJQBnPnKY9lezArjdP0ColrzZO0gIr/jXi4mLWqAjNqbKCphbsafOX7Hx5nAizBeOf58qoyAJLGRrN/i67e4TkVIEaMo9QioeIhV9tFHPyE9QKDC16j4sXKaYbtkUtuq1fIoJh9LR4mtCqK9EsKCA094tyXT9c9EGONJ/pZYtS2yap9HNFt3SMAnAYNtpT7b2xTfQsK1HcCZroyKJE0zWpE69lbrMPlnBCpab6pVLXQsr0qSOLef/2EZFQQqmJghEOFST0yiJIGKqbkjEVCRrMTjAtzTw0pIm4y5sMr4s9HUBpamsKyI5OLEzTlfFoDUVKHPKkglJ4LBcAxUXEZ5MwYqKP3ExZNABRkVnYAKD0pq1dh02u+VgxZMKHBUcEM9MjKihYTruVB0Vh00iHqz0rkcJT0cqGByhecgUEGgQx4Vm2WryE81lBgxoKKqAIcV6UxmpXvTuDF/HRfPXEAGmYhRsf/QQQwOD2tVdPkcfp79K43LbBr9fQQqrILWK0QMqKibOXmapqkGWJg0TAOrq2uSnRgeMlkpXgvvBd+n3wMrbxk0sbKUyR7aavP/AgT4zKhaIVTwNBpKDBKs2LN3j+4XK4o9sW/6ncaoSAIV5nlSMvmrzXX98DtMCrJKpFSq4OTJkxgaGcXjTz6tJJqPDV6/+TOkMbVnSvrgijsYJAgTa2JtdQU3568il+/FxjqBmWUlOyYnmdxN4+//7u+VJKL00/4DBwSIMXhh+6WhXjFz3B2BimYKC/Pz+Na3/9KAigMEPFgVY4FYq/RTDFT4NPXG66+LOfH88eMYnRhVX3jyzUE1BedktARq6Xe/+10MDwzi5ZdeDmavBhxJco1sGfq/1CGPjQ9OnhK4dvz542KWcONgmzdSiBsog8nls7i1MI8XnydQMahkJ9/jMXg/rl65gvPnzuHo57/YEaigR4UxKqYNgAkB3D/88IcCKubm5iL9V0qWEaigHNTU1NQ2oIJeJCPDw0oKi0qdmJ5/2UDFTku/b6oMOGliVPJP+Wjz4pfhAJRWw/bNYzBljAEMgoFGL+b/tzZW8OZPfoyF61fw4otfwN7ZSWyVG+gt7kE6VUwYQFrVV3Ldb2+7VfBk8POfv4Pl+1dw9LlfQbE4gBRoZm7sIRpvp1J5NOX1cBWL968rUTsz9zTu3NvEmdNv41NPHsLo2Cxq6JPk3XkCFQuXcPz4C8gUxtDMZnFj/hLe+9kb+K2v/ToamV58dPoiUFlDrXFX55ibfRJ/+a3vYX3zHo4++ykcOXgAueHdSPWMI9PoR7PKjVwF1XQNf/VX38Hjjx3GndsLGB8dxMQ4zZnJrOjD4CArtnMobZXFcjp99rxYA8YSWMPNhXkxFab3zWHv7hl89OE5FIsj6MmnceHyB6hvbeD40c9iYDCLiakZrKzmMX+rhKGJKc0NvfmCNiNm+Mf5fwtblZIq5lnBX63UNO9TWk3ySflsC1DR32+MCj6DBHcJGhtQsW4m9DXTMiZpIE95vazNowQ/+LzeuXNHDDbOtZx7ef9agYoG6ik7DtvIZ42+CwIUcnkU+9PyXyB7oNBLQ+6Mjs+hsibAIgYqyFpjhd3K0rLWGMYLlAuUmXY2GwEVPD/XEbZnZGhYCWQWNGS5NqAh1gsB34sXL4iFODwyrHvEtb9eZ6VhCv395jlEcJlADIGKja3NsLkOjApJYlmy3SsCyYhQLFCvR1JPNY6TSgVFARWUz2KivB4BFUyKe6UkgQoxCAsFJS3YZ7dv31Yy3oEKJc35nkjCMVDB+amXIAaMUUGAf2Cg35gkQfKA/WVrh0lb8d800+aaw/vs0lBcc3lPTS7L5lz+KBaSVrUBFRGjQvJXVijQCaiQLGECqIgA9gRQQcbWKhkVm2sYGKQcE8GYVu+eZEWrr9sOVLj0k7c3AioSZtpJoIIeFTGjYjtQ4eNZ638EVOQxNDyAkZ5pAyroU0GgQl4lySKTeHb7JwEVbVuU6KgPC1S073X8QDtkcbsBFS0eBMlJvJvc0E6LVPt7HwNUtFTkJ5LRndv0jwAquhkddLsGteFhgBAzA06+Ph6o6DYI2hrV0oyHaRPZjN3PoV11G5oQaoUDkKgnTkU53XGSfwRQsTPCEM1LHreo6Cx5N0KbPw6oSDyp+nZXgCR80OWf9FwHYKPr8ODxwh5Anw/yQT5mHKhIjoGPBSpaihHdu2J7C7qCCH4dLcBxSDwn2CLJ73c71k5ARTSiwriI5kEHRrQmhSRzYKKpaeGGWd9sByrUnVyDuL8Ivg56CqXrb3KnLsUouSeXgaqbLJLWpwAeONgtlj4T7jJijmtlrc7MTNXDKI/aFANlQd2A+xPYWsECRB5QifHAnuA5+Xf5GQR5JzE2WNHuoIuYPUyoWwJciXB5IJARQtkdMgzGCn9tAAAgAElEQVSSI9oS4A7mS1a5Nx8VP3oswr43GSqTOiYzVooO1ZoB91R2CElrFk5Y1TzlXs2vgudgfKEKfjJGnJER2PVK+oekPZPn5ofBr8VeHy6fKAY9q/1lyO2yXAZc8GosCW+Jcm8TC/UYezAn4woN5sOQSNKzcJFsfuYhBNyE/qcXCMEJen5FQEKsWiHppWy2Faj4ZpC+EmDDPUc6Mtb2OUbKCUHKzHNIrs6gtqtvgvyu1CfYd7EvDM8pKSX1bxhnYQ11n5Q4d6mBERgaYV/dqCsGsTEbAxEeq8VsHDs2+9f9Qv3fTFA4sOLfk6RauC/2zAZZ5uDlybbaZx6ZaT9MaPPos5+QHviD//BS1NKIghZYkf5GHNR3SqTbUtEaWOwMVLR+3pea+BjSeE9SjRV8JKOdBwcqwpKRaJ4/5O036EGAikTpQPg6ExzRKxGx20LaxpjuQo9u77vWlnX3qNDi2H5LWnYNrbJaXWP3MNluP1hMt40X4o9nVKiCdLMUDLU3tXlOAhW79z+mxDwXo2RCTkBFjmCDBQPyvCiX9Rkmx1ndx0SPkhWlkiZ6Tvz86Q5U1HDt6qUWoCLFhHo6jdHxyQ5ABZkO1i6+qJvtjApfNJy6xwQvXz1ZY1RYcsqMmBq1Cld3DVoHKhhkiJrHahIxKmpiCpAZIJ+Dck1JdlYzKsFBSh/lPAAxHvr6i0jlU0qkXTx7AZlmBnv27EWhvx8HDh8SS4EHd6ppL42saYSswIeJOJNdElMlGBkTEKG+t0y9M0xIsUKVgFBBfXD/vmm1s/qY3+V9W1xcVDKEyTCySuhNwKRRf3FAiRYmvRjEsVLYTbGTlUK8nl27p1Qp79UBJuNgdfG2yMeVEcbQKanNmxtrklji/cv2GBCzvraJUx98gOGRUZnaumxVMkFD3w/K0ezbt0+VGtTJzxFo0DVtoLSxIqkJJkquXLmixBWBED7fb735MwwODUn66cDBg2JUSHqKgepDABXzBCq+ZYyKAwcOIpMz5oXfEw9uCCRppmGAHwDd1197TRvXdqDCgbqo0qJpwS/H4Pe//30M9Q/glZdeUUWzKMGipfL4KWG5lA9a21jHqfcp/VTD8y88r/FsQAUrOwzgLDUruHDmDG4t3MCXCFQMD6LWqMnIi8fgdQioOHsOX/z8F7oCFftn5+RRIbZJSFYRqKB3BVkmHsgxeXry5CmxLAhUeKLNGRVz++dsDA4OisqdpOv/soGKnZJgDszaXAKMDPSj2FeIko42B7dKqUQBdmIz1M628PtvdHFga6OEv/vB97CyuICvfu04RsaGUan0oK84iXozJ3knr+DifGs/XLM6of6U7trEd1/9c3zhi09hcmoX8rlhNBtkVHD94zxHmb11NGp3cPvmJW3sCFTcvreBMx+9hWeefgIjYzOoB6Di3On3cGvhIo4ffxE9Aip6cP3aBfzizdfw3//m11BP9eLUB2dQyFSxUbolGaCZfU/gz/74b7C8ehO/8sXDeOLIIQzu2g9kRpBp9iPb6MHqxioq6Sr+7gev4siRw8ikmxjq78WuyRGMDA8in8tgZe0+Ll26jPPnL0vWZu+eWQwODOv39fVlXL12GUMj/ZiZmcW+PXtx9sxFDPeP4t7STdy9ex2PHTiE6b0TuHr9Il548Su4fbeJW4tVDIxPiEnCRKv555g+7dZWCeXqFvr7+7R+OaOCSwzn22wuowS0V9YTmPBNFsc4wQoCFZsbXDP5/AagIt1EvtdkiwgkbG6UJBV369YtAecOVHAj6B4NxqhoyMumUuXa6YyKGKgo9BGouCWw1kEXrufcnLcDFW5AubpMU+tWoIKb4w1KP0liK4/Fpfta/4YpJ8XNZqWizSif3WJvLwgeEKighwg9jCjHRfYC970EdAcHh7T2sx/E6Fhbw2aZ12wax5TIciaBJcQtqS5GhfSPyaDoj5IW1GJ2oIL3yxgVy0oq5HImaci5j3/j9ylzwP/zHpB9w5iE/eyMCvu8yS6QviZGRd4YFQQq6FHB51Nm1wQqQqUhGShcV2nU7kDF9evzun8e6xAI57/dKFvLQ5hDVVFIHWvFEwTE+iIdclkddwEqDM+OE54OVNi8bB5F9ONYWVrDxua6gIp83gA4JRwSGuLJ+aiFUdFbiMLK5PF93fOKQANktloYFfkcgQrzuyhXYuknBzv8XvcN5MRSGc7uewRUtG9rHhao6FZKv8N+tpmQ6/V12JNB8d7IN0wS4+8MJHTbXnbauOyY8+9srrzTlvxhgYqP295H8EACJegGJnUuIHND7g6V/G0eFb6Dtjb5vjOczYGKjv1l+8fOXdnlr91tMwwgCHOSWhLus9/WuCvst263MJn0jfYNHMfdxkcyuR+YXs4MCGF0y+2S4EsEVDCBbgmP6LyJhsUgyw6MipZ9vTWyRYoqcfadgIrkXNzi99FS2Bk3rivrpTsdpqXf7bLteKb3H1e/ezI+uo4kaNaWk0/e3zrXGxWBWYI7MiAOSeJk0RrPW92iwbTJFCpRHiRqJVMU5Jh5fzQOxF6w+2RARyxB6N46LUBF8CQwM2kzm3aPBa47blzNvaqtX9Yftjc3Q20ODiX8gy+TpIzljWkyRIxxTKo3roJ3RpORQgjcxOdibOE5C+Is5jtgSW2XPuJj4wUgvPVsH4sXKBHL/uN+mIVAkv4N98/NpD1mUW6ETBR+JiTi2Q+S29J8HQoaw3PI66cagtgjAejlMdk+xVdkPwSJq+g+JCZ37zsvhDPmgk0Jtu8Mz6+KqZz9pCjCxqSS+uY5Kt+GYM79p/+ZexV7/fbvlmPfiLB7Yd+zzZ5HYPGcP/MOCDm45HOOj1cBSUHtgOc3dQeOKduTqyAkCayGudTa7/NBPPr5UfWjGCHm/eL7c4tZ7NrlcRoYGyx2dI8R9+VUsSl94/heAvCQf0lol6tmxM+BFYSKDfNI+unjludH73/SesAYFbbytAdSrWn58EBuqwIKiQ3PrLVHE/q8acF1Mp6Oz5FIqidOrO/4XJDwefMAIgokWoCNAO/bDNgCpIhZoCaHvyfBBCXl/GXGTtYxTu1LrtDWKKvg2A7UcIPYemZ92NoSxVyJPu0oFGqnbw3o2sO+7eBJJ+AoHpcdwkNREVt1MJPjWAFHIviJghstwmaGFZlpV8omdbFZwgZlevj/TVbkcTO+oYQzPSqSZtqehOSGnz9NWHUwN/WcnB2ooEQJpRrc9FmV4UTqa1UlknvyOSUtJQdVrlgVaaWKa9cuY2tjTUnNvsFB+QWwYmJschd2TVH6ySowfSPtiwv7gEAF/+7V68mEOimDPFex0K/KSjOZZLVGFbXKljEqAqPBKncCkp9i5aoZOFFSI5ul7AV9IjYxOjoi6Quep7/Yh3JpS32/vroGaltXMzXcvnETl8+dR7qZwd59+1Ao9mPu4AGMjI8o+cFEGPuFGuUWmDHpD0lneALMgRheV6pBMIWSR01VfPIzxaIlGJgkWFq6r+pOZ1SwmpRABsELSj/R34JyUNevLaC3J49du3abwWjeqli8byPfhhQ9CKxaePfuKVW58nq9UrTRNCaKjzMGZvQk4UK+sb4qnwq2jZX/fFGa4v3338fg0Ag+9enPhHvBe0eJq0C1ladEGpMT40pEsepjaKDPGCbVCrbWV5SUW1tdxc2bt62CmBU+9SZOvHdCEiy//mu/hr3T08FM26i2DGbLWyUlIynNwn7xccRkvDMHmAC+fv06/uzP/hy/+7u/K9PvVIaggo07jnMPYAWUhWjLv98OVPAzPib9ezbdEUCx4PTVV1+VR4UzKkwixYAKJZgZiDfTWF1fw4lfvCcTteefN+knXrdtnCzxVmpUcOncWY29F557Th4V3JTIxKtpdOKFhQWZaX/hc58PwF0atbRVVPEevvWzn8kcm/JPDIq1MjQa+G//8A947LHHML1vXwQQcgx/8MGHApYIaPHF67xw4YL6/cChA5rCR5mQzffqmWPgzuco0rjqsBh7cs36yjc87czBMO0n15S2Y7VvOB0o2Amk2N6cJgo9GVWP+9iP51Yb/+2AhB8jWcXs1+IbXdO4zeDmtXl879W/QL53E7/xm6+gf3AYlWoeud5JpFIE4Uxv3/RBSIvhAusARhuTo9nE+TMf4NLVj/Dc859HsW8EmdQAGg1WhnOFYNV4BXdvn8bK4jyK/QPYN/MpARUfffgzPPPUYxgbn0O5TjmfOi6dOymg4tljzyPfN4F6JoPr187jo/fexte++quopwt4+62fY2woi5W1Bc01e3YdwX/5o79AT76KoVHgc888hYmZw0jnxgRUpKoprG2u4Nqd6yhtrGFifAS7pyYw2E8TZGBtZRFnz57FuUtnce/efQwOjuKZpz+Hgb4xXLt6E+sbJaws38e5C6cxN7cPc3PTOsaVi1ckAVfeWseuXaN4/NARvPfuO/LneOWrX8Ote03cWayhf3RE0kScz/hM8B4x+c35pVTeFJsrn6f0VV3zCyv4ZW5eLGh+ZbLa5XL83hPc4I9/lt/l76qEyxAAoK8PmXCb2CqR/ZcVyMD+onyg5G/C3OoVdgQqkCWgbbKAVtlG8J6fzaJvwI4RARWpDNY3N7ShovQTP0N5PVYKEgDl3MX1ybwwm5J+orwTN9OU6YuAisV7mg/JqGAUw2vNcZOZTqGoisMqLl++pCR5/0B/5FFRr1nMw8o9zq98xgnmcL5dWVuJdIsp1efrsz3nNseYKbolFAhU8FnjPamRUdFv8QQTEVtb9EhY1rWxYML1kMnIEMOxQN8iMhCbmuu4NnK9dkaAsVYthmzSTDtvMmC9rO4P0k+8ZjJ3tO4GkJqSV8ZSzKt9jJMIVLj0E2Mlvs9r5jhxQN83515kwPvLMcTPeRI/CVT4mGKfGFBgcZbPick5zNgWZKdyfV1DqbQZMSqUBElqLSeBkFCNygIHtou+LF4x68CKxwN2HJMusKRCVRKfvb28z0UB5rxWekgRxBAgJIDH5mu/xoFBemr1tzEq+HzQTLtVttPnz53n6W2Re4eVJPwpEX7vlITsdIBUu1nytoxuhxWjE7uge+v+kdJPHfYIXbLKtu0LqfbwGd8idu1jXXfnfUjnS+mcrN/hsg1499uY3CJ1+b0jUNGWkN12vuS2b9vltP0hki5K+Br6AbtnnLuk8+3Y7V+zvbDv5UMA2V793nIRnSGSdgpG5E8ZgAg/ry4/bMBDi9qKFpMJvW0BVMfbZ7fMqoXdVDk6SYKbEe37nW0arjPSxPcqQcug2j5dX+LRg1hZ8jFPePV0itMkYeRzuzMcEqbhLTNGksXS4So7zRP2NwOA7bkxwKklIdpyXMuntLMbFAN2eTD8GpSCCDdR+wsyITz5KjAgmB2zCJAJ5BagxHEd+1z0CDBJG0xxmBDnXoPFXjwP13XdF64nYiTQJyGAA8EPgtcsb0XJAiUGd4J5p3Uj5FzkhxCSwl5JzjW89Tk2jxJKXZKBwLXDX+aRZftM5RzC/Vf7MimxTB0QT3aoKvZZkMiFMXgsSGJIQIUzTezeOWhHAMYMty3Hptg9yCdx32T9lVX7ZJgdfBa4p1GiP0sGhxlii80QzLm9CFHMQcaDZHyI4W6V9WxVxKjQeh8AOYIU1arYsy7NpWIGXZsBTDa/kKVhwIYDPMY8sQTWlpi45qVge9HY1NtiCjNXt2ORiWFSUcp/Ke4ws2mPJWSmnfDz4Hf+9D/FQMXvfNNYDpact5FHQMvjB+2JxTwx5oiDT2yLJfbN18PlliRvLGANyIpBY/MnP6c9eLifvDZ2HnMQJk/t/WztSAI4kV9JeDgYq5IB41OX9Yf1CeNpslI89yYptlRaxX8eG/o1REp6MECLBaDxyxAhB0IeARU7RwaP3v0E9sAf/K/t0k+J6KNrKBECxyjx7knukIhvASvksBsdyeaXOMKzBdO+p9yVnuNEBOi/aubpvAS3LJjR4UOb2oCKME8mmtCWpEqeO/J7YAVGPMEkJwiLKZIRa5jkk6tbhEcE9FhBFROUyQ5uBzzi97qFHq1nTfZZ4vdtfdmpD7e3v/XWxywKW3TsXek2JoGKWhWSfgpSPcaicKDCPSpKoEcFN7HOXEgCFZJ7CIwaTvIyrK5TkoFGnNkIqPDErpJB1YoqMLM5AyoENFSqpu9MM+02oILSTzGjYgqN4Dngm3aBH8HDgdJP/Lt7TDi7guOW0k8MMnrzRSXHmSRyoKJeLctQO3ksO47dd1YNsJ0EKvg9nm9jvYSRkWEz28pmUSSlcovyUk2sr6xJbqcVqEhj795pFPoHsP/QAQyPMjlkARjPS+NqLn6WoEoJqGD7RCENwbsW4QYXfANECFTw/lIvm0HV6toKlleWogQ8k0NMYjEZ4kAFgwVSaW8s3MSZD08LqNi7dw+72QJtJhUkQ2G0T/VzpkfBIPtjYmIC4wQ9BIYwgK1KX9MDHIIKJY6Xes2AipLJRTG5xtfq6gbee+89ST899cxnMDI6EjEVGPj4M1+q8RobMhlnMDIzvVd9xGuvltZRLPQpcUgDbZrH3ru3qCrl998/Kemrf/PVr2J6djZIPxlQkc0QUNsSY4jVwy51oSCX9zvS8qZHxTX8yZ9+G9/85jdx6PBhyck5UMF71A2o4H15g4wKpPDC888LkOoKVKjSldVJ9YhR0Q2oIKOCySi2/cR776FercijggCQ6evHQMVWs4KLZwNQcfw5DA0OoJ5qosJqInkcQB4VZ06fwRc+9ysRUNHI2hxhHhXvYI6MitnZCMBJAhWUhPLAjM++PCoCo0KBXRtQwWddYBDlZAaHYpOyHdbhdqDCn4NOX9kpmdVps/lwIIWNyt4sgQqrFPfxzuN4Ei8JViTbmAQwHKDw79M3pNFIo7pexZs//nucfP91zO0fxZe/+qtI9/QB2WH0ZCgv1IsU2RUPBFQAlc0S3vjJdzF3cBdm5w4hlx1Bs0nWFu8/k4Jl3Fw4heXFGxgaHsL0LIGKTXz0wc/w6acfx/DYDKoNMrVquHDmfdy5eRnPPfsCeopjAiquXTmH0yfewm/++q9howK88+57mBrtRalyH7undmOwuA9/8e1XMTCUxlb1Jo4f+yzGpw+KUbG5Wsfq4go2t9ZRHC5iYmIcYyPDaNSrKJc2cP3qFfNYubWAKtLYs3cOn/705zDQP4yF67dx5fKCQPTbd27i0uVzMiM/eHAG/X05LFy7ikqpjMmpSRw5fBipehZv/fQnKA724ktf+TXculvD7fslDAyPKXHfV+Q860BFVYl1Sj9R8iffSzPxhmSaOE+bmXZB8yvnHq6L7nPD+Y4gxcBAnwAPvl+tGAuC1VbcC9KHyIAK86jg88xqf8rrJaWfOL64CRa1P8GoYBtUxdYGVBCM5qaOcyLnE65T/P76AwAVrP6jFGALUJHvwSKBinQKI4ME9VOobpUjCaRigXT5Gi5duohUqqH1hYl7yS90ACrIGuBatLq+GgEKZFy4lIEl821eItAgQ8x6TSCSsUtM+qkvyElxs1guM1G+bEyGfLyhdUaGmWlntbGcn7+O5aVlrTWMM1xDm+dkyCWggn4S/JFhOCT9xLEw0D+gxEK02a6U5QNDcJ/tc6CC18hjkyVBoIL/dqDCk/6cB/i+WHSBUeFAhea6lEsSxMBnPI8YazE5b/nvDlRwPC0vJYEK61OOwSSjwucg2+hnxLr0seyJAX4vWRDic5yZmTPRwf5nP9A0nUCFARg0Lt8ql8zkPPSbJWcyqqYcGOwViDLcs6/NTNs9KqwyttN1Rn2RrJwMf+wqp9StBr0dePDjdAG8LXGYfHky1SOW7atS9zRk50XvIXGN7mXuXdZUl9zpuH52LYF/WOOMTnuvHRZ5Wwg/5gOtb8cJ4fa/JxP/ifc6MBGSfb3NOjASQQ6jKpnkZize3lz+oQvzpOuVdQU8duqKtqMliAu+N/ctux0+gggS+/jufR0Z1nZqQsf2WtW8J1ijiuHwfcVrwcPQkp9WaegJesaDHgfxd5+XlLIOD5slbO2A21qeLMjzNvNvTI4GBlkEBrlkVMt3whETz3wyVmyPG/3f9vF24/HWRoaUr1oVG0a3XsyOQIVkmAKTOfgUGJhgAImd3gA+JlwdBEnGl74P9kpvm1cTwAdlcwRM2D5EvgxuCi2gwbwleLkmMdR57Ji8UHj2VEhpN0+SQO5lKKaEvRcllkPv+GHVjmC4LGnGADCYf4JVoGstCeunMUlMpYHrmPqackbBb8L9H+RPEbFEzPPCi/+SQ92Pq+OwQI9+lVljYnihQXxtZuJtYzUex/ZEWMEXYxjJNYfzScaqbv3J8ak2KC/DmM6YKtrLBfks9qkMs2mcHQq7BDbIy6NzsaquXebZxuSNrpMJ+9B/3pf+7MWPTnx/PV3I71j/m0+XCqtcBkuyYHZv+Lf//IcJj4pvUl2C48ruh90fXr+BRoozBI5YIY+zXjiMrBDCQCG+pGwR5gdhmCyMDXJP7Eu2gbE8AR2/d+4Nx/+zwyVNFlg7bBOlutg/ZsTtDCUygeyc8TQR94nFaO65YcAQvxnEt1pk/LyvTMrbWNKMmf3f3uePgIqd1rtH730ie+BfBqiwpTQKBVKmTRc9SMlJOFrXExuJlrXr45LohoK2bCr0lYB6RMFV6+0xf/DksZPJ/UT7AwqyI1ChWai1nS0bigRQEVOCbQJONsFkNx781fnTSbmnNsDCg6GOp+h0tBC1tjGpDWimbqgFG2JUhAlzG1CxzUy7BEo/cXOdTM6ySaxssOREkF2iR0Wlos8xgZBK9aC/byCSyVAVQGBzEKhgYkAVHNWaDK2VnCmXce3qZWxtrkeMCjIfuKhT+okyJqk8z+kov9H+XKOQppsaTaH60TfK/AwBEiZvCFRYNWcMVDTkrRGACiVzLZCg7BDvOemlrHxgoooBD5NXTIozwcdEHoMR0T9ZId4EKK3BKvZapp5gVKSxd9+0qkIPHDqEgeEBBUBaSFmB2svqZWOcsP3UPufLF1/+btUCpOAaIMKqAVZq9AUGBYGKpeV7kYEnEybUQCfDgEAFZZCoGc7vrCyv4cOTH2BoeETJ6HqTYIMFEHxZ1Yc95/UGKyIt6OG/ya5gcpH/Z3W3qi8SRp1kLJj57CrKBCpkimaVMBsbJbz99tsYGR3H05/5rNplNN9moOUSaExho2wSG5QoYTumJscxuWtSgU11fVV67GYayz6qyZ9jdXUdP/7xTzR2vvzlX5WZtnlUOKOCDJrYo8KTgwqQA6PCKlIskf9f/suf4fd///clIUVcywOynRgVrLp5/fXXFfQLqBgb7gpU8DwMAHkR3//e9zDYP9CVUaH6lmZa8l2/+PnPUSuXI48KaZYGoELjInhU3L6xgBeOHxdoxgoqByo4e1y7dg1nz5zB5z8bAxXNLJQYpcfKO2+/g4P794tV4bNNO1ChzYlAwKqkn2ZnZ7FrF71C2oGK/drcs6r7xsINHP3iF6Nglfe62ys55yc3jZ1Ahm6f3WmG9uD3wWbxJnKZlJhS5gljLBafa3wz2IlV4QCGlp42DwvycRrNDFburOA//eH/gUKOcjBbmNo7ic8fexbZvhFk04PoyQwj1ewNSzM3QtykWlJv23GbKaTrKVy8cgLXbp7GZz/3K+gv7kI6RVYSq4wy6ElXMX/tBFaXbqB/aEhm2vSo+OiDN/HpZ57A0Mg06ihqvbh47iRuzl8woKIwhno2iyuXz+D8B7/Ab33t13BvZRPvn/gAeyaLSKVL2LNnGhmM4e++/zomp/pw6crb+Morx9A/vht3FqvY2mhiqDiIsYkRFEcLqJZqYnrRz+f/Ze9No+O6zmvBXXOhABTmkQMGzvMskeKsgZKt2LE8tJ3nQbJj53X6vbxer9fq/tfDj16d/HlvdZLu16vTncSxEzke5EGyBkrUTEqUSEmcCRIECGIiQADEjCqgpl77+8659xZQIEVbyWp7qbxkAqiqe88999xzvvPtb+89l5xB57V2TI6NCvOuaeVGNLeuQjTCpHASV692YHh4FFOT0+jobMft0VvYuHElVq9aDmLYl86fQWN9A9as3YBIpBQz40mc+fADlFbGcPDIEfTfSmBgeAYVFTWy5rCKnP2h/g9cw2ZF+kmAiogCFQTwLVBRFCuWNY3yPlKFXszvc47MoKQkJmCFC1RQ29f47oj0E4EKn6wjBCrIhCKQXFtbq0wBswnXTY1uytPcSFGyTmSklFXhBSpK4kHcujUk8whBFwIh9Me4G1AhRZP0s5mblfWQ7ZqZ5nyaRZRAxciwyJJVlFUYj4qkrAHcNHK9sYwKJslLSotFNknXeF2bWWXPfmJMwIT+xMS4sDblmsiQo0k31xhzzbwHfDZGb992El8WbOC5yCBbAFSMKaPCC1TQKJzHpIE313huUAlU3L49KoUFAlSI1AHXNjV0z/nzGRV8ovr7VPqJ/h1BGoeaYgGu8VxnyYCkbBjZC2RUcBzwejkmWKhBkILzhI1BNOnDsUSWC7WtVSpzvkeFZZ5611ONPd2EgHe+0uswIHXWJ+s62xSPFyMY0g2+yj/pyyYu7JzEtnjNtD8+UJHG2BgZFQTuyIIKy2Z8ZGQYieTMAqBCGRV+lJZGUVpWgrLgkt8cqNAJT+c9ZwZcbB1ZpGDqHoGKvGS691Ry+EXOsWi9dOEV518aqNCW5rf17uf8/yFQUcgs2XNZ80eCJg/zX3cEKuR5MmPL2Q+66+wnAVTcqd8LAlyFxpkFKhzfBqsa4HI18pPrCgYsFnJp4vwe7jeLLEQ6yJglmypjmWcEMLDJazP3eIAK6U1jVGxBFgtsuAl1e8+MLs1iT5oXuDQxqSbf7UjQBL3GaJ5xYH9hot8ewwtkFABn3P6zwIR7wAWMCc+os/O/Z8IyCeVFgCNP4t8ycp1kvOk3YWkYphuvislr3afTlFg9Gex8r6wATazLXTZyvXrP1cjYsiokhs3mjKcCmaYq+STAQYGXmiK7kkOs/injPuAAACAASURBVBelApGtVYaMC5S7Ruos+rPV5wQVLOCh7Vc2AO8Zz891nm2018b4hqwGu/e0jErbz+KzYeY7777NAl+2XzT5rJ5REsuzbwwD0fp/MBCyLBYpqJxTXxBN5rvAjJ4vqzGbAW8EqJEEfVb2ucIM8Iwr693AgkTGFlaiSnxeZH9IkAXqfzWrHpxWwqrQPkj2w2lNwjv7ApP/sf1pgYb5QJz9vDyawoRkX+g9UKBCJb4tgOJ+X2WK//kH6lPF1ze+Y9i/UtSgRvD8j/eSxYyM7Wbn1GtTeFkGWGHsLIwWI8euR9PnWAzHDUiijB56ZlgzbH3GbS5ITKvFI04lvSkFSlYE80ASd4qUlOYO7LMgrBGn6NI70HU9sGbZWhhogLdAELMpLbSVNmdzCIV5rzQXNX9OmF8P8ClQUXBK+fSPv8s98IkAFYLGuwu4C0rwb4x87GKUD1Z4Jw7dHJnF3ZOwXxgALdw8/EZAhcwpC4EKTZTN/ztnFJ0i8l8eGu+9ABVyGBcpdis9/qWBikUCGM/EnX99bnmN9ou+q4GIoTAKUMGkh0pcJFOz+YyKAkDF0pXrpQJUvBJMJTmPy4UgWkSwQceLTd7yM5RZsIwKm6yQ7zIRPzcnCX4CFWwjFxL+jRV4s8kZASpmZ2ZQWlaG0nicwk8y1ghUVDXWISBAhUksezwDuJKk02QYuOaRqtmo944mWlwkI+Ei8Wtg0oVgk8hVpeitodRSJqSEmid0WIIkhlGRzWF6SnXHrewSE/VCRw3RyJRABZkZWUyMj2ty2J/G4M2buHalXYyrly5dJsmW1hUrUVyhlZpctBnUk5HBxY8LKZNBAlSYQM0CBEyY8DngIsgEopWAKjVJmcmpcYyNjRj0nkDBlANUsGqXAQ6TGAzEbg0Oo+1SG6qra9HS0iQBH2W/mNihJAoDJgloJFDSJJKt0BEGSCwmIEO8tAgBmqo7uQP1xuBiPj01KW3kSxM2fgEXBKioqMSmLdsE8NCg1GPa5gOmU7MYnxjX82cZ5PlRXhZHSWkposhIcoRJId4vMlo4QzB5+atfPSeSHIcOH8Ky5U0iHcV+Zhu5b2HCa2qKyRxWfaoxsiTLrNGWYS4QqHj6n36M736HQEWrSFGpJqbKnFlGhXpUGCNyMYfP4s033pSxQ6CiXIAKDRx5He4zpBVmApjlfHj+1y+gIh6XdodYfSparArCSQ0OadZZmsGl8dEHH4qE1d69DxjpJwtUaGA0m8ug/Uob+nv7cGDfXmEB8P6xwieb05nUAhXbt22X+yhBml+F/yjX9f7772FF6wo0LV/uMXnM4ZVjx7B27VosX7bcqe4Sj4qz58Rgm0AFpx6Oa5F+CgawgtJPgJif0xtj/959jpeM1W39OOuyfbYldL0DwGHnPXvMOwEehYL1+W3R7zNRmENZaRx83uwKY4+tCUYXsLOJRnss7+9eMEOAiqwfuZQfZ0+9i3Nn3sa2rU1o7ziL6ro6bN65B8WxavhQgkCghFaDWlFlVzi7DBmAWjdifvhzlFYaxJnz76K6mmDkaoSDJfD7w8gijLA/hb7uc5gYI+MqjuUtGzA0ksDFC+9hy5Z1iJc3GI8KoKvjIvp7ruD++3cjXFyLbCCIzo423Gg7h888ehiDw+O43NaOhroSRIt8aGhYhlSyCO8e/wjVtcX48MNX8PBD21G3rAmz6RhikWoUhUuQTE1jdHoY7ZfaZT7r6elWVlo2i+VLl2H1qtUoq1kCXyAs1Uu3Bodwpe0aZhKzGBq8havtbQgEMti0aQVWrlyC4qIguru6sH71BpRW1GFodBbZlB/nPnofVVVFOPjIYfQSqBhJory8SsBlARqgmsvJWSaPk5hLzwqjjZXilG8iUMEKLrKZpHI+HFGgQhLNJWatzQmzjX4MBBM4B5LtRTCCayU3fZyLLFCRTCQdo+e6+jpZD23SnpX9nNdk88812+jgcu7gsTlncKPFCrzSkqjM8WRE0PeBxx+fmJDvT80kZB4qiikDxJp0c33Sx0eBCsqZcQNIbyVuziPhIEZH6FERQEUZ2RZ+kV4KBEPCDimOFck81tnRIe/xusUnSYwmNSFCdgfll2aTs7JWsPo+OTcjj4MXqOD8znWJSQs+IyPD6o3B4wgjwRhrMvFBU+5IiIBOUMBRxhlFsYj6F0kyQddeF6igNnRExpUCFWRDKVChAKN6/yDgE+mnqGFUcC2gRxHnXms0bucetmN8YkyBiqIiAf57e/uEVWKBCrbLC1TY+YrH8AIVXL/ypZ+YGMho9aoF/k1mhXOP1fm2a62Nw51kD4GK0QkkktPC7FGgwlRuekAKW3HJ9nDeJ4uFaxrvoUoS6D1U7WpdH22hCceyZblY6Sc+J4wbKHPAY80kpqWQxQJRdlwTqCgpjSL+SQAVbsBhpth7AyrumY6wGOjwOwZULLrOFkjK6mfvIXHtrIp32rsUaMGi5y7c2oLJ9E8UqCgA6EhTTKLfLv5OgLG46fhi8UUhoGLHA9uw84FtKC7V+OJ6+w38/B9/5XbCvH5yatm8CgYmLnrgwd2478BOKah64WdH0dPZ47a/YOwkgYNHvii/7xeF4jwJb+0h7SOR9VkAVKiKqU5pxiPD7FGdOc1k8u2cpq0wz7YXkJg/NLwAg8xfC2PE+VXSzu+eqWM+YMHfV21YJWdrv9juySt4esQ5kAdisvtvU5jJd5pXteCL3/oyYiXFOPHKW3jt1686SeuahlrUL6nHQN8Ahm7ecmYbyzoRyR29KPV/4Nxt7qOtCmdcYPdRUuwg5sNM7moC3rk/9j4bIIeXL8laqHKAzPeSuFe2N+Mxxifq77DwJWsjjyUG22RX6PqhXkaUXFbJQP6N8ZSTAzKSYTJeJPHP74RlX8fj8fqUvZfTvTsZi8mEs9+TSn16bZn+53pt1xoBVwz7gGuXjSmY/3Akf8w+wiaYub/jdTM+kfb6da9npa8c4+wUCx4jhh1gyDWmWwT0YYLfAuHcbzHxbu6ZDnu30JfXxr1tOsM9pQJMUpNGSSmRwFTgiTGhBRrYTjv65u+DLGOFe3j2va7xXL9V8skWQkjRoykoW/goGSBL2qn9630eXXBB75kFR57+viv99K3vKpvYFnIREGCbNXY1c4SAWPP6z/Gf0XNbBpDNP6g0mSBE8kUpxOC+OpWSogm+JRJOhpXMCcfrQSPxjAEpBLi00lw5ypuqZKXzmgda6jhzAVD18qBcmcv68BaCaP5EpcfU/1MlLr3P0adAReE1/tO//g73wCcGVEhUYB92TyBgaWt57AF3FbfPbd7keEegosCi5qFCujHI3RgVBpCw1S1moloIVJj5y4ngvOf/DYCKBZGMN6JZZGO02J89PhtuqxZhVNx1jBY6CSdNXb7c4Nil0woyLpqIuhBzUU+m5u4KVCxfvVFkG6wXhA0GGIQwSUCggufzJm+5gQ34QyL9ZI1HLdChSQoaaWqFvQInc6LfPZOYRO+NLiRnEigpL0NZaRmCWaWgltfVoWJJHQJhk1y2C45J5ufI1sgmzf7TSBb5WbGpSH4qMyfJ6XAoKkwAbq656EgglWIwRTaEgjhSteDxwSBAwEVpcmJSEiTCTslkJEnFO8HggrJE6VmVyJqaHBeNcyoYDg4MiNY6E21Lly2XqteW1laUVJVJ4ocLGBfa4iIac3uAitISU0Gi1FY+cxo8BQWo4HkEBMjmpBKfgccUgQqaoBpjKCanhoaG5HqFuRAMSh/wWujtcKXtCiorqtDS2oKyslKphLSglKUrahUOq7BNcGVo8Pb3ktIiqTLn9fuYcJKKYWqdQ5J5HBc2WOKY4VgiUFFeXoEtm7eitrYGgYCOZ2WHqj7ozFwKo+NaHcsXxx3bzuM3VpZh6dIlEtBaGim/w+TfL3/xLKJFxdh34IBIqnBTwESdGFSLNElKDeNN4s4GtjboFzoqfOi90YOf/Oin+OMnn1JGRYQU4HyggkEJE5g5I5cnm7RMDm+8/iaC/iD2CVARl3tsq6Stj4tuhdXEC9kAfv3cC6iqqMChg/sRCim9mfkq6T8GR0ILhlTrnD3zEWZnEnhg7wP6OYcqnJW2p7I5XGm7LJXEB/bvk/vDXuXGxQpYEKhoa2vD9u3bUV1FEMvP1kib6LVCoIL+FM1NyxwqMZOSL7/8MtatWycyT3aeYXX4hXPnBaioJVAhrKM02tvbpd0rV6+UzQuNdTuvXcPOHTtRW1PreNosNt3ND8LvBCp4AcpCgfddp1TzgUIAiPyNTBtfBiXRGCpK48ZkzWjcc49mpOMsIOH9V4N51wDSC1QwyM1wM5PxIZWYxhuvvYDZ2UEsWxrHtWttaGhcjs1bdyEUKYc/QD37GHI0LeB3pF0aPLtroXqZEABKZ6bR29uBvv4b2LBujUj8BIMC8yHoS2Ogtw3jt/tREoujuXWDMCouXjyNrdvXo6SsBplcMdKpILo7L+Fm3yXcd/99iBTXI+MPof3KRfRcPY/HHt6P6z396O0fQG1dHBVVccSKy3B7eA5d7f1Ip5O40vYeHn5kC5pbWxAtqkYmHUcy4UN75xVMJ4fR3dUuY2xqakbknVqbV6K5uVXm16xU8ulmpuNqB/p6b0ryu7enV8ycy8qi2LylBc3NdaipimNiNIGWpjUYnc5ieIqU8yjOnj6BpXVhHDy0Bz2DKdwco69CXOYsZa755dkgo4LgQzqXkkR7LBpDhkBFIilVU9Mz0yjhXBIOCXuLz3JxjN/XTVMsFhG/Bsu+0HlaGRV8WU8cy8bgOKBfUP3SJaBRH+dPblojQfWSYMJcpJ9o9k0mWSrlGkMaJkK8qFhYGWTLlZbFJawbHRuTxDJ9PDgnETzhvCv+MJk0JsbGROqPY4drSEV5uVTFzkzxmtSLYmx0VLwe4mTNSYIhJcwCrtMEJniN1651yOaL11daElc956xqXMeKmbgvEi8OJu3HxsfFQ4rzANtA6SfOiXatZWEDvzc8NKSMg3RKmBhch+bSCgyXxEoQNl4INBcfHRtFUXEU4aBbFUnmBsENnlPkFAJhh1HBeZBttUCFPCccWEE/ghGyIkMi/RT0+9HTvRCo4DOmQMW49IFcXzIhQAUBLIIXBJLIUOC95n8W8Lcb/ZnEjCYgyKggiFOsPha2gtRWz+bNdbI8alyiwIPGw/zZVg1roseP2yNjAlSUlMYQCpONSMkMTTZbAMLOP7rppvTTiMRBIiEpG39Nbvl4TyRhpLIbbJMCFZRqmMvzqCB4xPFC6S0WPPAZsdclG3bxX/GjNF4kbftNpZ9swVJe1blJIBSe4xdLmt9jMn0+UJH39UXTuB932dGt0G/ZpLyTfdw6KnvORcGCe+w/ycTd44V8DKBieXMjHv38YZENm/+SuW5iGu1t1/HOm6dE1sP7undGhSc3buMCT/FXwV2tARQ/buwx//bct28Hdh+6X5KwUvySzaL9Ugde+sUr5pBGS99zAnsMWX1s+0zC2AtUvEig4nqvYRNovFDwGozk1YL3Frk/0q/CojDxh6n0l+pzRUMNYGA8zuQZcq/DKfqzWJg5j+457D5W2+qMqAJtmf+ecAY8fpY2EW3loLwgZaGpwwtW7D60G4c+e1jmxeOvvI23jr6lCVLTovxpwOy/nSpBtycXAhVv47XnjzlN+ZP//k/R2LQEt/oH8V/+t7925IusV6BUpbNXrPSMmdM16W4Kacw8LYVdpJcabX29T0bJwiSGWZhmFKT0/kkUxP1wSosgZF+h94vXLmvGImAt2yDPnMgkq2yPgBXCsmDhn+Y5rL+BXetElcJNKmkxFT9vEtoCYOSy6m0QCRvwRMeDSA4ZHz/+bpma8q7x0LCsAtk/G9kreoYJW8A8A861zWNH230nZYzl3CJ9xT14SNiwPLcAQMYvQ02rdaRyl2WvQfIlZl8sBWcGlPGOMfo9cZvLnAjbL3JcMGbZho0guRLxsExLHJbOpvOuwY40u7YrSKRV/SppZUzCzd7Mft7u4+fvreyeXa7HSDC5oIWCEyr7pHEIP/P0990k/x//KeU5Z3U8iToFjb9NQl+8OeecaUi2MSyGoTdJSAEtq1zBnIi9Bv5LoIqgk42pLZjBXID1v2CeQBUgOMY1l2OlpcRc3QBu3r2eu0fzAPOeuUakuozPqlWbkJxYJqf3gwWTIWWPcAyTwZFlEa5RyJAiT3qyZtLweYGmT820C6xFn/7pd7oH/uJPDkv7CyVTCl8Yp06jaegEJ97wxpmuzBSrC5PzkkWtMFDhIqz6fn6RhlkNCzRKwyRPoCQ/Lg5UGGLivOs2319EfkkX7/nBsjc4yw/UvAuwcx00nTXBlhpy6Mv2/WKx9aL3ZiFfWJtYsLrFtm+xgH+xXYhuEpxFh2ZkupK6HhVMeAgFLiXJlzyPigKMivlAhV20OCnHYlE1ODI+EbZaXD0qQpJosIaaFuhwgQpWfzCQ4eRNoCLkABWJaReoCFmgoqEe5Y11CIYjimpbDwWzAWdgP5eeMYGP0gmt4ahQDtOzkuhmhSUT9wRR+BlWlNKjgkAF+8r6XbgJBp8kgRinUJ6E1eNMPvF9VkOSQcGfqdudFtCD/hUTYnAd9OUwOLgIUFGt8lO2GoYSJOxHynGFfAGU0EhcFkKjoWgqVBj0WIkt/uvLZkVHmwvw9NS4JB0s84HJqaEhSj+VCTjE4IXBAwOMgYFBtF2+gvLySrS0NKO8PC7SJPwMEy2sCuVLkkk08/VUgfDvEghL8jWDcCQk8lJMeLHyhmOKC7JIkHh0Ixmgzgcq6utqhe3Ax4AVoErFpfRTCrfHRp3nje2mNAmNP8O5FA4eOCDVswwIpNqEQEVyFr/65XMIh4uw78B+YV+wirk0Xir/sSKJ95n+FKxstXIrllGh0IELVPz46Z/gu099GytXroQvHBBDbfaDBRuEluwFKgzw5gIV+1FZXSY+JraaxXq98OEnrMDkDbJBASoqyytw+NA+6QcmszjmhFHBgFimNL8wKs6dOSOsB5ppW1DKBqic7RWoaENfX68DVPBgwt4xc5kFKnbs2IGqqkpjOiYO8lLV/t7Jd2RcNDeRUaHLAPv4lVdewerVq9HS0uIkvphwO3/WBSo4Pniuq1evyrOzYtUKB6jouNqOjRs2YsmSJY4EigUZ7L+LLdJ3AirubV28tzDAAhUZXxpFoQiqyugbEXRANdo++MhWkUSt6vV6NyI826JAhVSz+eAnaymVwszkMF499hzK4kGUlQZwrf0SljevxKYtu+ALlsIfLEYoUopMxgdfzm4MbCrGu14woTmH6ekxXLz0ESrKS9Ha0iLzX85fgqAvg4HeKxi/fROlxXE0tW7E4NAULl86jW3bNyBWXqlAxVwIXe0X0NtzAXv23I+i0kZk/BFcvXwefdcu4siDe3HmwmUk0ylUVrGKm7rHPkxNADNTaQzc7MbURD927GjFqrWrEI1WYGY6hEQihwuXz2N8ehAjt/pEhqehYSlWr1qPmuoGREL0x/Ah7cvI2OO8S0+dsdEJmYe7OrvQf7MPNTVxbNjcgtbWRjTU1yI1SweOYsykfJhIcCMVxtnTx9HUEMGBg3vQPZDGzdEMSuKlkswW+bqcJnNp0EzPBm4CKW8UixYrUDGjQMVUYhqlMZo0BwWo4LNsgQre3+JiAhWumTYZFVwrrE6zF6ggUMoXPSoaljTCbxO7gYAABbK5Ns8dt9lcB2yBgcgDGKCiJFyE/pv9CHOeK4uLoSYT6RyH09NJma8I1HLeLYoqE0IMq4OcUMgiSQprghvOxPSUALkhf0BkfcgU5LwuSQACJ8GgeDMUl/A4GXRe65SNINmQxcVx0fflpptzGpmDIo00kxT2G885Z4AKrnki/SQVZqYoACoDNTI8LBt7TZyXyDpDuTv2R6kBKvT9tAtUGIkjkTQcH5ONI++tMgKC6O/rlevhGmiBCju/yhMT8iMYDSEaIlBBuSg/+nr7ZczJ2mqknzTOmROPiuJiSlup9BOBCp6Paz4BHAtUsEhDmYTufJNIqNyB9fQSQIXnNFIX3jnEjSX5fFtJBJWhYCJDgQoFlxW4CGD09jgSySmwgICAN+8PQThHesTMRQpa8PsEKoYNo0Llx9QMlGkrF6iw85r0nyQ+8oEKFqbwPTIq5gMVXkZFvJzyaDHEA42/kfSTd++QD1Ysumos8sY9JtPzko/ud70J0fkn+hj597yv2OTnx16d7nQJd9giFDz+ohuaRU6y2Ofv9aJN8vpu12yBCoJcIp9iTZJNkpLzBOfg7ut9eO6nRyVBZl+/DVAha7eASK4WVCHpp+VNS/DoEw/JHHDqxAd45/X35PSLMUbn354vP/kEmlqWYXhoBL/+8YsYGbo9r0s+BlAhiWz92gOHDaNiJoEXf3oUPV298nfOkYuRUSVGKZiMdhn6+Y1SoEKSfDZdzsILU5XPii7vvkGSm6ZcXJ4bU9EvbTIHlrS7aaCtTi40Nu4UCyrI4XpzKlDhmvrqPXXHdWHwU+/dhu0b8egXH5N58divXsaZkx8ZXMAzB3hGmjtNmPftP7kcmld7GRVv4/XnXUbF1/7k61izaS06r3Tgh//H9504UsBpstwITMix9F5oYlzBBwEVzDUymf3Et76MnfvvE2bGX/7P/8kFsSRI1kPIfWDlPyVsTO+zmI7xAX+3bArxZzAsyEXHjSmCYntk30xTbJHGUVaAbT//RtlKttVK49i4XdYbE9PY/S3HgazjgYDJU5DRWiJrFdst+2djVMyfmUhWxonxNzBMD8lqcZ8uxV4u+4Pjgn9jV9h9mRfg4bVIW4zMD5PojG0oByreHRZn8ZLO/BqrsQ3BkO6FFTBRyS2V49JBIbK/clO5E9T4TsIRYTswJlU2BeM27n8tO4FxGBUi9Ha6M4mbm9L9R56MozHSVsDG+iyoybmMqnnztgIVCkjYPbwtlNB/uT81Y0eAygx++LeqrMDXV79Jicug4+dGmS7H2Jpjl/cop94VPA5jB87rFnCyUlNshwW+NCej8wPBXDtXyNg3DCN+j6wLAhXsP4mUjL+JbRv72XqC8PqU7aAeWlS00A6x/9h7RWaGYco4k522xYJVTn9b0It30fS19dsQsNQjavMpo6LQ7P7p336ne8ACFXZyv/vFeIEHM6E53Evvt/W9BUGKk+8375uHV4MPC4Z7mAqeQy4ar+ZhFIuDJvZQXqDCvW6vO9rCiNyDK3ha9BsAFSbJLzOLWaU/OaBCl5lC5t5ONFHoBi+2AfHMru6ic2eggsE8ExU0JhUz7bsAFVbuhqcSFkFxkS6yIumUEvSYnyFQQTmNWKxEAg0NLFwmB6WXFH1mAEYWwyyKipRRQSPVxNSMw6gI5QJS6VFW7zIqpNrPgBVmlZWFb3ZuWqu5jHa7ABVkVUiF5hxYzZgPVGjFusOoMJX7PKat9JSfJZjxmcQ75TfSwhRhEoMJHH62KBpxgIqZaVYUBkXTfjGgorS6QpF4k+AsKS6RQEWACn9IEmgiA+EFKoRRwSQHwQatNPHlaGZaKonT6ckJ3B4ddnwmWLnb398v5uFMOLHPGfDwdbN/EJcvtwlQ0dzcJIyKaFHEJKZ8ItFESREeoyiq2ud20+H+q2WAlDURsCYWEx1wa4RG3wgbfOmYyQcqtm7Zhvr6Wq0mJhAT9mtix+/HDIGK0VF99KSSYhZTk5OinT47OYbHH/+sXBsDwbr6ekMznsMvfv6sABWHHzwsQAXvHY9fXlGBIqnKodGtC1TYak8vHZWsg56ubmFUfO/b38EKASpc6SdKlZEFo54raZdRIUFPDm+89oZhVOxHVa1KP1lAwdUgZ7CbyWNUVFdWOUCFbhRMhZHPjxQDc39IfCbOnz2L5Mw09u3dK2PIAidagQTMZbO4evWK6Kwro4Kgl5rOK23FSD9duQICFZUVFRzwAhwyKUyvmPffPymyT63NzToLGR3+Y8eOYdWqVWhtbc1jVJw30k9kVLBPed+FURHw5wEVVy+3YcP6DaioqBDGi7BizOZ0PlBRKHhebM2z87I3WHfWEG9lzDzAbf7xCm2AXaAig7A/gOryCkRCNLbWDTqBCr8xZbPB7HywYjGggtIzClT4QZsYX2YON/u78M6JV7GypQ651DA6OzuxZt0WrNmwDXPZMALROPyBIviy1IT1rt3cdKgmKz2CMhlWLWXQ0dGG28ODWL16BSrKK+EjUOHPYaCnDWMEKkoq0NS6Cf2D47jadhrbdqxHLF6JdI6MgjC6rl1Eb/d5PPDAbkRLGpDxhdF28Sz6Oy7ggfu24sNzl5ALsXo9JWBnTc0SJBNBDN4cRl/vNcTjAZSXhrBt5xaUxqsxNpZGR0cfOruuYmSsHyXFMaxYsRorWlehtLgCPkTocEyxLWR8KdlUcy66fq0DU5MzIkvU3n4NU9MTaFxagzXrmtHSshRLly7F0MA4gv5i5AIRTCW5WQ7i7Kk30LIkhgMH9+LGzRT6R7MojZdIFTznRa5DyqggUDHrAhURlX5KJOhboUBFnBXwfj8mKZOUzsgaZxktsWKC4OpRQSB0Nsn1MB+o4HgjSMF5lWOCbIiGpY3wh7QCneBA0Mr1MIFDWQBupOcBFRyTnCuLAmE5RiQWFWkkCitYoCKR0E0X9Z05dxIw4BwwNnobwTDXNIIzCZHU46aUkosEKnh9E+MTMqfquqFzDNcPghJkMfDaOzuuy7rATWYsVuoBKgLCWGEinyAPN9oEKmZnEzI2mUwhUOGw2WTu0TVdPCq4Xot5domaSKZmZb4tKSo20k8BeBkVoaArpUAmCL8j3iM8bpaG5f0iPcW1ScygCZCYc0rMG/QjEAmiiNJPoSCC/oAAFYwNuC5bM23LYuS94332AhUEoZik5Gab5tRcCxWoMCafJn4kUMF7Z4EK61HhBSose8Gdm5hcUTkTowq1AKhQ4EKBipmZSRQTqJjHqPCCpxao4P0bJaMiRWkNHYMEKpi0IuRnGRVsC7/DIht56wAAIABJREFU/psPVLAghXEWEzm8z1PTkw6jwrJmLLhWXlkszI1Sf8NvAFTkC8D+qwIVeRuajwdy3GvO/rcGKu5W37TY4imbv0WuaTF2xKIXt1hSe7GTe/ao+Xo/eV+wQEWsOIpT75zBO2+edt5nlfNDn9mPNRtWyPP39qsncfb0Ref9TxqokBzvvP1yExkfTzycD1SYpOmdut2+99S/+zqqaqpw/sOLePlXrxb8isZHnrdcW0K3Ls8CFZR+2r9TZAtf+tlRdF9XoEJeizEkPECFHsaaNC82NsyxbGrBJDxF/s+TQvUCrgTSbbLduRhj2Gz71fv3O0mDLgpWkIVoIyOHzVpAwsyTz5BumQfSiE9AgZJHo13lGV9uvzrHsF1mcihs63ygwsuoKHTDee3WJ1CAYpEP0r7VmEOvSWRbPYbWX/jml7Bj3y7cujmIv/wf/5NzaKdq3Nb+G6BCsQ96jagHIvfXkriXIjzrI6FlXPNxLIHQU6wgV48qxlBSZc//sQbL7PvtWq9JZz2HvX86PjR5nmaCn/4a4q2kniKWkc7zqJR0ysgyzcqaI4WYZBtIexV8t+oIvHj+jcdmUpzH53XJHiVDCaeoI6lkk/u2YJFrlsb4rs8Gix1lrXXknPQ5kUeA12FqWkXGidX7hlEhgIDzGJmnyySxM1nGVurFyQIvBTQ0Ka8JeGVgsgiQ+QaRDBbQxfgkmDZaXw6nqj8cMbJD/JwxSqcfl5Ehts+lBUDy4oOcymVZFoW7f9G2i1Qn98C2MIseFT90PSqe/J76Q/B7jG2Yd2B8IoUQZImIZBKlu2gWrmxd9o/NMamMmftUiAG2GFPrMaxviv3Z3jubm1DAg14hxuvDeG965dLm7zftuDBTnzxvSoLRa+DLKUQzjB4qJ8yKAb32i4JxyooTJokjt6X3QNrlgLs5fApUFFzqPv3j73IP/MWfHDLNdyc6jTsKBxL67DhLtkm2K8JQ+DteKaL5PVUIVNBJutBr8aoNz6edry4EEdwtiWr+aeWSCxgojLlImwqxF7xMlEIeFVaayelhRUr1xAUYFZaoYj9vLnjR4Mmv9yh/q2XO8YkNShNYecaD7TdOsGqmTcNmI/00NycLCJMq04nEokAFJS8IRNgkK5srSRJ6VLAWwCTTrU8FgQommphAtx4Vklg32v62up8JIsZaAlTEwkgkJtF9/Tpm5gEV7LMKw6jws6qB0kyWUWE0CJnUT85N6SKquhZG9okJNJV+YoKIpo8EAajnzc+onAaZEFqlYZMEXqCCVeGMQJjsYaIhnWb1bLF4XVAmh+MyEg4JUMHFOzEzJcFRLBKUitkrl9vkXEuXN3mkn5R9IEEFpTBK4xIcso8YMLLvRApqVg22OLzE14MV70ZiiskcVnqJHngkgikCFTRBlcqUoFSXDg7eknaWlcdFYkmlmFjJO4iLFy6iuroGy5Ytc4AK9g0lUSToTKXEY2NggAbdqufuTbjaahB/wEo7qIQF/ToogSKmsbOzTmUHAyQafJ86dQoV5RXYunU76sioYKIo4BdTVBsQzKZzmOQ4Ms8tgTT+d2twAInJUXzuc38gHghnzpyRBOWq1askgPzFM78StszeA/vQ0tIq1bgMLouYHCmOif+DHfNMsDn32QQ0Yq4KP25c78LPfvwMvv3Nb2HtunUcznmMCjvmpco5q2CVVObMpfHWm29LWw7sP4Ca+kqpulVzLx1f/I5sLMioYABkpJ9qqqpw8MBeCVoZiJK5ahkVQrzO+jCXTuPiuXNIJmZw4MB+NWQ3xnUSSAmjAmi/ekXG3oH9e8UYmOwcL6Oip6dHJMko/SRG65QLI3CILFKzc8KoIIDV2tJs9pU5mT/IqFizZo0YZ9sX54azZ85JxX59fb0ao8/NSYKdM9KKNStk3iMjpu3SZWzeuEnmBTKS+J+MeZG6yt9Mzp9L3Q3vwgnTBp12M2bHjd3w2N/tN21Aa8/prfyzn/G+Z6WfWO1eVlyC4qJYYaBC2GvKqvAepyBwYSouOQcSJPKJBFQGmdQc2trO42rbKWxZ14DbI0PovN6JLdvvw6oNWzGZzCFSVAE/aOTMai3dmMnd9xHt4KbWulhkMTU1hnNnP0RtTYWAT6FwHNGwH303LmN05CbKymvQ1LoZA7cm0Xb5PezYsQHR0gpkUYzUbAg3Oi6it+c89u3djUisDsmMD1cvn0N/xyXUV8cxlZyDLxShaBgmp6YwPDSJTDqCJQ1LMTUzhOVLK3DrZi/27L0PkaJinD3XiatXu8WzoKYujnhpObZu2Y44z8l209WdDxwCyAUymE3Nouv6ddzs68f42Kj4nPT19qK0LIra+ko0NS/F8qZlWLq0CR3tvagsb0AgVITJxJzMmx+9/xpWNZVi7949uHEzh4HRLGI09TXrgDL7MsLIIljPeKMoEhXpJ96b6emEyCQS6Kb0E4/Jv/E5jhUpiMvnmUk0VouTRcE1lWwCDmkyt/iyJuxMdHNO4rgfunULjcuWIhBR1lqIYIVUg2UEoOdznzIbOGd98DAqikNRDN66hXA0LOwyX5AgypT6NUxOOx4VlF2jhAHnExpOS7W9ASriJZRYCiAxTY8KAhUBkTkkKEE2nq1yI1AhoERxVI5/vbNLxi0ThWRUiPlkhokKehHQdD6GmemkPOtMYHOdZT85jAqPmbbeb0iSn9/PAyrSWuhQHI2J9BPXCPqUEJCJFkcQEUaexoK8NvXNUDPt1FxGigUILBGQoTyRrKcEKjKmspSMikhIgOxokAxCYKD/lrAtWcFpGTESK8zNCUCmwESxgN79/TflGvkf7xHjHyv9pNWHKr/ANjJ+4Mvef+tRoYUbKrPgLU6wRUEEKnQiNnJzBtiRdceYXlI+a3R0HNMzkyiNxxAO20SDu8G2CS6d21S2gYwKXhvvdzBIfxBlVJAVy/PbRAa/Y9dMenpRYqwoGpPYIBgMi7kppbcsUMH7ZAEKHoPXGC8rkgKXOM20Q2GEwhH5HtcxR5LLVH165+q7hsgfDztwD/OJJeAXP/G/OFDBqzFJxoV7o7v2WP4H7gQ83NOhFukPWw1e8Fiuv57ztm5cnF8FqPjcIZl75gMV/FB9Yw0e/+IjKCsvxfmPLuOVX7/pHqoAS8DBdAooVVlVZO+VOMPF209OMjqH5c1L8JgDVHyId94go8JNJs+/7PnD70kBKioFqDj6q2PycWev6CS7bXzkFgdKXZYZB95zPPCQB6h45mV0i0eFed0FqJC0sbOf9bATFlyE+56TqDW5Bfm+cx4D6xi/RO9hnDs8L/bzfsZ2szemWnSfXZARokezMjILL6NwDmMxRof1H8jDjMx126r5/PbrTWpZ3YonvvUlkaM9/vJbwqiwDAf31rijzrlG6UsLMJn3lWLtnEaAZwMskVFBoMLLqJBErlSvq4ST7ImpImCq/PmsMf60j102rTGsshJ1/dAiQHNKk8DlZ5hTsNK23Mvan0UWTOSfXABB9j7OeF3Y75IbNmbKNsnsHUqS5Db7f5HwoZyQSdpLy0y6i32hVew5ATPIhFQ5Q78B5aMm8a1ggjxvxhBc12zNDYiPpInnGeeo94UWbri5r3yzdybghRFg8kbyfZFJUokkZVLoS/YFUl6ieRT2l8gkGXlplXbUGELmesse4H7NyK7Z/QbXW2HEeKRm7XOsAJEm3C0gImOA12ikofRcrgE7z8k2CWAjfhZZWatFStKY1Vswi4374d+5eTKaafNz7j5Lx44t2JMDGr8aC7LpZwnApA0oo0CMY0wufiXcP2s/iWyySFApIGLXQPnZyIdZRQpbCGL3g84+0TPJW58z+x6vnfdCjmfGpP0bx7n0iwHdOBbFb9KR2lKvUwIwLCyVwkM+owQqsupXIayjT6Wf5k/Hn/7+u94Df/EnBz2X4E7yHwcUcD9jg4ZCveFWpi18tzAo4JI2f4PenQ9UyCJjQBgHAFE5FrtCqs6kJwhaIP/Ea5gXLBf4TF4g4QA6HlktsyHUYMtbH6JttNUM+TJW3uDMPYOc3gAVsiCaighdqOznCgdL99KrbvBtgxkDYglyr4lGJvRT/I8eFXOzHwuoYNLFghA2eGNig3rVXqBCpJ/SuoHlppkmrUzS2IpvS+lUoILmUPSoUKCC1aisBOzu6sTMZD6jgv1V2dggHhU+SSRQGkflcazZclbYCNOq++9TNJ5BCSmA6lFBb4IpYVQwicCKTr5PqYbUXEICGQtUyBpqfCrYkwyEuIBScoSJBlbNM8lFAGB6UsERSmJkKCNF74jkjAzjkqKwJIuZnOU1LG1qFlBBPSoUqOCLixy1wLkASyDkD0lFqoA7hvLJz9Egi0Nnbo4m0mSCpODL5jQpEi3C1MSESD9xoeXCzITJ4OCgAhWsmg0w+DJARf8ALghQUYtly5aKwSUrQpngIVBhX2xDMpnG9etdcjwey1bHaABJnwWezw2+eH4mbSSJYl5c4JnkYJLu5MmTYqa9fdsOB6jg9yNRNeCUPslA5Eos/ZQG2Ewk0vMjOT2KI0eO4MaNGzhx4oRc/7q1ayVx9NJLxwSo2H/wgJg+89mjjBWTjzGRiaI3Cq8pKeeyiRQFb5WMwzmtq+M6nvnJz/Hk17+B9evXU53J8ajwPgsy5qUUXg3TWIH9tgAVPgNUVEmgUsijggkh3QUE8OILR1FVUYmDBx4Q6ScbrFqgQoNSyqCQUXEGc8kkDh48YDYcHMNaPW2lnyxQsX+fAhVW+knIuj4f5gMVmvBSLXyCbydPvoMVrS0i/yRaw8bY96WXXpJ+pR+FfRGoOHfmnHha1NbXa6Itk0Hn9esSZFLyxwIVly9cwqaNG43WuVZs20BY58N7zThpK+4EVOQBDuazdmxK8LgIyyKv4ou3yZ9DIAeUFsXEF0aSnR5GhWzaPPJP3mfItnE+gCFy89aLU35RI11htZx8DeOj17Fn1xZcvngB7Z3tOPzIZ7FsxVpMJTKIRMsR8BUhl2U1EpE0Tnqkj5N6rhscHc0ZtF0+h9HRW1i7ZhWCoRh82TSmJvowcXsIZZV1aF6xGQNDBJLew47tG1BE0MBXgtlEAD1dl3Gz7yL2770fwUgFJpMpdHVeQWZqCEXETkNRJNJqFCwJ4Yp6zM0GMXBzEPFSP9ata8R7757Avv274Q+GceKdcxganBLgtqauHN3d/Xjk4SPiH6SUd60ok02IPyeJ97YrlzB+ewxjo8O4fOmSzLHNKxrUvLuxUTwt6mqb0H61GzXVS+AnUDHDCv4sPnr/GNavrMSePbtxvS+LW+M+RGIhlYSjRwWBikxWmBPUJKbnjBhtG6CCXg8EPKcTM8KoYMPop8FxTqBCKxpzsoZRDtECFfRn4LV4gQqOA86BYrZNoGJoCEsIVIRDMp5oABkNKahJoILPfYqsw0zaAbI5b9k5mNJPBCpCkZCsD75QQI7P73uBisRMIg+oCBOo4Nw+m1QANxRU6adMWhgF7HNuzAlU8MXjMZFNsKOoKCJz3XU+31nIsyxARTaNbJrgEIGKOIpixUgYoIJ+EhkBHNTgU6Sf8uZfA1SMjDgb6VgxpcRUU1j7OoZIMCqbPPqGTExOICpm2kYykECFGIX78oCKgYGbwhC0BRKcW3UDT9ZODj5K7YWDiBqgglAAGYece1kwYNck8dlKpTA5ZYGIGGZmptHX1y9rkI112AZrpn0noILHt4wK9j/HEMehFJU4utDGvNGnSRc+H1pAYz0qVPpJi2sDGB9zgYpQ2CZLPF5lefOTJiYsUMF4zjIqeB7xDTEeFXZus4yKXI4SV2Pi9UWggs8uv2uBCgU9dJzascprpEeFAhWNAhoVAiqsPIUTGS+2wfEGx/e6bPwrABWLFXEVXuJc3fuPHfMbkIKflz2F+BPcK6PBnO0TAyoWaf0dj//bAxU865P/9iua7F8EqNj1wDZs2bFe2HR8/lmZTcPqt185ickJjeNlndbHAus2rcauPVtRUcW5ShNNk+NTOPvBRZw68ZF8VgGKhzTGcgas/nD+w0t4+dnC7Ag7/L785BewvGXZgk6jbOqLP38ZPZ2WCZHDrn07sGXXJlm3BDzOZDA6PIpTxz/A5TMshnJf+UDFUQeo2LJrM/Y+/ICwp2mw/dIzR51r5y1qXtWEBx7cg9qGGnl+OVcPDwzj+CsncL29K7+dkkowe3OPrwT/RGblQ597CCvWrhBGH18suurt6sW7r72L/u7+vO769n/8DiqqKvDBidOobazDkqYlTuX3YP8gjh99S2SR5P7k/x92H96DrXu2I14e1/s6O4eOy9fErHpyfMK9rwYMaV27AvuPHETdknpj1pzF2O1RfHD8FE6//b7zee6ZN+3ajEe/9Fn529FnXsD5U2dVZsmkqbft2YFdB+4XNowdI+NjE3j/rZM4+fo7ZkApY0GAim/STDuGE68Yjwpztif//XfQsqZVrvEf/urvPNeZQ8uaFXjk80ekvSHZv+QwPTGFc6fP4vXnjonXEQstnnhSJZ/mvybGJvDj/+ef0HWFUo2aJdi+Zwf2PnoANVIopmOb8dV7b7yL18XkW2VrBKTmCsOks+WcGDTDKb4xz7Ywabj3NDJDUl1ujs1zyrpGGUICAdIKb87D+BIYloDG55pnsVJJPBYLSfhifKYJapVtsjE81ycr42SXBMYx3KMI+CCFADQHD0kMw3WWbELun/OK8EySmW1ljGTBGD4PBCpsQaNeen7exx9SU27bbhmuxsNCCwCUcS6AhY9tSGstrJPA0c/r3kBHmjBrzH7anjsaow8CfRLnHEaHBXIk2W4Myslqt0AFj2dVDhiz2J9FDonxmBTI5Xta6X3QdvD+Kbiha7tl/XCEP/0PrkfF177F+2TNuAlkhU1Bmvo4yL0rkPIS2TAxFXeT/vxd5Zzoc6HG2RJXmHFmk2gyBgxjg3+T/ZmRSbPDTU3iNS8hT/G8NZS5RgFwhLWjeSZh+Bo2B3M08t0cATCyQbjf0nFq/S8o3SW+HdmMwxzS+TotOStQQlqKcVKfAhULZqtP//A73wN//j0FKvJBh0VsDpwkuAcCN9+9Uy6ID1jh178wUJFXvpJXq5CvJ2lYFXYSXjjbaV3BglferJg/QzKJ6V0ztRrETs7uguoFJWTiNofJZ0ksdmrz+bzveBkVnzBQYbEKaafS7VxGBSVr5j4WUNG0ZpMkVSzYYDfQnHjnMyqkWpwazWOjUo1H1gI371b6icewHhX5QMUcYsVhB6iYnph2pZ+yatBcuaQRFUvqiRoYRoUmdbiQyHlFS3JW5HSY5JJAi0CGGGoGkc6mJIHDDTWDGSbKrQnU3CyrWymnpNWMfNkKSPmZ0kTwi/QTgQpWkWryvwzjo2MSANFIk0AFE8Y8Hheu0ljEBSp8fixrapLEljXT5iad32WfsLLSqZj1cUNfZiS1mPjRsSFAhZ8BvwUq0uJREWV1Z7QI05OTGBm5LZ/XpMGESKYoqBJn1zlABatAL5x3gYrKynLZXDA5xGpxSzvVIEzplj29vSozEonI8cmCICgoj6SpOLDnttUbNlmhCzu16RMCLtBMe+eOXXmMCgIVtno1m/MLA4bnkcB8iv4gsxgaHsL0xG0cOnQQfb19ePOtN6XfRDYlHEFPdz/Kyirw8JGHsWrVaoQiYUk+ssqTWTUyKnQKUTDHtk/3XDkwvyuMis7r+Ok//0yACppHg9WpYhymlGQBKCw7wqeapRz7yZkkXn/tDQGkDh08iJr6KglEed3qD6JVqQy65wMV9KiwQAUrV7weFQQQXOmnc0jNJqUPbBUN6adCxWUFdiaHq1faRBpr//59KIsTqDDVuoaZZoEKkX6q5LPApCgDT1b0pwWooD8FWRLsGyZM2XYyKqyZtp3pyCI5e+asMdOudSqDCSQxWFu5ZqWarE9Ng0DFxg0bBMhi/xFEamhocBJ2nxRQMR+4sBsZ7/GlWsejXWyfM3tdeW1h4M+q5kwWsXAE5TSmpna9ASoChnpfCKiwST4b4Hr/FRaLSAwQoNDKIMrvcO4aGxvC228eRWnMj11b1uDkO2+jvasLf/iVr6GyrhFzKR+KohUI+MiYCZlAgDq9NOO0QAURFsoXjePUqeNYuqQW7e3XMTM5gl0712JmYgzxqno0r9wqQMWVi6ewY5sLVFD6qfv6ZfR0ncXGjSswMpbAVDKNirIilIVziIZyiBaXIuULIZvxIVZMgDWC8+c7cPnCBaxZ34hVK2rw8ksvYM8D9yFeXoW2tj6Mj+UQjRVLMnxoeBwPP/yImUtUdsDeC26PKd1Dv5PkzBQGB/pwvbMTlZVlqKsnqyWBquo6rFy5ATVVS3HtWi+qa5bBHwhjYjoh5s4fvv8Ktqyrxf3378bVrjncngkjUhREPE5GDyWLtFqMsgWcK/gURSNFiEVispERRsXcrLAOy0pp5prD2NiEvFdUpJX7fMVinD/pU5CRsc5EmNdMm8lrvjivEYTlekjPncalS+EP68avEFAxl+YzrUbaumFygYrSSAwDg4MIhinLFBUvHR6bz9bk5LSMI3pUJBNJkWdgEofsBhpQM07iukfpLfoyJMkm4UY8GMTEpMr3sH9sJSDnLa4RAlTkIMwWNWlUoELXTwKmPvkegWNKPzGpMDY+pj5QUhGXRhkNvGUN0bWFfggc+5ZRQcCfa5HIFRqggutSOBCRjSNBpQnKEhaHERY5AI3XeO18cRMuOsXpHPr7+wSooJk2/6Ya0LKya8IpEpD+i4ZDwqhgv9C0XddlBSrsXMH1fWKSCfqouT4FKqzXBO8P1131rOA6qtXPNp6gFAv/RqCcx1fmB5mIus6pUbYWL9g5TCodPUCF7pTzPSoKARVhynt5imL4NcvWsImHOwEVIj/hASr4Xa7P/I+a1PTiUKCiCJGwJiMnpyYxPa1sHFajqnyExiPKqIjJM1IaaPg9ASoW2S7d4c+LAhUyGO8RcbGMCquR6WRx73E/8S8OVMigLdArNtE97y1b2m3+fDdGxdqNK/Hgo/skAfnBybM4/pp6ROhZc3js8w9i3aZVOv9OzUisFi/XuW1oYBjPP3MMoyPqy8at4padG7DvwftlHNM8l0VKxSUxSbpzjT//4WW8+sJbqG+sxb6H7kdxSTHKKxhjBzA+OiHzdPvlDrz7hpv49l6hvc0Pf+4wGpbWS5Kd56Jc6myCfmwzePvYOxjoG5SvfeaLR7Bu8xr5eWJsUpJ1pWWlEotzLnnzpeO48IErd1UIqGhZ3YxHPv8QSuIlctyjP38ZI7dGnGZt3rUZ+4/slXWCye/pyWn5LM9BoPvNl97C+Q8uuJdhC/zMvdJ9s1YRf+Ebf4imFU2SLGWinH1WVlEm88Dtkdt45Rev4EbHDTkWD0Ogoqq2ylnf6FPIF5nQLEwj4PDSMy+is63DABU6lh7/2ufER4KvKfpGpVIoqyiXoiICHL/6x5/jtvH74J5s+wM7cOizD8n8zX5j28j+5nmYhH3/zXfx5guvy/HY5k27thQAKnRUHX78IQFJOM9Njk8iMT0j96SoOCYFayeOHccbL75mB6EAFZRlskCFeFSYZ+LJP/uOvH/9Sif+4a8VqOCeYvX61fj815+Q8cG1m2ACx2Ap5VxzOVw934Z/+i8/kM8f/OyD2LB9k1wL+5r3kEAW94VHf/4ibt7ol0TvrgO78diXPgsmunlfJ0bHpd1kenCOP/XWe/jlD37u5s1NAY7xaTcqE8YYWpgaGrNJUZ/xtLA3lkPC7v91fGgRoAs22eHkZm1sTG7jZrsO2mp8/m5/Vi8C9XHUwoISua9WDos5D22fgiZpJsGN0TTXNnl+DMuRx5CiKQmZVZZImBOm0JPrl+QHci7rwDIcnYeCLJSQ6Q8BCowngYBkmvi24IqVYCKLnawKiTNA1qXKS3EuE1BCCAymiNiwJbivcuMDY1Zv/SZMYZlNyPOY3B9KrEUmhlHUUB8IPa4wPmjybIAMtoX3LRSkxK0aZ0ufU85JFDVCTpEof+ce9+nv27gKIFDB4ytLRFEYjl8WZ3KfKjElczXzihAY/ogslNxTle2yCU/xIGEvOkbm1hNQe19jFb034uNlgAsLQAlzJJU2fhhUNdA5xCvXxn0u8wgcz6qCoL4hPJ4FwRxghN4xxl9H8xthke4OUtHDSlUZJi2PIXkKgr+szmUxGvc5nzIq3PXk059+P3rAAhXyUObFoYVT5fmai4UC1/mBoyKghV/3ClQsFnB72uH8qAvYAtqk4btJxZhJsOnEpptSCyjMb2/BEP1uQIW7Xpo11tVQlMh1/kHz8R/zncKbAwFCeIHytj3WfH+Ke9xYFLhJGvx6ARZT8GIWGgUqdIJkZX0ylbwLo2IGLeu2SmLFBhuWZsiFhhV4WhHACmqVdOBCoMkGbkrLRMeZrAC+Jz4WmbQkDHSRZkCgiTn1qJgS6ScGVqVlZVLNGRSJAz9qli1FZWM9clxsufEVaqUusjynJEFAQ1suZjqGKfMkyD8X2EwKk9PTYtLKBYvJWZuAoXZ2ao5MiYzS8XhGcx4eJxBi8kI9Kig/RD1tJtrLCVSMjcqtJRuBptwMDtNyrDTixVEFKi4ro2J5U4tomjcbRgWDJKnySM1JwoLnZ7KMCQKVpgJSc7PGdI4SGxGpvJidS6rcz1xKFn2p3oxGJTk2MkxGhYI0TNrcujUooEe8tESkIET6KcvkzQDOnzuPmhoyKpahqrZSwBYeh0l29oOVPQsEVD+Sw2tyagI9N3ok8CGLRHIoIpekVSCsgLXVH3xG2Q4GeBLYMBmWnMXx42+jvKwCu3btRG2tK/3EwIzJMd5bHo9JHams8PmkcpULPSuQp8aHxEi6p7sXbx8/LuOKgSgrzIZujaCmpg6PPfYYmlqapW8YBhJsm5lmcpBVzhlJglEuywUqtF5ITKNzPgEqfvyjn+LJb3wTa9eukWSWpQSryZmOdUkoidYrfVrSGB8dx8svH0NNdTUeevBBVNZUSDI2wqVPAAAgAElEQVSQSb3bI6MIhgJYumwZSrgpoEan0EcDeP7ZF1BdVSVSTTQkzgcqCCKwR7SK7uL588KoOEygwlQQOUAFWTiZrAAVfeJRsR/xslKRCJM2MiA1jIq2K1ewc8d2Be0Mo4L3nWbaBCoo++RIPxn699GjLwujQpgW5iXSTx+eQXNLM2pqa+Sv7JuuG93SpytWW+mnBC6fv4CNGzeKGS2Bm+tdXVjR2iqSURoQMjVtXvOC2DuBGPY9CboNO8YCUjYY1rVN+8EG/l62RSGgwllnGDwjLXkk+lQQqOBmV4J4VuGQMi1Ag6kWMhVI/ACDWRss21yN0p3Vn0Leo7eEfFcDY21nDtc6ruDS2ZNY3VSN5Utq8eobr+HW6CQeevQzqK6vgw9kU1UrWCHJS1ENdiqvJTIQTVR6VVxGf98N1NdXY2ioD6taG9DX3Y2auiVoWbVNzLTbLn6E7dvoURFHKhtFejaAgd5O3OxvQ01tCYpLq1BSXg36AsSDaSSnb+NKexeCRaVYvWYjItFSjNxO4tzZKyI3tfeBdVi9ugFHX3wJmzevQePS5ZicCuL8+R7cHp9CfU0Vysrr5BnTe2j6wAyCdBYiUdbX14PZxDSGB/sxOjqM+voaNDfVAP5ZJJMZrFi5DlVVy3DtWg9qa5fCF4hgbGoG2eysABXb1i/Bzp27cOV6EmPJCKKxkLDYWJ1K1gPlCTj3ckzyuZREdITSTzlM00x7bg6UQCwvoyRfDmOjYzIvEdCwOs40mWYSn+AEQXHOBzy2Gr1yjYgpYDc9LUAA5+Lbo7exhECF8ekhUBEx9Hp5Zpm0pvlkes4BKsSY0EgElESLMTB4U+YBYbGJ0feEzBNcr6yhITfjTHBwLabhccRIP/F3rg0yN88QYM/IsVgZL0yJkhKZizj3cs1WmaeYA1QwluBmNlZcYjaIKqNAVhuvNzEzKzGASD+lVRqRcydjA7fiXmV/2EcWqOD6xmPKhplm2tmMAOiswqe0Y2KWptaTKIpFRMZKkh85iGQVH1L1h2DVJGQetEAFr4WbRVn7qZHHzW0oINJPBCoioZBED319NwVoIshvzTD5TPKeTUxYoCImLE0CFRZw0PcnJGGiQIUmGezaYYEKjjOuWQJwELAJ2mSDzhXCpDMxrgtUaOyr9fOuZ5SVfiLrUxgV05MoiRME1D71vrzJH52LjPRTWqWfRM+bmlhSxakAjZ0X7Rjg5xhnuUBFVMAKPisEKmZmlI3jZVRoUUAApSL9FEWp//eFUVF4t3Snv35iQIXVRNFiV8PONDd8se3EnXCQgu8V0Pa/90v2lsHP+/ZvD1QQVNhx/2YBCoYGR/DCL45hZGjUOc+uB7Zi94Gd8iwKiPH6+9JdG7euxf6HdksB0Jn3z+PNl7UCnjHgN773ZdQ11Ii3wy9/8hJSsykZ049/8WG0rGrC1OQ0jv7yNdwQ74ccmlqW4tEvPCQg3KnjH+Kd10+aVbxwZ91J+sl6VNj9++YdG3HgyD55fk6/8yGOH3tXDlpdW4E/+K8eR3VtFW50duNnf/8L52TzgQoCKA9/7kHEy9hHQ3j+Jy/mgRQNyxrw+Fc+g3hFHN0d3Xj2R7+WxGJlTRUe+9IRNCypR++NPjzzDz93jZDnAxVm77lr/y5hbXBP+NbRt3Dm5Bnpo407NuHgZw4KcH7+9Hm89MxL0l4LVFTXVsva+M4rJ3Dm3Y/k79v2bcfeR/bLfN5zvRtP/1//6AAVBAn2Htkvs+H7b76Ht156Q463+b4tOPTZBxEpiuD08VN47TmV0mpc3og//PoTKKssx41rXXjuR78SACQSDuPRLz+O9ds2CNjw/D8/K4yMxYAKjtimVS1yLAI550+fw7NP/0LGeCgSwVe/+zW0rGrBrYEh/O1//huJp/laAFS88KqD3X3rz769AKjgXP1H//U3sHbTOpFx+vH/+yPc6h+QY/3h17+EbXu2yzrxwk+ew7mTH6kmfzaLL377K9ix15V+ktSD8THgHP3v/qf/Fo3Ll6Cz7Rp+8H/+vexZCU597Xtfx9rN6wW8+fHfPI2OS9fmLR6apM5bT4ycjTeOtkb34sFnDJltQQL3BTYWdtQ4LENF1hq3UMUC97YIgee1a7EqIKiHhsoWqkeGBS1kZbN+CIZ9RJAgZXwsuLZr1b6ZPH26Z/Gud/xZkvVGMtNN/FOqOCDvaSGfF4JltooMR5NUp++HieVtjCL7TEl80zMxI/GmSGSZPXdA4hZlsah6h/a4LabToEKLDiTGIcvAMCL4LLA/pKjOSFkpsKOFIN6X3SvxbzyWt3BLr09loeznBPxhnkdoCq5ah/oppvHPP1SFCL7+zVMqAcq4mUwD9q0WZJClRaaBelTIdXn2bJrwD2GO12BykTYOYl+J5JMx4HakpYxfiJQYyj1XLxeJYRzWhSvtxfiWYE1eTs90Db/FNtqCINsv0tcij6weKnzx/gjoYPatUpRLtokB4vgcMF6VvJuRrLJMHi3qyX4KVMybTz799fegB/78ewfy6HJ3Z0TnR6vezy+W9OFmp/DrXweosLNHPoZhgQqV89H51qDVtrF5QMRCAMYu1u6U717lfBMtXRE8fWd/9nan9xR52MvCHYIAFVLib89pPiPn8QJDvx1YQY3JBUCF2WfIIi5SS2oALIyKxYCK6WnR4ybNsnX9NkxNT0lwaimHNihhct4m+5VuqbRCJhuYAGBlCysbmSQREMMg+RWVlSoxIFTQtCx+nORnEwmRfmLFfFm8XP7zBULI+QOoaWhETWO9mAFbOQG7+RdJhnQK6YxqYKumIymWXBh1w8xED5PkPoRkU02DYeaI01KpOissBW+Qo0GMBiE8BpMB3ISzkjObC6C0uBwVlVWYmByWexuLRKXKnZItBCxI8yspLcbgzT5cuXRJJJqamloQKSpFy4qVKK0pQyisFf2soLDVtqwGCfhoRkrJjZwaZktlAIEKlWbgIirgD2mrNB0tLpF+FumnkREJSPg5JsvIqCDzg6agBBb4Pfb7rYFb+PD0adTV1qG5pQXxqnJJSlEaicfTvmDylCQWrZQQ+qL0dRpDw8OaVOL7fg1A7DPpTQJLlbBJDEllVmIGZ8+elaTIzl0q/WQrVm21pup1UzM+YWS3/OJvIFVSgwNIzU2IITOBio/OnMXMtEqszM6mxEB66dJleOThhwUQ4qaIwQqvmdJio2O3MXp7VDZsBAaYoLcBpA2M+NmeG9340dM/wrefegqr1qwWgIH3gC9LLdb+55jiXKSAAxNzL774oiTzDh8+iIpKlU6ZGB+XapKArbCR1LShQeeCeO7Z51FTVY1DB7khVaCJCU+t6FEDLjIqCPRdPHtOgDXLqLCJLWkPAaxMFm1kVPT1C1DB+y9VJkx4ko7q96O3p0cAtJ07d6JS2EVMEVP3lIyKFN599x20eD0qTFXR0aNHBWgguGVfc7MpnPnwQzS3LJcEMscBfVw6O5VRsXrdKpG3ol5928WL2Lx5kyR051IJXOu4juXLl6OZnheSs3DFBBWc8czTnt8LBd3uJ21Cz8z2Vk7QAN8cW94xqoCaAtNesGL+OQhICGzqg8jlxOOlkthjvwd8WmWcEVYXtXO5GWGikIk/j7yTiY4VqFCfEgUEta0EwWQfIGALQY4Mzn1wHP3dl7Bl/SoBRN94613MptPYc2AXamoaEQrEEYlWAAECJ6z64ljhd0kpN9RyAUTTePONN9HcVIHy8igC/iw62tvR0LAcK1duxq2hcVy6cB6bNq9CuMiPsYlpTI6RQZZGTQ2vtxiRaCUyuQiGBm6ir+MiouEcrnf3YP3mrVjRshZZxNB/awKXLrXhZl8H9u5ej2WN1XjhxWNYvaJBjNV7b6XQ0TONxMwMkJnG3j2HDDCrpoh2Fcz5fJiYTuLMRx9gdmYC0+NDmBgbgs+fRn1DHbZs3oju7m4kkhm0rliLeFkNOjt7UdewDFlfCGM0rM4mRPpp54YV2LRpG9r7EhhNhkQGrqy8TKSf7PNsDY55P1XKp0j6khJOXDuYlKbEB58lJqM5H1EyQCrGyTAspk8BN8yaMOd8xO8zEcbngJWW/CyTMZzzOT/zcw1LlsBnqt04l0a55imKhQyy8swSELWMO64DfJ//FkWKcbO/X9ZPVvVyQ8oEMt8fn6B0XlCS+cmZGbmmubkkxglUBNnLlH6imbYaW5NRwRfne/ob8fgEzGXjODdn5NponF0i96jrepdUkBXTI4m+RmJoyQ0mQZkS8S8g+EOmB5lTqZSusXzO2fe6Ceb8axP5fgwP02NJDRZp0K2VfSkZy0wCMvnOvyWTcxgbnURxcRQs+uN3GEvxPBzznF+ETekPC7NsYnxSAFtumuW8xmib94MbT0pn0RuISSu2v693QJ4XMirsZp19xPl+fGJUWCIEuzkmenv7lBFGpkeS93US5eXlDnOOfaqJIsgcyOMpUJGWe8IEqG7WueYqUGFjLbvuyo0RdZ/CxUS2cpHjkuOKVcI8rs5pesz5lapWPmp4eETiJ+sRxXYIGGLMH+2cKPMcgbQIpb8ywpwlo4IJFwJ2HLK8dhYz8DmwjBmboGCytLQiKvcm7lvy+8OoWBQUKPxG4b1XTskU98KoKLQBNEmkBYVVzj7pDhvh3wGgojRORtvCF/u0r2cAx154C7c9IAU/+dWnvoAly+rR2X4Dv/jnF+yjJP9+5omHsXbDStwaGMY//c3P5G/cRj31p191ZKSO/voN57asWN2E+/ftkM+999YHcky+SQkoF6j4AO+8royORcv15r3h9ah45Vmtwrf7Uso9bdq2QSrFCVIoy0KThUe+8BA2bd+IkaERfP+v/tHpGC9Q8frzb2DP4ftRU1cj680rvzqG61fzZZwOPnYA2/dsExmoX//4eQz0akKcw2nr/Ztx4NH9Mifxu1fOXzWBlX5ACwxduYa9D+3F/QfvF1bICz99QYAPuZpcDkeeeFQAA0o/vfKLl532klFBoOLCBxfw0k/1Hun5s3j4iSPYev82Od5LP3sB7Zfa5bzf+PdPYmnTUly73I6f/d1P3O8gh89//QtYv3UDBvsG8Pf/+9/Ke4c+cxj3HdotgPyvDRghzQYEkPnKd/9ImAjvvnYCb7/0xqJABb+zYv1q7DuyX4779tE30X7xqlM9yvPsfXifMHd++cNncP1qp3yOZtpe6SfxqDAvB6i46jIqmKx+8j98B61rVijT4i//VtZYvpY0LcMjXziCaKwIH544jfdef9f4P+Xwpae+IhJQ1qNCk8osJFT2+3/3v/4PqGmoxenj7+OZ75t+8wFrN67D4T94WI5PcOfK2cvufVaagZvsNiCpyGAZsMImui1Qwa0O13YrL2SNmaXq3cT6JpVj4QIZSVynbDzOMSOSP4YxYedOnsuCFoyl7FrD/ZJNdDMm48vmKFQWSKXEJSEeDEmeg2u57H9EbklNry27QJgExgzaPs38iE24657FjFUdsSoF7MlPKcCgz4es08xhiXm5Mh7phUVJTcs+kcIXkUDSfQr3AeZhcPZxEnN6jKXJdGBBjPgspG0yXcEPMRH3SElKPxj5b7v3tXsifYwtGKCMBSttqvGD7pPEu8QU3fLamEP52dPKGObrj55ULy7GUHr/cojQ3NtcE/Mj0tdGMs7GGDwWr9/GmzanJMCLg8UriCPG8iZ+5Ln4Wd43mZMclpfKcNn7aQEWWxSdt9+zM5kBziygJqodprhNgZSgY8gukszi8aG+XioNpv3N54CxEvcAAraZ9glIIsbbnwIVzoD59Iffnx748+/udxIa8zkUtqhGp0qtuXIq+GXSdINmXRwKhVC2eqpQgF0YqLDnkwnOG5h5ki/uKmTa5AUCzJ84GcvkYSZ0712jZrSZ6Z3r0Gs0SX4ew3hKaBvs6pEPNrh9kH99MiH5mCBxj6cLwzzmhvdwklCTE3vAI/O3+Z0h5Al12vD6U2iHzWewOGkaaYK3T72iVvl/N71lFjTvrTVxjZF+MlXVAlTMIkkGgJhpT2M6kZRFm0kU+Y9moEkFKqyetk3kW1YFk+sWcLAgBD8jiRK/T5gTTGAwkGAfe4EK1Q/kgpNBNk2pjQhmZxK4IUDFCMrjFaJjzcSbABVLlqCmoUH1LU1iwwIWwoTIpCXxWQioEMpfJo3k7KwYtTJxwrYxThCAI5WUBITQV80iZ5PnsnD6WcGaE8BmZkaBirJ4FcorKjExMSSb9mIyR5IJZIz0E8EgGvsN3OxD24ULClQ0tyJaVIrWlatQWl0mchNeoILjk/eDY7k0bhkV6j3A67ZGliIBYozJ+TMTJlwQpycmMXr7dh5QQakmskd4r1iVxOoZPku3Bm/hw1OnhNHQ1NyM8uoqSXQxuWHZHHJvPAu0BSpsZQn7g9VZlGXSaltKgmigZweuBFTGjMsCS6ptnpaEdW1djSP/YSWlRK+b1ryz6iPBYyid1y/tTqcnsHLlSvT33sTFS5cxPcX7pxXRZC40NjbiyCOPoLK6WjRYBSAQw7UUxkZHJMHG5FRdvWrUsl9EIdrkizkGerpuCFDxne98R4y6AyGOO9dkTemlBBLmRLLHLzIiQczNpsFkPhM1hw7tR1V1pSMT5VSOCGhA4DCjFb0ICVBRW13tMCqkMsSYaYs6rDA9NBC6REbFbEKkpaz3hX0mOX5YNUQQgvd+3759Ut2rVR1Zco6kP3t7euUzlH6qriRgwwoXPQ/NtN9/7100ifSTMdO+K1DxAZpbmqRan0HZ7GwanZ3KqFi1dqULVFyiR8UGSValMrNob+9AbV0dWpubVcvfUGklkPuEgAobfJto3wS4hvJsae0fA6jgsJZEIXIojtHnplRkZDj3BBBGNsfgm3OIgrac27mu0TxNHwplh6nUk2V+sEpNq3I02NaNqMyNZgGYnRrHu28eQzoxiR3b1sPvz+GNt98CR92u3btRXVOHYDCGcFEc8EXhQ1gev3RmDtPTE/IsxUvL4PMFce1aB250XcD27eswNzsppvHLljehuXkN+vuHcbXtCqpr48j5UogUlaC6ogGxIvr6KKiczhZhLhPCR6dPYfJWD+pqSjE8NopN27ZhSeNyTM/60X9zTPxvopEMGmtjWLNiOd546zTixTls2rwB7d0T6B8mmBIQ8OHRI5+Fn/JJ5l7Y+0TwsXdgEFfaLmIuOY7k1DBmkxOoqIxj46YNsvE5e/YCotE41q7bhKJYGbpuDKC+fhlS8AtQkU1P48ypV7Fny1qs27AZbT1TGE+GxYenorxcng2vh5LKs9FXIixABTc5BKc5tzABTLkoB6gQ+UMF6znmCSJR+5sAI6v9ORfosSIincakAp89Hseus/wcpZ98RvOX/hDhANmGGaGQs2JrLsf1WgFits8LVETDMfEhUvYDzdV9wvbg+JmYmJJNVFEsaoAKGkjOYuz2iAAVtOqm/jIZVZyjuc7zJdJPE+OykadEE4/JPuI5OMcXRfU8lOBijEAQnGuQbD7FiJl9USxm2pRN4XcIIHD+5Rhi//G4DptNgHg+WwEHqCBLi6wMC1RQJq+YQEVE5aKSCQUqSkqKDFBBMNqPsdFRYSeQocn7EgoWCVAxNjYuwKIAFQY4V3k0VmkGTdEA5QOVrdJvgAquhWyDTZAIY2JyTMaPABVTU+jt65NxJBraMzOSrOfvXFcsWKBrJpmBSWc9Yz+oR4UWX7B/JFlizDu9SRkLrHrjeDtn8G9W/pD+GBxfZILwfnE+spmUwkBFQOTHWLiivhLsR9VdViPVfDNttpPXJWba9Kgg0BKKyLPCKY6+IWRU8Fj8rE0gsQ/5c3klTcijiOF3TfppsT1TXu1Y/mazkAi3mdvzP6i7qIKStQs/6P7FeoA5JbfWo2Kx9PgdMueLncduIO7Ujo/7XsE9p9mrzd9ymkSTPbSVfiopjRlpJcs8hACYnOM4Vm909uK5n70sLFseual1KR77/GFhk713/AOcfPsDZ1/FH/Yc3IX79jIJnsALzxxDX/dNef9L3/ycfJcMqItnr+DimTZhaZhaB7tEOVe+vLURj/6hZVQoUHGHu+B8z/oTP2XNtD+6CAtUKBbhHkX3jvq7dE8uh0fuAlRQ2oeeCY3LGkQa6ZVnX8X1K9cX3LGvfOfL4pVx/VoXnvn+z919dg5Y1roUn/3yYyIpdPKN9/Dua8oW0daZKgyJi3T80dfh0GcOSvK1/0Yfzrx/FpfPXDJzqN7o+bfbAhXnTp3Dy4ZpIZXouSzWbF6LI198TBKxJ15+GyffOInm1c34g69+TtbUd189gROvHPe0Cdj/6EHsOfyAsMyf/adfChuDCfzVG9agt6sHP/jrv3fvgflp5fpVcryRW8O42d2/KFChK6dlyZoiSnNRTFYe9AIVP/gZOtsVqJjvUUGgwvbDN//s22hdTY+KTvzASD9x/v/Ct76MLfdtlfF86aOLeO/Nd9DX1WsKKd2xYUFknufz33gCO/cpUPFX/8t/dpgFdjx9+z9+FyvWrcLM1DQ+OHEKp0+cwq3+QbdKXuJc9VKw6xHvg00C2/2d3SurnA7Bdi3asbklFgEKQ0/WM+1kd89uKigN+1lHk6nSl7WHSXY1oeZ6biV7lDXBPYyeRoyXjf8B/5WCC7NXVOkhK92jvgcEVqQ8KK3Xw9/DwRCmpqdlz6YMaJoe+6TP7WDltVopw7k5FgD5pcDSeRbdJ1MYFfbpsH0lDAIjvyuxgEmGB/yMPUJIJDX2YuELCzMYb9q4UvJS5oK1T5QJaoEh26fSz+JGrhJc7DPeDxZhkDFsC3ztfdC26zjmsRgv2GIYjc2UWSBgRpZKHCmJucWzhNt8I5XFfmGh549+4DIqrPQT+9j6OPA4jI8YL7KgToqSTPEfYz8189Y9EHM1lJO0zAOOL37e+mdY+ScHBLNAgOM/oQ8kcxgCdhkPMFvoaQEjBUDc2ShtYi8FGBRs4Bhx9u7iFUlDdgXE2Cc8tgW4+FkFZJRFIYCWsI6VSWKLUCSm5F73U+mnBWvRp3/4He+Bv/juA+4SryUM865IK8AXVtOYz9nvOAHjvO8vCBa9f7DHMJJF8itPxknZPsiqx+s2oBDgYYMvnSDc5ha4FjPd6/VYAyv9nHzPJuYF7PAm/L105QLXIAdw/07Gg6aFFrbBncTy31NWmgkcbbyQ56nEAM6CRfPM4swGWRfBRRgVskGYH+ryfPMNz917a2+r2xyTDKPEkjAqFBgQwEAYFUzAJCUYp/62ABbTZFLMCFBhGRVW+slW+dnFzSZpeBlS5T+ndEyaaQujorxMkjQ8Hl/WiKm8okISKHIbDFDBRXIukcSNrg4Po6ICOSL4/gDqlixF7ZJGReBNFbx3gWZAMjtHqQ9F2b2MClmcMinxlyBQEQ5HUVlZgUCAlYuGUeEBKngMLkKSLBapHC6iwNTMtAAV1JWvqqhDvLwc4+NDEgyVxmICVOTSaSREpigluqID/b1oO3/eASqKiuNoXbkapVVlYuDpBSp4PiaimKwlUMHFUemlWuXgZVQQqLDsBgtUTI1PCFDBl2VUUHqqurpakgsWqOCIGbo1hA9OnUJNdQ2amptQWVuDmDFVFcktk5xRiSOVobBAha1IlUApnRZfjMFbg7Lw2jbq02GrIFwzT3u97J+GxjrU1taYhFJQKo9tYoPJWFaaWKBC+gXA8NAtIJfEipWt6O8bwJUr7ZicnEEywSTeHNpZIV5fj4cefkgCg4YljQJIMAhVTfakmHATTGPAwcpTgjVMlOreWNtM6ScCFX/8x3+M1WtWwRcwcmBSVUtDcgP60chMKlCVUZFKZXHs2DFp94EDe1FTUylJRnsPNdBm5T0hAwZqfgeoqKupwf59exAMapKISW45l9ghcxxqsCNm2rMJHD50yAkubYJbnu1MFhfOnxfZsQMHDqismDlvirqgZFR09+AyGRUEKqoUXBAllIBfzLRPnXoPTcuX/UZABdcA9kNHR7fIiOQzKi5h06aNiMWUUXHl6jXU1tViaeMSTdpJpY6+7gRU3Hkp13nSvmwgrkk+pQXbxB8/463g8h53QeWrGRuMp8k8IlBBgFWquPwE13gsNb1V8zpdK5NzUwJG6EaH1UUM8jn/Ecigtq81ynU3DgpU5JDxZRHI+DE+NIK3X3sZVWVBbN3aKlXLx9+9BF8I2P3ADpmLQuE4otFKbnfgy/mRSE7j2rUrKCuPC8uIHhIc42+/9SJqaspQXVWC/r5uATLpHTEyPCkgVVl5Mcqr4igvrxOj7omx25iaHkRlRRX8wXL4giU4/f5JjN28jnBgDqFYFBu3bRUmVnfvCGaSQMe1DrQ01WB44CoefeggPvjoOm4PdeG+3dsxngjjfNstqcIOYha7du1VwqEBi2TDairoLl6+jJv93UjNjiMxPYSiogDWrl0t0oBDt27jRncvKigdtW4TwuES9PQNob5hKeYyEKAik5rER++/in07NmDN2o240jOFiVQRouEwqgyAOx+o4Bggi46ANtvFZLsFKkpKYguACgvEioZ5lJs9ZVzQq4LLuAIVOWF3MdJgItmCFfy3ceky+E3ynOM/ZLR9I8Ew5tIpzEENDBWoYOJfK+U51xKoIGuOPzM5zr8TFOCYpiG2ABVFBqiIRUVK0AUqciKrZIEKFhTYtYNABYGkyip67GjMwPWDyQD6LPH56bh2TeSw4qVxYeNx08YENpMT9O5QoEIBDs63fE+KAQhUlJFRyCpCTYSz4MMLVHCzXmKBCjJTcgQqoqBBtBeoKC2NIRTR551AxfjYGAIBn7BI2P5QqAg3+2/i9ujoAqCCjyrPz41mOBwUwEITLkBPT79s7i1Q4QLTaqZNoILXTKYfvZvY92JInkhgctJ6VBSZqk+dVXguxg/8l5/j5pYG4fmMCk3E2BjLzkeW1eHUG80LDSV54/fJuLNABRMgCjpofJ4HghrNbPY55SJTGUo5qgE2YyK+mKi4K1ARJfNIzbQFJBsbFZYOgcrxergAACAASURBVAo7liyjgpWGZeVFKCbw6W+UREQhM23bV/baC4EzC+f/j5MW9nyrYNLcfd85mvnc3dnr81tkqjrvvFDlvavn+PjXcZdL0GObw8kaKHuHRRq0yGm18Gfhq7DY8N3aX+gkTnWIbpcWacfdPCroP3Hgod0CWFw6dxUv//pNafT6Tavx4GN7JWl+pxeZBJRy6r7eJx9b0tKIQ488gNr6aufZScwk0XujH2dPX0RPl37Ovpa3LMFjRvrpfUo/GW8KB2xccHLXkJlvPfXffN0wOC7i5WdfW9APNADffWgXWlZTPlbBce9rAaPiwd2478BOM7dqLE5ZuOd/+pIk4eVOSV9rhz/1H54UCak7vbgOvPfW+zjxqjWJNiBFgS8dfvwwNu3cpMUnZn84OjKKyx9dxEfvfuiYG6u0TRZMnpNRce7UWfFTsC/23/IVTXj8q5+T/QnNnslg2LBjEx75wqPO8Rdr9+TEBJ57+pfounYd/+bffhPNq1rR1d6JH/3fLvvEzoveY9g0Bj0fHvvyH8hbR595/v9j772/5brOK8Fd8VW9nHNCjkQGCBJEYpJEyhJp0RItS1SybPesnu6emX9g5if7l169xu5Za1ZP25ZsSZREijmBYAAJAiRA5JyBh5dzrPfqVZy1v++cW7fqVYGER93T8kJJ4Huvqm4699xzvvPtb++Ns0dPi5QmF4Sc1x58bCdWb1KDcysJY/dDFt+r//wibly5Lu1PoOKb3/+WFBR8sv9jHKBHBdeXXg++/z//GJ3Go+Kf/5bMCb0vZD587U++Lp/Ze07wqa+rR7wkLp9R1gOLBCRJDYip9uYdFqj4jy7JH/180fIl+Nq3/0jkn7QfpMWP5Nbl6zhy4LDjA+LkE4T5a0AE6XY6V9uxQQyyOY8bsIrzms5fpmjNVMLrwXQtKFI64sOn32UswLUO9yFCqMmEHIPrcMa6lNBxpIAsg4frIrM9mQMEzAUoyYrp9bxt26mhcabgjNdlGQPyrJLIavwYpHiLyWVXAZGyIFgNr+xHKRSjb4P1zTCgjHo2UpIpqV4T8h2yVZm4t0wJA/Q58zPZ7pbtqZkxe09t0bGYdAtopGsZy8DkWtYm4dXgmiCMJtXZRlZVwK577PrVxtya61BvB/GFMM+sZUPosQzYIwuY7ImEq5Xnf67POl/f/UlMClDV34NG0yofyquyMp+MaRlTqhm4rnml6EvkmixByRiP0z+D/ovxmOZmzPVRJps5LesfqeyTzNxrDch5bPYtno8FXywQZI3Oed4256L5H21/m6O0fc1ZpwgjRJ8p2b/xXCOLREy4KTVmJK/Y3uzfjIktqCjskntAhXvYvff7v4YWUKDC/dIHL/MqFIXmbOP8mef7WW8Z4CP3+4Lu2qjSJtRdySH5vNAxlX6oL/tLoWswg07ehL3dg2sfttxFy00yx3B+zXc8WxdSABTIOk/XObsjavemhW6B+32HyueewbOTaxIMZV135twzC7fcyUIv2Q3pyNwrAIUFKlTP0DHTjlmgYlbQbgIVEco+GaCic+V6/V28GawGoAYXBCrcFd2i702D3MlJASoor8OJyDIqOFDz2JR+coAKTuyJpEgusNr/5vUrmJ0eR0VZpWFU+JD2+tHQ2mKACq9saydcO2nwuNH5GZOEZNKYjwaTDxnpJwIVqSQrAotRU8Mq0jSSKbITFLCxE5hUIQToqcBJUKcpBgZMykQiUamcr66qQ2lZOaanR4TdUMZkMHUz4wnxQhCPCjIq+npx8ewZeIVRsQTFJRVYtGQZSmuZWNRzo4ErE55WEoLJTkpHuIEK3ld7LQ4oxCrbZFKqGoVRMT2NiTGV/eC2rNZltW1dXd0CoILMBAtUdHZ2oqbRABX+AErL1KSP+5G+Qp1J8RShD4NWetgAQLxGkkkxZbvV1SWmqUw4s6pAAlerj+qSnlCZqJSYE9bW1jjXpbriTI5oQGeDEp4Hq2T4or66FzGRGSJQcePGLcxMz2FuLi6AG5PvNGfe+8heTE3PoKqqUiqWmQz3EZBMJUWy6rac66QwTVpbWyXppPJN+vR037yF3/z6N/jBD36AZSuWCSPDUm1tYlMYCom4UKK1Wp6U1RT2v7tPkl+7dz+EuroaB6iwQI8yk5LibeFhUJjyCaOisb5egAqfXz1YHDNtF1BB0OP82TMCilH6yRp82QWx3LNkCmfPnhVt9j179jjG1ewrMdFD9aK3u0faavOmTeKnIQEtr8Hnkerro0ePKKOis1MSi7bek2yR1atXo6Ojw+lnsWgMp06eRGdnGxqb6gyFOYlbt3pkPFi2KsOouHDuHNavWycVz/Mi/XQDtXV1qK+tEw36EkrImICYyd3chN2Xmcc1yM0YzLkXKjYZ5E7A2edlATCRezCdjrR/eoDKinKRMmOisby0VJ5FAhFyzmKSrWPvdGQMN7uuIxQKoL2tHV5fAJ50gOlwI//ExZAu6mzlDg9NaTBK/3iSQXgTPnTfuIJPDryGjRva0dbWjOHhFD47dghFpT5svX8LKqsaEAxUIByqRjpJoGIOp04dR3NLkxyXYBoXA11dl3HixBGsW7cMY2OsxuczX43S0irUVFahKORDgjI0ySIkEz7c7rqB6ek+rF+/CfBWIukpwtHPDmN66DYS86OobqhD+5LFuH27B6Pjc6iubZaEcXtzJS6dO4Rnn/ljXLo2hSsXj+KhnVuAYK0AFTQFXbm0HS2tix2Q0EnseDzynJ4/dwYjo31IRCfg8cxhyZJFaGlrxc2uXilOoNdOTXWjABVefxi9faNoamlHnEDF1BRi85M4c/wAdm1ZgyVLV+Li7RnMpUrkmaiuqpLnn/MSn2n2Vc5hPAcuoumtwHtCmSHOHQTsCVRYMMCysThuc1FDuTcxrI7FZexNxHXhJ5XtSIv0E19MJnNfFrBobWt3pJ9Y3ecXneYkQqwUJFCRVuknmeOiUWNmnJF+4hjP8ZqgK7/DhJQAFRH1qCDLYz46J8l4Vr5NTYyjSDyYtEqOfksWQNZr94MJHv4koMAOL1VhZM0RqChWE1oCFSxCsIwKznmqS+0VRgXbzzIqRA4SKmXH+YKMClsMoPOJFpuwup9jKRd4JcX0zmBlIHWcM0CFAPrCqJhBaTlZFspWSJNRMTEhRQWhsCbdfd4QBvr7MTk1KSwDMirEfypH+iko0k8KVvCzntu9Mo5aoMKCNWSEzMxOO4wKypcRqOCcRzCcsQ5ls9RMm4beKpuo8Yp6NHHxyyIQYVTQUL7IFkVoBSRBh9yXtJHxu9AxUcchBSA02cU+w34nVYtkeEgVoc41bmDWzutc1HO8otwWq1/JcrNAhQKHGZlNng/7AD9nf+a9HBuj9JMCFQE/Tc69GB0ZQSweddifbkYFE3lVFcUIF/kR8rX8YQAVElC71yxfZgYyUfiXQhIy+/tvAlToqTivgivEQvjIXV7DnYGW/ECFLocyn+UDK9xAxdHDp3D4o88X3IivP/0oVqxZirGRcfzqH16WcdgCFSJnNz6Z99nijsioOPTBEQz0Dekayixh121ajeUrF6OuoUZAEJt8OnviAj58x1bxA/9SoMJeBIGK2rpqnD25EKioqavGE898BXUNteprNEz50gkZRyprGN82qfTT3/3CaUYr/cTnj9twTOE8cPtGt+M/4VZV+MG/ew61dTUikTdvYm2ngY0GP8ers8fP4tSR02ahWZgFxG5Dc+yN2zeibXGbSCpxvGd0PTo4gvde248e8fdQWSI3UEF5p8wrjbalHcKeYEHWZwaoWLtpLR57WlkWEyPjJkFtAjTX1mRUHHjrffR39xUEKvLFffY5Wb1prQNUvPu7t3D++BlHzvGZn3xHAATOCTQlHxkcloQ0jak7lnaKjwmBCiv9pEDFM7LuOWSAClsMR0aFA1RQ4ikn57Fqwxqs37YRzZ2t4othE8sXT52XY2gRnqZUnvo+gQr1qPjb/51ARaby392u23Zux5rN69DY1oySMmVJsiiNAAjBHTP0ORkFxqgeSdQrCMGcghRpSHJfK/1trM33NTmfYQvbB4vjnIDxJv/D40qSXdaWHgFdGLfwpYCFrjelCNEAJlJcJDLIyuBULwKNt3g+1sdA50Yr78u1UcJICLkMsV2+nlbuUJgXpgLeqj/YeVzXfXpdEtsxt2IKBSxwwPwH50oWlvCEWOBhvQ3JMBUmvmGOCPOEcYLN1RjWiAUMyMy2OR+Vp+J6IQMoyLGNH4MaTmsxqybJ1cybRRdca9r1lO0//JlJnKucks2pOOsw4+vhSBjlmRMIivz65yGne33nB3OOTBTPmXGXBaj4JcbXNua2TF0Wyur6n+CK8QoVU2reY6H5OPdfyVvsQdo2+gxnZjcFGBy0wylG47HZ9ja2kXY1a357f23/ZNwkrAmXX5heoN5bthXjZ0pmsn3Zt+jXxrYQyW7DKBXgyIBqbAdlW2g73wMqFkzj9974Q2+BhUCFPjSZVz7gIfe9L/p+TitZ1oJzJDcwIKWPLvmjnGS7s6usLH3mXeftQj4N/ELulG03z+wzi/Ugb+cu9CzT5G6BCq1EWdjG2dVSX6riK1fhyUbCedvIBlwusMX1vexqJr0m+aa5PEsXFsbKAqCC1ZFMfMQwF6OZdlSTMAacIJNC2BQGqOhYsU4SKpQU4HVa0ypODGoWmdFStFWf/C6ln8rLy9XA08gUWSCDVZqOyREn5bhWaw4PDqG3+xaS8xGUi0dFlXhSwOd3GBUq/cREhho9SaBgzIqUUcFEiVbHuz0qOIlIciCp1Z7V1ZWy61QyLgtrBud2n1IFEVCpAivhwuSxSj9F4fEWoaqSif0SASo4KVWUliLFZFIspkBFSgNWh1GRpkfFYpSUVqJz8TKU1lQiGNLEAJNPwkTw++Q8GGxUVStQIVJQBtnjdy2VUCRKJKmRDVSMjyqjgi8x0x4cEoNjtq+YPYn8FeT9Y5R+qqMpbSdqm+qlYokTKYEKMaGWgIzG60xiUK/dJPJMQMrzYiUM3+f3R4aH0SsyGyo9UkYzVFOBYiXCpILVABX0faDmu61O5T7YDmw7PytPGAQYPXYrS8KKzYAvgda2FvT29IvpaTSaQCyWFE3Y48ePo6GpEXv37hGWEBOHTCItWbYMJeEQUgnK4UQkOUPGAc+LyTjKDwUCCs4w4Kb00wu/fQHf//73RfqJMl1eP+nQ6tNh+5wYl1lfFAEqknjnnXck+bt7905hVJAmypdKkFHqTPU5LVDBpPIbr78FYVTsfFCMirW6RE1VrUcFq0foUcFkf9wAFbY/2HtugYoLFy6gu7sbe/fulXvDvi/SLMbvhB4c1qOCIIEkvAjUeCGGgkePfoaO9nYsWUygggGf0qR5bWvWrEFLS4suSrggiSVw+uQJtLa3oLW1yRiHpQWo4PmvWL1cZJCoz37uzFlsWE+goigLqKA/B6tQigJBAS3Z3ywN9wsBhNwpKw3VtRczOksnz1RWFRUpQGgBCvfm7mPljusqcyApUfnHROS1q1cwMTGGrVvXa2W6h1VdrD7Siip5hpJxfPzJAUQi49i8ZaNUiofDZUinjA+OIyOQK9FIszYCGEGkEx54UglcPn8Uhz55E48/uguVFfUYHBrAp0c/RWllJXbs2ImiUClKS6sR9JUIsHry5AksWtSOlpY2ZeQkkhgZ68OZ08fR2lKDYNArQFFFBZlNRZiaHMOtrmuoqqlDS9NSJOI+3LxxFROT3di0aQvgU6DiyOGDmBi4iXRyAr5QAHNxSsFMob5xEcor61jih0R0FEO95/Cn3/kOegZ9OHXyALZvvw/+4lpMTBfhyqXr2LFto0hWZar3dM7jfaD/xPVrFzA22gOfN4bmpmosX74cly53YS6aQnVNBbp7ulFdVY/VazYgmQqgf5Dm1J2IJ9MYn5pALDqB86c+xq6t96G9Yyku3Z5BFGWO9BOfDZHSM0AFx2KbrCegbRkVwjScnRX5IX7OOY5jk5Wrs9JPTGbRm8Jtps0xks87Kyl5dQQquC8LWLS2t8s8J/OZABVc5CfkWcgHVNi+Kyy5YLFIvHGcE4k3mmhPEShPClDhD7Dys0g8bQJ+Jq2imJ6YQBEXhFK5qKCBG6jgAoqsAEo/kdlnixF4fm5GxY3r10U6ilViOl+ojBmfG8o2MYlNzx62kQUqhCFmpJ8y7DkWH8hSW4AKJtAtUCHjG4EKSj+VKqOCYzDbWKSfysIIBE2MlvbJ3ENGRVFICw2QDmB4aGgBUCFVe4bZahkVHLMzQEWfVCJajwoB6U0fodcRxyfO/wQqKP0kfxerzCXnKLYHmSyWEahjCedzZZ1K0YRIP+mcJ1IXyWygwj3+KLCqAZ5KxylQoYkG1aTmmMc+xXPgnKcSioxVM8kim4TQOYzVjX4MDw9L+3JM1nutElSFgAp+h74XGaAiLAt0XuvwyDDmDaPCfX8F4AiwwIPykn6EPE3//wIVd1oMmsEou/6oUCa/0I4Kf7/QfPb7BCrsGsGRDjKn868ZqHj8yT24b+NKTE9FsO+1D3H7Vi8WL+vA41/fLUVBn358DJ9/SmNnW8dmGiXPrcpdnhE8aWptwEN770dbR7MAjvtfP4CrF1XWp21xC77mYlQcOqCG3faVC74oXzLzuhNQ8fATu0GfCibdabR986rxl8j1qCBQIZMnYIEKjjHHDh2XcWLzg5tkbObfh947nHX8Z3/6bbS0NePapWt45Rev3unpyP6sAOMmH761bdc2bNu9TdaE9HR47ZevOnryP/pfM4wKN1DB/rtq42o8/tRXZX2k0k+fYumqpcI0IFPm0Lsf4+hHn2nC3Mg4OyfpauRnfvQdLDPST//8nzPSTws8Ks1SmvPMqo1r8JVvPSm72//S2zh//KyM0/c/vAO7vrpX5s8Db7yH458cdeKWXU88jB2P7pT1yKu/+B1uXr4ucagAFd/LBioksZ1K4Qf/4c/Vi+LKDfzi7/5R5p58cSnvZ2VNFb7yrSewav0aOf4Hr72LT9772JGweer738ImC1T8H/9RpYIcBo3pIIbxrsleoG1JJx5/+mvoXLFYis5e/tkLOH/irLOdsAqgOvw2OyGV7NAiBgHNbbaEa3TJPSiLwOmUcmhVROBLwAojLax/k3XMeVnnWgW2gKBJFvPeco0gXnssKDE+ECyi4/FsLELJJh6DQAlfnMdslb2OvXpSCv4r0C/SuAJMqEeXJLplfaMAiXoOKDhgJRGtn5wtLBD2gSRcPKJWwWIzy+TgPliMOBudM4AE52wWKyl4InO1aSuROBIJXPWoc4AK0/B63QyxNdbSWIZtpmbT/JDHZhJd5nsTM1jjcZ43YzJZuxlJURtTsl3cxVIKzKrxuKx1peAi/yzyq59lWGvf/v6cFDdK8afxvVU/P3qlpHRdbxgcWgDhk7YTUMoYhfMXldbVol22C89DVCYIJEk7aQGnMk+sjrwW68ocKKwI7f/ST6ToxsQ32mkd1oTtg3qtjNMo4xR02lnuL9nFwgbieWkejTGp+gnq+fH+67odwiSxvjK2wER9xoy05j1GxZefa+598w+jBf76Jw/IiWYPFHcGHjJkgnxJ+nzARjYyaSlemZS5axtBI10TaiEZo6yQzc3AsNJ7uk+7mMu+G5Ye534395rN9s6UaCej7O+5oY2sIECkn3Ku233OBbRm7T6+HFCRp12zAuSCSwgTNuUDZqTVNJiQDJoe44uBCjIq4pibj2KejArKPon0k4IUVv6J7y1Zs0mSB5Ru4CDMBbmla/KnTVLbiYyTjhuoYPLbVqxaaSgyKmywwkkkYfQYb924iemJUXhSsSyggtJPjW3taDDST5zQeK6iy01tbJM4jifUo0IN4UlF1cS+TCqppCZr4xCgoqamSrTecxkVlj7pMCokYGA1vQIV1CtPI4D62iYUhYsxOTkklSAKVMQQi84jFp2V4INVKjTTFo8KAhXtiwoCFZLwYgWGABVknWQDFTZ5xmvmJChmnAbpLzKyTmKmPTJqghcvJienhFFBaSPuX+S1iPSL9BOBimNSyU4z44bWJgEqGOAQqGBSjYleC1SoLrUGkNLehmIbDIWEMcB+Qb3ukVE9PkEASlERrGClvAZXOkErUMEgUJ9/nhdZHwQMRKZIqJxK/7XMDsvKIaOiOORBQ2M9err7MDQ0gkScQaUXkcgcDh78GLX19djz8B6piGVwFKMEVGMjmpsaUBTwy3my/8zHWCk9K5rulCOrra2XoJiv2zdvCVDx3HPPifSTL+BzKnFtf9O2iVHAx8WoyAYqamurHEaFBWtEp51BFiuUWOVigAplVDwIf4B9l0FdBqiIE4Dz+B2gIjY36zAqhJ7ssA80DD9//rwkevfs3YvysjLRYOWL0k9yfV235Tvbtm5FQz3ZJl4kiFJYoOLIp9Ivli9bKgbx12/eQl9/PwiAbNq4Ue4jmUAMZP1ePwYH+rF122a0tTXpceJp3LrZLbTeVWtXSrBNL5GzZ05jw7p1olMeS0RxxUg/UYKMC6Seri4x62b1Mw2G7XXdzQzNwLa3tw/nzp2ThLGtkue+6E2zfv06uTYrp/Jl9+0GKmTeS6fw4osvoKGhFl99YpcYM4eLyiHFUvQsMUBFMsW+OYUDH+9DKOzBsuVLUV1NBkmlSEDZNemCBBZ1YWNxRGMJeANBScBybPzkw30YHryJ3Ts3CkOrp3sYH350GEx479zzgLAzKoobpX+fPPk5Fi9ejMbGJkxMTEtSMpGaQzjsR2cn/SfCMr6xiHJkZArHThyG1xPHrt0PoyhYi2TcjxvXL2FqphcbN21EylOBlC+Mo58exGjPZUxNdCMSm4OvqBjNzYtRU9eGyGwC85EZnD1xEPWVkGdodKYcnx/ZhzVr2tHQthyRuRJ03ejFfSuWAH5KImXr5fJ5v3rlCrq7LyMRG0dpOIAHHtiC8+ev4sbNQbR3rEJxmR/dvTdQXVmPNfdtxNx8GiOjU2hu7UQsnsTU9CSic+MCVOy5fwOaWzpwpXcW0XQZSktKUFlRoYCYAWP50wIVHP9zgQqeE+Vx+GJCWKSXQip5Q+o5E9XSr2MJAUNpMs9nWFhnBLZKOA5mgAom1Xm81vYOAQK5KA74/Cr9RJahC6jgc2SB4lyggh4MPA+OnexD7PO8Flb+c5867s+JXBm9mGYmJxGi8SIX6Qao4LNgWZN8n6wAsuIsiCGLSUojBYoQKtICBTIqeF7KnlA9YVb7ccwtLSWbUoEKHt8NVLiPqWyU/ECFlX4iUEEJI5qV06OCx47Hko5HhS9gYqu0T2IPsvHIXpKqwaQXI8Mj4p0g8kz+gMhsScLDSj/5fcJqcAMVvd39siClnJltb1mYxuOIzE6JAadb+omAA8GJaHRWvBvYrwhUaFLfxreGUSEMQWWfWqCCX1E95gyjIhuo0MSKxl46Ylmgwlaxclsem/3UMip0v+q95V47CNCeJBiRC1QQzKTUYzajwrIwLKszG6jgdRZJ246MjkgbsC3Zbvb+8ncmY2qqCaD4EML/wECFnRBcgMVd+0eYqDzf3PLfGqjIlWVyJ2ILenXfNQ5TaIM77SjfZ/QH1BWMs57K87Uvw6h4+jtfE2DCzahgP3z2R08JW0HMtH+jskKZdkhLrD0+OuEcf+uOjdjywHoZv99/5yBuXqMZtK60Fi/twOPf2CMypUcOHsdnHx+TzwoxKgpd090AFc/84Cnxj+i6cRsv/vxls0u9y195+jGs2bBKGBU//7tfOmu/Byn9tHOLsIzf+d0+YVJ8/dtPYPnaZYjOzeODNz7E5bOXnWt+/KnHsGbTamE5vvHbN9HfrV4d9kXpKTLeuX7IeuUBKr77V3+G2oZaXDl3BW+/mJFx4nZ/9OzXsXLdKgwPDOPnf/uPXwqoeOQbj2LTA1skPnzrhTdw/eI1kZb7/r/9IWob6nD90lX87h9+a2RwVAKPfZ4G2WPDo07X2vPkI9i2W82036SZ9qVr5ilNC+DxZ//mBwICEHQ4uO+AfEbpJwtUvPvSWyL9xLjuyWe/iQ3bN4lH33/56//LaRJ+xuM88IiaaRcGKg4K00OquVNpPPfvfyJABj0qfvaf/ousNeTYzzwh4/6BNz/A5x9/ZqRx/HLd3/2fnpNrpCn2a798yTmHp76XH6jgF3Z+Za/4d/BevvGrlx3pKE4mK9etxtM//BNh6BN8ef/1/ZnrEnkpk6j2MoFMQNsm95nA12Q55xV5mk2RkClYN/vRJL6drzi8iqGw/dQYs4tsjpGGZiGlSAXx+JL8NRJTRgKa+2BeQdZWaa731OjYFiFpLkDnVgtSyDlKMt+yrnXA0SjCGkmrtJNI4sp6TWXOlJ1BeSaPxGhSNCAJaWWAcN3PxLxsY5LljJv43FhWqgVhdH7X3BPHA2EsmOviNRAUkiS3nK4yIxSMU/mnzJzOI+u12PWSMvL1XkgBJgtgAppcZ7GSlSnTxL3GbFp8l614wu9ZJqWySAqN7x786me6dubrme/NSR/hvVHWP4+heRnLJhDFT7JjhcFFVoyCS1IsIYwK9UuzniQCvMh3MowbK9MlOQOX/LvNN/A+q4IBPfE0xtbCO5M3M0oPzpxsADftPyqPZ5UQCJqwH4jihgWlPJoDkwyA9ccwzHgbqymbROM2d3GcrD/vARXZ88m9v/7wW+BvDFAhV7IA1TRVZXe6THnynGkhhyng/jM3aZ6hVsknmf8YVy/nTddO8gEoFkDQiUJf7vNeeFwuiPJVPGRr5Lm9MexAmjugFmofGsjmAzbyXVNmnFbE1nUfjH55wepf59Jy2iXvuJ97rnlAjFzwRDR2cm/+Qo8KekJwEhWgImqAiqiCFEzk5wIVy9dtEQ1sAhWavGFCQqsNmGThIE35Hk6kTIJwQnIDFUyeSGI9Nu8g4RWVVeohzoGbYEdMjUqHBoYwPzsDJOdBnwQyKuhRAa8fTe3taGxtQZq+DXHK/MzKuVgzVJmM0lqtDKzUnwAAIABJREFUqBUUGaBCaKgGqIjHKFlVIudM6Scu4i2jghWJnJhtIKGJZQ1eFKiIiIlnKu1HY2MLgqEwJsYHJJlYXlLiABWJmLIzwmXFGOrrxeUL58V3or29U4CKRTmMCmuQaoGKdIpARdUCRoVlkDBwYDLCAhUMLNkW05OTGB0eUZ8Hv08kQNzST0qvZYWDRzwqyKhgJXt7RztaOtslucLvsFLUAgbWB8MCBmxnvjShosEHuzC3pVwI/UlYOUKQYWxkTCSGmKCoML4XDlDhYXBrpSuUQkwplpbWVhNEEURSpg37miTRAIyNjqK8LCCSSre7ejA2NgH6pfl8QWmTd/fvR01dHfbs3SOBAwO0mblZ2WdtdRWaGxvk/AXoCmggxaQ9n4mm5hYx2OW53Lx2HS++8KILqLCSYwQQWPlqQRw3UMGqVgtUBIVRwSQ2+6tWUCgbQ4EFNdN2AxVNDQ1ZQAW17i2jwgIVNNcloyI6O+N4VIicilkkMJCKJ5K4fPmymMhuv/9+AYDYhnwGk0YuhNdMeaitm7egsbFRE3duRoUAFW1YsXyZMJ4Gh0dE5/3o0aO47777pI1E3oYJTJEPGcaWLRvR3t4iQ3s0GhczbS5EVq9dIQl5yiucPnUaG9evE735WGJePEYIUjU0NGA2MotzZ85gx4MPqjZ+jqnsl53BlY2SkjGFL9FGNXJoVt6FiYbc6iAZdV3zau5YngtUMAnS39eHy5fPYeeu9ZKYrK1qhgfs/zQn18RtOkWD5QS8/hg++ngf5uansXrVGlSU16K0pEp8c5T2bdgfZhynJF5iPo7JyAyCkqQNCuCZmk/gjdd+jcqSSWxcvw3hcAOuXO3G/g/3Y8Xaxdi0ZR08iRDKSstx9uxpVFaVa/W4x4va2jrUNVSgvIwAhcqgpdMBFBdXY3BwHAcPvovq6hLs3vMokCpDMhHAtavnEZnrx4aNG5DylCHtD+HoZ5/g8ulDmJ0eQG1zA1as3oC29lUYHJrC0NAE5mcj2P/mC1i/ogHP/um3MZtuxNEj+9DRUYVFS9eiqzuCVNyPJW3tSAkg5eEQKc84n/vxsVEx0R7su4ayUj8efHArRoeHsf/dg2hsXo6GpiUoKk6ip/caqiprcd/6TZieSWJ8MoLm5k5EWV0+M4Xo7BgunDqIhx/YiPqmVlzriyKaLkVZKYGKShm3LKOCPzmG8Dm1QAXnOiasZmYi8lmoWCXtLFBBtoL2IzV1LQ7TsDopc0UsSsPAtC7q06ks6SfuS0yM43EBKjjPcVFMHf+gl1TypCRjxFgxRf8lmnynZLxyAxVFgbBIvGlFv0pLESRRRsWkASr84jtDkIXAamRySirFWHzHRZ8FIyxQwX5OoIIeIgRw2TFlcRak9BO9jvQ4169dlX4dLi6WxD3nWFZRMllAoJFABZNiZGGoRwUT/Qq4cEzKZlRoFaabUcH+6zAqknEUG0YFn0sCFZMTEZSVhSFAhcRDOiZZRgXHAYLYBOfEt6G0TKrqbPJc5JMMjd8t/cRFe0/3gNwDghEW0LRABT0qwqGQzJNsMzLXCDhwzoxG5+RaeT8oBaUySWZcEW8KMhrTwqywQIWCGZpM0eIPTTC4Q3w7VuUDKuy4yHYhy4HxhHpmMHHACkZlANrz0CrSHKAiyftIwEE9KjRhobrXdgFuEy3a/9zST2RiFIksmBuosPeX7WmBivLKsDAqSnAnj4rsqs0vLgSy8fuXnSEsUzr/97PWG1ml4XebzS90Pneb5DcDY87uCqeMMpWlTt8wCaZ/DUDF5yL9pACBfd3/0CZs2b5eAMfL56/jrVfedz7b9eh2bNx6n/TZE0fP4uAHR/RZSAM79mzF+i1rxYT7zZc0MbtoaTse/6M9Mp5fPn8N+9/8SMZhjjA79t4vIAYNYt9/6yAunbsq21TVVuCpZ59AZVUFzpw4j/ffUo8MzeNbkZvM+UpC0XX+d2JUPPGtr2DFfcsk8f3+6x/i2uUbci7379qGzQ9ukBhZgIr//EuNI5BGPqCipr4aT/7J11DXUCcJ9jdfeBujQ2Oyr6Wrl+LRP3pYDLO7b3YLuEHfDr6WrlqCXY/vlPFq38vvZoMYeagTT37nSaxct1J8DyjxdO2CAgKUgvqjP/2GeFHcunoTv/vHF5zEqmVUcA3x3iv7hXHB17I1y/DoNx9HWUU5uq7fwm/+6/OSBOeYsPfrj2DTji2SeDz+yefq+aCDOnZ9dQ82PrgFt67cwCu/+J20S0tHK77xZ0+joroSXddu4Y3nX8X05JRs85U/fkKAh+jcHN749au4cVHP2S39tO93BCpOST96+BuP4/69D8p66pN3DiijA2msv38jdn51r/gTUkbrNYdR4RFpp29+jx4VlH5SoMJ6EDz3737sABX//H/+vSTCq+tr8exffg81DbXounoTL/3st6DPB2OErbu24+FvPi7j6sfvfIiP7LUDePxbT+KBR3ZgemIKv/1/fonb17ucnrZ87Ur88Q+/jeKyEpw7dhqv/NOLAlrw9djTX8NDX9mNRCyOV3/xEk5/dtLZTpLujBeYcDUeDlKNT5kmzhOsiKdhs5Fkkl7vgFgqVaidUxPHsm408a6sz817nANZICDzUIJMSnpPaHGeFDcyjhfZRo2FgkUhkTjlPmxinPGHxCustDeyVGr0rX5N1v9D/DBcZt66RtO5za6ntD/pfMR/9vuyfpN5WhkN6gXBvIpW29ttuPbzSUWBR8AKsonsMyprOybChU2qIIdsx8icoIVRI7CJdcEpXECFyDqJoTiZFbwHfimaFFaIAXoksW+KH8QM3ezD8c8wZs/yfVeOiteauScqUyQeIoaF4hq6dJ8AnncxKr7znH7Xsj+F3WLYErYdmXuxxRf2XlmPCmEUyb2m/LZ+T+W/FHASE27jJ2JrjNV03HVmzj1TmTJTzuL0H3veGhvpp5ZxKscjyEOzbJ96Q9rPtF8rasQ2531X/ycjJyZ5Vr0vFoDh35J/IfvI5E+EbXsPqMjtSvf+/kNvgb/+8QOu/L7NZrivKkdfaEHe3wIVNkTKkwDPk+y2gxt/OtU6Fqxwl3fJqeQk2d0JdQcQMCyMBWDFQqCCCy2CFe6XGubYY5nfshJMeaSfZOGXq7/kjE8GrHAfJV/78vt2MFSwRdpDM1w6YOdQNp095gWWlAq54CX+H4WAFfPtLwVUmOSXMdMWJF6ACtW85gTPRS1/UvqJyZMZAhbWp2JuDss3rJdECGnHNKEWA6ykGgMlUkxysCrVmI7ORYWSOSHsC2pml8vnXMxTyoHIOQfziuoKePxMTKVFBmd+bg4jI6OITM+IGTX/rigvR1k59bE1QdzY0oam5iak/F7Miw/ErHhYMGliE01psBKQE5xqUvp8TEqwqs8rZtpyHrG0bFNXRwNh9pOUAC487wz6r4ZOSptkFYWi5dRQnInEAF8RmtsWSSAxOd6PRDyGimL1qEgz2TUzIwFDcXkZhoeHcOnieZls21vbUVJchqXLlqO8vk7uMQEAtrvoNBZRS5xao0mUSyKHFZgqRaLX45MgiBOrgESGwkhpEe5ncmIcY+NjxmzKIx4MTPzU1NRIYsUv0i9MLPtEpumzQ4dRV1ePxUsWo7q1XirveRwmnphosiAFE+bcP+8dF2x2UmdbM4i0SWAyFXj8cCgs/csHryTs6AfBtq+rrpFFFQNbBho+obtqcMsVHZ9zsi/a2tpQXKqaqbxenhP7Ke/z1NQESoq9IhlFHXFWjRMcY4DJRcM77+xHRWU1Htq1EwTE+MyTIcS2jqfiskioqCgXFgTZHrxn1NOnFBQ9VWrr6xAIhnD7Vhd+9c/P469++hdYunQxvCGlAWu1jLJKRKMyloDHqxI+DCi5gN331ttyP3fv3iXeGNZMm2AAf1eASaWf+AwU+cN49dU3hPHx4PZtInvFoSqRSmvi1BdQSyBTqXPx/AVJBO/evVvui03E82ffwAAS6YQwWghGbduyFQ119dInyAiKUeM0lUJPdzfOnzsnn9fX1WtFO6uCvBBWkDXTXmQ8KjjqcGHy/gcfYNWqVXKPNECmrm1KJLcWLW5HU1O9AhVzcdzq6pHKn6Ur6EHgRTQyj9Onz2Dzxg0Ih0kLnsfVKzeE8UPDd17riRMnsGnTJjQ3NxsRdk3yiREan1ZZ3Wj9UJ6R0wma8yVxJOElZn2kF+s47gYjCAJ4Od/kCRQkgW5o8jwX+4+GzEc+/RSRiW7seGidSM6UFDcima4Al0UJ7yw8CXpSsMdRYmgWR44cwvTMBFauWoG66joUB9nXg8LU4tqH/SLtMaaAZqzlWMPnVsa3BDA+Noz9b/8WK1e0YunSVmFWfHbsPN794CM0djRhzfJ2lJeUIZXwIuwvliRBfTN9dYoRm4uB8jVdN2/g8tVr2Lz1AVTXt2FkdAaHDu5HMJDCY499DaFADRLzfly6chaJ9DjWrl0mwMXFa7dw8vhRRKf60VhXjg1b70dr5xrMRYO4dOUa5qIJtDa04e1XX4Av0Y+//KvnEElV4czpoygpSmL16hXo6hlHSVkTampb4GeCFj4kPMo8YBvdunkeV6+cRBBxrFy7DiXldfjVP72AinAFOhZ1orKxSqrQ+nt6UFldio2b7sfI6DxmImk0NbciSubA9DTmp0Zw+fxn2PnQBlTWN+Nm7zziaY5vYZljmEzn+Kb+SSkjtacVgkVFlHliX6aHUQzTM9MIhH0id8eEMJ89NZZWunpxcUAT9kmyGuZkOy7GAkE1UA8XlzqMCoIJTKDzWaRHjh3nbBU6xzqOlVJ5nwLm4zo/ScUZzbRJSw+R3RCWZ53nwn9kY3Bu5Dw/Mz0icxcBWY6T/FyAipkIKH9mq+Tph8TxgWO0JMJpvErWRTHHygplMMRVhk+kn3gd6TSuXbki7UMJQ3ot8Hn2GkCQTARrps1tCIil0mqmzXGDspDuinu7CCQApFV/9KQoUap/VBloxSVFaqbNa5yNIjIdleS6P6gLTMZiZKnwfO22BI0GBvrl2mj6bQ0PdYHM8Uur9vTalAXABXF/35A5B2VUyPhDgCQex/g0vRmKhEnCOW+gf0CBi3BYPDvoh8F7x7jIDVRwDJmNzsv4wvvKsJbfCQXVhDKR4rygoJACBQqAaRWn6ksryC1hkSRH+L6+p8ydoaFhGUfZvuIB4tPFs8pzmBjVsO84qXBc4TaUMODcKIB1Su+RjYHsdrayUuU/PVI0oB4VKhnFn6Njo5idnRGQTeImH+MWnccJ7DKRy6KBEjTeQfrpXwJU2LTDl1vlFTaD1u0zkknumeT3BVTkO0cDRuRDEgocNm8Bl12j2UnMta0UV90tRlKoOfNp+zizb8GN8s6sd8Oo4Pw1OTEtsR5f7P+lZerzwn46PDiKt15+H6Mj486xOP4++fSj6FzSpkxQjh0zs9LfOX5wTD322WkcPpDxvdixdys2b18vzwB9dmamZ1RGtFTZZLeud+Pl562XgjbqU8+S0dGpz1s8ge6uPrzy/Bs5K1XTv+4CqFi0rENABLIa3M+yVEibSmWe31sv7kNvV5/ERw88fP8CRgWPvH7rOjz02IPyrF46cwlv/W6fc37bCcLs2KwMvFgM05PTkogrryiTeL3rWhde+/UbGVaFqTLPvamMNb7+nSdR11gv5zs1OSXtweQ9901mxMfvHMC5Y2cXABW2InzK+CxVVGnhEAGMfS+9IzJKVpYnUBTEN777FBavXCL3ZHZmVtaQJZSTLS2WMe/ogU/xsWFHsF02PrgZe554xMytlEGckrUGv8+2PPLRp/jorQ/Mkt4jQEW29BM9KpICHjz13J+goblBYlKp9gelcANyrUzcMzH9zguv4+znpyXuzAdUsO34qH7v36pHBYEVSj/ZuHTzQ9vwyDcflwQ3Y5DJ8QkZa+n5wXlqoLsPL/z98xgdGHZuw33bNgjjI1QclueERQpvv/CGgCx8PfrUV/Dg47tUdnh2DlPjnOvDKKssl3a8cu4Sfv6f/mt2hE0gXUy1lQFiE8X8SWBDqsZNsZRICgkokCn8sWwGzjlsL4ItZLzzxer0KCWOzbgr840ZX+ya2K6BeU8tAM5t2HoaJ1GSmYUejLUyxs9cG7IPiuyxJPEzoLYk4yVfk2FpqD8WC8s0sWwBRdlK5IU0oS3Xb4BIqyzBv6W4kdJURrZYPjMMBn4moIrxsbMxCBmMLKCwL/X/ULajHMM11sqvJj3EdagtJmCfY4zHGETkz6SYQ+WxpT0NA0SySj6NlfT/jO3Us8Eey2JKBFmsBLaNAZXdsnAS4Xk9//OM9NOf/pCxHk20tT0EfDGAgG1XglC898KaMTLeolZg5Jdt/2EbSjGH1yOFIPq+ynYJAEUzd/Gv0DWdjVdkrBTzdJVusMUacnzDqjEX7fRVXrPEgOZm8Byt34m0lhNDWcYLARhln3JcYJzIeynyVBwPfAHJF/DFsY9xqMb6upa7B1Tkzh73/v6DbwECFfqQ2kvJLDz0HasSaL6UD6jQ7IzZwcKUTKHg1w1AuIP8QgwCBQVc+zfm22Ia6pFsjDll/am4BxHi3HPiqoyTSQZkyFy/fS97G4vk51ZiZcb7zPcF3eXAywheztHdTXJMwc2BRX+xAAWu0AJIqqdloMtBffOALjp4Oq2S5165T9K2o5lEHWMhHbBlojVARZITuGVUkOUQVxNpy6RwGBUuj4rlG9ehp6dHqi78fi4+faIPTeChvLJUKw7NYpkBERP+42Pj8AfIdiiThLeVC+ICmudUXlUmbrQCnCSSmItEhLXBRFw8Oo+p8XFJkBCoIKIuQEVzK5pampHwQsAUXlNVVRUCAVawMnFMmY2YMaXVBTwnegtUqEeFG6ioEeknamoTHGBQyWS4VhRqhb8FKnjL/DTTjsxmgIr2RfDCh4nJfjHQLisOC0iRisUxOz0l7VVaWYHh4cEMUNHWIUDFkiXLBKgQWY6iIqniEdmJoHpIsKKREjVikD0TcfqkVI1IlYiyWSTpQ5NTI0FigQrui6+JiUmp7qR2vgIVhsbp9Qnz4tNDhwSoWLR4Eeram0TyifeHQEV5OYEKJozYrgz01EgwE+xpAMXKXHl8PGyfCEZHR6SyhRXADBDYN9jvmai6ef26JPKqKiolWGJFqph9svLAmsdTyzMUQk1tjWjnszJUFpdzc3KfWc1aWuyT6uD+3kEJRBgQqf5mAm+9+Q7Kyquwa89u1NTUSpKf1bQcQWJJVllPSJuuXrEMNfQUICAQi0v/Y5sWl5Wipq4e3V1d+M0vf4u//MmfY/nyZfCGM9WlFsCRYJC65UZbU2TMCFS8/Y4EYDSybmhscDwqGLQxEOL2vN6UJyXyXLPTURw+fASLOjqw86Ht8PtVb5VmwExoVVRUwReklIlfthegYm4Oe3bvkuDHSlHJPaCkVTKOmzdvoK+3Dw89uEPkvXjvGCTPxeISMHbduoUL587j/m3bQNklGT2kEsgAFUc/E0bFksWLnIUh79P+994ToILSSYWACq3WsR4VMaxcs1yAirnIPE6dPI2NG9ehOMwqqXncuN4lQBr/8R6fPHkS69evF4YFr82O4bljeR7I2Rm4C9XXZoAKjfRFIsC1CPDKNFAYqLBUbqFnmzlLqvJDRXjvzVcQKo5h69Y18PnLUBRqQMpThDhi8KR8OuVBTbNjsVmcOXNSvC06WpvQ0tSEYKAUHm9IQBSSHwSsEH15PUc5d5k6daHIPnvj8gWcOv0xNm1YjuamdviDZXj/o08wG49g8ZJ6VFaUobqsEjVVtQgWFYMSetMzszh29BiWLGbSJonPP/8clbX1WLdpG2YiCRw5fADJxCy+/uRTCHgrFJi4eBpp7xSammtw9sxVXOvqxfjYCEKeKNavWYF1m+9Hdf0ijI5HceX6Tfh8IbQ3deDV3/4CXgEq/gxzqMXtW5cxMtiFzZvWYT7hhT9UB3+wCoF0Qozc+Y9zwmxkDCdPfIyJ8T5hXLQtWor/++9/BW8qhEXNHWhurUdxTZkkB/p7u1FTV4F1ZP6NMgFFLfE2BSqmphGdHMbVC59h5+5NKK2sw+2BBBLpEpSVFYEJeoIRTGZboEIXGDr+W+knC1RQPihYTOkgSgxNGXAgLOAl709piV/GSa7Rp6eVUZFMM8GvABSBCr6sjwDZbnwRlLPzjQUs+EzLApyV96m0jAfWFFX0jGnSXRSU+ZesHgLG4SL1RGDynHNIZGoMPso0mIWTjhVxzEYiMmewR3L80nlUgQr2NY6VnDt0HjCsBmOmzUIFMhIFqLh6VX5yDlOvj5gCFSBQUCqJfCb5uI0FKiwTz+7XAvA2VmHbcEHJ8+K1cRyNzSsjygIV/C6ZjRaoINuRbBS+z/nODVRwPTrY34/p2YgA026gwno3sM1ssl3ug8+Hvr5hSbZQIozzmCZP1IhRgIpwSMAZtnVPd4/6LIWLRYN6emZK7h2lwOx8rVKXHsyZhAzHdVKICFRQ4osDimU+WFaFLsQzWtr821Z66mcK0Nj3eKzh4REZRxl3KVChgIwdq+14J/c5pT5eIgeXYHuHDSCSYUvaY7Cfch/SVkEyxshuHJN24LXaNuT8PztHIMwAFSxI8JNRoX5i1TWVkrwIpxsUqKBklJynAlDK3igEVNjK3HxLuUKj/u9p2edKcP2e9rhwN4JA/R7AEFNVv+AAd9r9nVD/u7lgG8ct2KbAATjP5ZEPyv22lX4qKy9ZsGf2f44zN6/fBr0h6FHhftk+v2P3Vqy6bzm4D2W3JsWU+uTRszh38lL2Nkjjvo2rhIlRxT7LivEU56Y5XD53DZ8e+NwU7Sg1g3dt0bJ27Hlsh3yfr5uUmnr+dV3f5tzW3GUuGRU1tcZM+9UMG8SeVOfSDux4eDvqGzWW4/zQe7sffd392Lpjk8ToB97+COdPXpRNyKjY+tBmkX7aZ6Sf7LJy91d3YuP2DZLQPfrx5/jsgDJMmBegNNSWh7aIcbcURcl8PIvLZy7j8IefZUs/CVCRWxSouyotL8POx3di0YpFMkZoQjQukk+H3z+EW1duamLaSK/8+H/7qTAtLp6+IJK5TW3NKpmYSmGwbxAH932EW1dvaPLDePRIXJSGsADWbF4riXbxkCObe3gUxw9+jtNHM6wAvcS0eEFwm4bmRqfwa2RoWEykTx85qWt7Y8K8dss6PP7HT8g1kVFx7vPTTv6FDI2dX9uLtsXtzn4GegcEENj1tb0yPx9+7xN89DaZHsgCKg6/d1AAEU2eekAzbSv99Iu//Yes/MKSVctETqqhpVGLFAABe66eu4z3X9knQIPNW0ihQSqNbz73LazbtlG+z+++8cuX5doIbvE+bHnofjzw6EOoa6xTTwZKRk5NC6jCfcr8ZF+m72phlVa6s++IpI8BDPM93Sy0YyW6MAcMaGGNsfm326NCx331irD5KV6LgAku5n7mnPSk4kwOc86mpJCcmxxJ/ql0MBkXLP7T4hP1gtICK7tfKQATz0v1UOA6kvOyfE88MdSsWs9Z2QuWXcDYxoJrdn/iZ2Gq7QUsYOGZyGxqzCa5lIDfAT8Zh9h5j/OwBWLI5M1XsGrVPIRxzvtggEWVrVIPD32eTWsZ83Kud9j+vB5J7pt8lj1vnpMyLSktpTuQAhBpK94L27a6HlHGQCbP9Ot/yphpP/sDNUFn29uCFMmrENgy8k6MEygxrQU4CWe9p4V3+qwS8JMYkCCTOR/r+SBFGobFw9Nlfkr6UNKwcFhQKP4fLIrTQg1hu5iXAlLZMZQUfJhiFVsAYiWjRLmA12AKV8QjRDxBMrGRSGt7tKjE3kdlwSpDVW9NZsy8B1Rkhpl7v/0raQFhVCy4FsWh9WXTJ/bPDJBhEWAtIzWff8mq/MyY5wJCnOPlBtZ5kujOOTPBb4AKcyUumMJ8a4HrtF6fM0i6gQ23lFWmYSTwdb5v53A3uJDbTjnXYJEQ523XNZkFa6YRc27IAuaEmTMMXcwmy5ytnPXVAlQpd8eZe5x7DAMC6QCYUdPVQNAGgxnDKGFUGDkm61EhBtpW+skFVCy+b7UwKlQ/USvyWUXOpHplNc2yw4JOM0FLFgEnYTIqfP4ilJWVOx4SHPS5gGa7lVeVZwEVk+PjksioraoWj4XJsTEBKsqZ0BY9SC+ahFHRjHkkMTk1JcmSysoqrbiMMVnNBPC8CSq0YpqgigNUpFQuKcOoMEBFOumwKZiotmh/LlDBCZZARWQ2BniL0Ny+SCrcpyYHkGZCIxRGMjaPNNke01MS0CujwgAVqQQ62jqlAnfx4qWoaCBQ4ZP2I1AhFYdidh2V9mQVE5MnTNxYqQ9OzPmACm7HwIpeC/SI0CQBjUnHZHsm5ITJwPhb9BUDotv96cGDqKmtE6CiobMNpWWaSCOAwESSTcjz3sn2pC4amSGZbgkqGOkTHo9ABasshX1CuSVWc5Aa66VJrF9MXq9evYqBvn60titDRqtHFKggo4JglTwjYsZehoaGRscklkBSZHYGZcXKOBgZGlMJJiZQfAH5+ebrb6O0vBI7d+8SECZYFMb0zIxIhrGvT0xPSCXw6lUrsGLpMgQZRNIQjknPwQEx4K5raMRQ/yBe/M2L+OmPfiyJeV9YkykMdKWvW0aFABWGmspEViyOd995Ryp7LFDhZlQQaNAALy0VtGQSjQ1P4MSJ0+IHsXPHAwgEvJicnsTlK1ckqFuydBmKBbBR6igBhtjcnDA2LKPCAQ1YDYs0Lly4iO7bt/Hwnr2ora7RCptEHNF4QhYDTDJevHABD25/ADXVNXLfk6zy8KSFUUEz7fa2Vixdstihp/N+WzPtjo4OJ+Bnovf4sQyjQhOgady8eVsSeyL9JEBFDKdOnsLGDfSoUKDi2rVbwqZwAxUbN25EU1OTVjHnmLfpsO5WI104uX8RUKG7sFTuzOzG35hozfeSfVrDQHN8LhKYyKSkTCoWw1tvPI/OJTVYunQpioqq4Q9WIAkmle2cy4C59gKvAAAgAElEQVSVtHLKzc3j2tXLGBi4hcb6arS1LUIJZaDobWHYdEnS5AnQmwojnbW00ICLnvmZGZw4/hGmJ4ewYtlypFNcxKZQUh5EWXUZSsuK4PdSWo/AsgceHxlTJbhx7QrqG6qQSs3izNlTGB0fx8Yt2xAIleH08eOYmhjC008/g6C/AvF5H06d/hyT072YmZ3AwNA4AqEKzE7PIDI+iPs3b8bm+x9EuLwRg8MTGB4joyuMloZWvPKbf4I30Ycf//hZJAMtGOzvwuULx7FlyzqESqvgD9Ygnub8kTCgDAGYOdy6eQG3blxEXU0ZFnUsx8tv7sOJM5exfu1mdDS2oba2AoHykIB1/f3daGisxurVGzA4HAWtWJra2qRCzw1U7N67BUUllegdJlxUKkAFGXlcyN6JUcEWZxKMC/fJqQkEi4PyjLCin2MxWYaskOO4UFrCqvIQ4rEUZqZnRTKKBpRkL5D5Hi5mkk1lozgXkQnBsZJ9PR9QQfkgC1RY9iMXSkw+yDgeDEpCmowBJo/DPBefV6pKOR9GZkazgAqO4RwnOE7beYTjeWVVpWzvMCo8ZCZMyjzA/XP+sYwKzqcEcPj80KNCFoVuoEKSC94MUDEfl/FfJMagTAmOI04i3TAF3UCFw6iwQEVU2WvWo0KAerKCIvMisURPSl3oE2BRRgXflwS41y9m4zQHLykulnjCtrVdMC4EKrzo7VVGRWmJFmIoYwMyrwtQURySz9iWPbe7BYAvDoUwN0+gYlqAG8pB2blbddM9mJ0jqxTSp5hkIzND51AmXZRRoVXTmkjIBSpsUsSOYblABdkRjGNs+2peT6Us7Hdt4pbMH46kZBMyqVNconO8FA+Y77uBCiv9RMAhldTiA/apLEaFA1Sw7RVAIpBkWStVhlHxLwMqXDVWWYO0HfF/D0n+vKO/CaQLFCcV2iSn6qnw1+QTo/333xKo4OiTP69c+FTvtkkLJK4LXnweoKIQZpJZMxW4iAIbFiqms/vLT2LJvnC7a6MslL38EwbkwqhDat9MPJF7avmaVb4vXaFAo9tCuQUf5yQmsxaX2fu78+28y5t9B6CiMOHGlaQzmQuud9xm2vteettJDIuXh5Hn0bAoA1ToY+M6Z/Mrvd/yvqRwT5PZNkmrm2gFekZCxpVSsTsyx7EV7faR1Y/NXuR+a3Ld/dKCk/ynpAoMmgbP6qdZl7XwGs1ZO/1QGNq2VNUmoMWIOZNIdi5QJg9Vf5BtXMWNHP+lkMqdJzKwiVVksACSAAlZha/Z18hqdH7HWUsbPw7rT2mZD7Zx5Aky44eVZVJTbJVEyr3f6kOg60VxeTCJe3lGjdSTVq5rYl2BD5WC5X6l2p+JedO86llBQI1J84Cs98misvJFbD9bRGAlQ7lvYfQb7wOpvpcVmAIxApAQ5BSp4LiwTFl0onJCNJFWTyhenZWsEtNomjCLzJG5WU7Tah+2b2cKECAxCNfIvAYFLMyzw+Imk+TnblSGiYl9sn/U9FnayPhEaPtYhgVjK8tG0HvANR0bknkEfTZVpsrtUWGlnyQfxcIqA/AEjGk2j0sWHM9Xi0oNWOS3MlrqUSFMCAMsybHss2rYK3b/+uwYloiLOUpQQQtfFECwZuz2WePfEnNJsaGyfTKPvI4j4kkikrSGzeoGN1iATFWBJI20tT9RyUPa0Dxb1kfDsmLFIN287gEV+cfFe+/+AbfA3/xou5591kToZki4kvx2XDeTqFK9chL0eYGK3BnV2ZF9tLJAAPdEXTDazWIq5PdSkDjdRgquQdmCFM7Un3sNMmPnBgY5VbECLkgokA3mOGCGu9TIACEyeZsgxJFickKKgkuWQkG2mVp08WlAmqyWzroGc5+MOXZWgOFAVe4j8fdMcGYnHRnEDcVYJlhBy430kwUq5uclqcwErQAVkYjIQLESh3+3r1ouPgdsC5paUvon4A9Kgr2krFiSFEL5TCZF6oKJdibMWcleXl4pSWatVk3oz2QCldWVAGXZOcnH4hjo65MBvqmhET1dtwWoYHKd8kd0XOYE09SijIrZZByTU9OorKgSMEMnOK38j8ejhlGh7edmVLBa0Zppq/RTDbysEEEC8fmYnBuTRwwcbOWgm1GhQIVKP/mCxWLYymz5xEQ/vKk0SkJFSMwrUDE3My37DJeVYWhkAJcvXpDkJIGKknApOhctQQUZFX6fVK1mAxXzkrhjpQGTHWQD2MCX52MrAsSjwphaM2HFwImeFKNjY6IBzUpJ/q5ARYUEMUzCZoCKYRw++Ilo1lP6iUAFgSV2L95bAhVsBybeqbMv0lTGyFsojqaSk7IituKU7UNJKZ4v21qCzVRaJvCwYYtMTU3j/f3voaqmGhtozku/B1br+hkYEahQwysx05KEVwmqq6sdo9i5aARlxT4BHaYnI9IvmbxnRXEsnsDrr72F0rIK7H14Lxoam+EPBOVcqENBBtH4xCiuXL6MpoY61FVXo6qqEo31DRLAEAAbGB6Uvjs6MorXX34df/7DH2HNmvvgDwdV+onyTXH2NfWFEONRr0kqyTNCRsXbEoju3ctzaJDvsq/Ltkb6RCo/RAoliWgkhv37P0BnRxseemC7yJvQv2GacmtFNOtl8jpH+mluFrt3KaPCDR7xe2mvR4ykKe+0d89e1FRWKehESRHKuCQSuHzpkgAVu3bsFJBAmCnGTJt9l9JPrS3NWUAFr4FAxerVq4VRYSueHOmnRe1oaq5TUIRm2re6xbdm9Rp6VFByQYGKTRvXZxgVt7qlopvnwATbqVOnsGHDBmFUsC/odJfRh7XPQu5i0D2tF8zFCPDhmgVcAa3sz0hK5QsRZBHlYlLYvs3+X1tTi6AviKHBLhz+9B0sX9aO1rYOhMM1gK8U6RQXDXZRzXNQ0zqyp65dOyNgRX19A1pa2lBSUg6/jywlDxKUQzJMQqk34yJYVmEpGTejkSkMDFzH8GAvqsqrUM1/VUzCBzCLILpu30BsfgItTQ0I+MsQCjcC6RLMRqaQSEUQj88IW2J8agINTS2obWjGlfOXMDzUh2ee+RZCgQqMjUbw+bEj6O2/JMetrm3Hqvs24+aNG+i7cRXrVq/C2g3bkPSG0dc/LEu0olAJqsur8dqLvwBi3fjRD78DFHXi3Nnj6Ll9Edu2rEdZdT3gK8dcPKDAk5fXFMHwYA+uXj6HcNCLlcuX4NTpG3jp9bdRVFaJzes3o7OxDRUVpfCEA5iensTgQDeaWmqxcuV6DAwSbPeiuZXST6y4n8bM6ABuXj2GPXu3whMsweCoFykvmYBF4puj0k9JkVWwgAUBUz6r6sWgQMXcXNQBKpgIiUTmBJTgPwtUlBRrZT7BcDIq6KOQdoCKNEJhSnx5ZUzmWEmggot4Mioss8BS9TnGckwnsBlPpGRuEp8KAhWm0pSARWlJWNhgmignu8ODmakpNdOeHhXgQr0uYjKGcqyg34bdB78njAq/X8ZJqfDkvDapQAXnAT4b3I7bUMaJRQICVFy/LmM3qe7cNyUQPcYjigtyYVQYoIIShB4vF/UKVBRiVFByitdIUJX7FDbIvG5jGRV8PmnSTaCCc6Q/kGFUEKjg+MNtufDn+RKomJqaRHG4OItR4QYqRPqJrEaiHh4PevsGZSy3QIXGbQpEj8+QSRAWRgXvS19PL0JFQQT9QQEqIrMRuXelpTwHXfBrmOrBrFR3Eqig1IVH2FhkwnDnNCu1QIWtwtOFspU5yMR8NvliEzD8Ho9F4NsyKkTCQIY1k4hjjs/IbchxkhyUWNAwKgwcyuB8EVBhAQeOaW6gwoI9Y2OjUkxAxiP7noAVPpXX4rNBvxxlVBjpp98Lo0ITGAWLh/IM6F+YDF+wTaFM452Su3dzFANU3NX61F73l9+oIA5SoMDKyeJ92UP8C4CKgvetYLa70Ayf/yTzsd+/CA9asAp23sjjF+L4KGaflwIVZsmec2r5eo0DVORhYORZ5josDVthnRlonBHHDDyu5NsX3Md83aAg0KNVcHn3WGgbMlbtFhnwJ40f/S8/QU19Lc4cO413f/eO5iqcxKQa0WrdisZpdvxzjm92KgnrOwCKjtqCzYeYY2j+wRxDYYMMeOE0ZwaQyFx0vvdM3sCO+/mACgt85NzrDLCVPdZnTiG7vd3trEUwhn1rNrDsGxtDM2HLedFJfVhJHFvxbaSdbK91PzsiRxtPOEl2NhjHcjcLIisON4lyW0QgSXWTRJcWMvfRetFJFsMAPTaBbCv3s67TdX/JNuUrsx7Qwjhl/uucaIsyxJcwSIk4rsNYQGHlFFn9rnOs5DnMepJ5EcYXKjGlwAPndX6u6gtULlAmB9d7UoFv/scGtsUdtu9aAEQLIplAVw8DgVmM7wePY83BM23pmkfSZFyrP4a0CU3BDRPEtidjQO6fLwVimET3CyhhcxsEangvuaaVNjZxmbKomLjXZ0yfM/2OfVlZL16/wzrw+fDLf8zIV/3J92mQTVkvAi4K8EhC37Ap1MtE7wMbXQsiCJJlvEgEZGIEzT5HAMNIcStgZsdaXRuy/VnUw+eW91xVMZhHUBNtvlhoqOdARQPtN9Ycm38zj8JrkyJXs+bk9prvUDUU7Yc2j6j9lUCUZWxw/1wP6H7IOtHvu+N6/u2sY+95VHzBjHTv4z+4FnCACh2Zc+fKPIwKF5Ivk7ya72Qes9xAmpmazKdyAAPdOoGBTZQ7m9qJM2c7J6EuJ+t6uHUoz/aLMMHHAqDCXKJJ2C8AK7LKG9zNYYwDs5L69hzs+Zi92Z1KqZEbyHF9P0emStulwAKlEKPCsB2yEmzuXYi7tOsa5FSsSaRrysoCatz3z0ZqGeYIq+XyAxUJw6hQuaP8QIUyLFqWLxUNfyY5mRzg5EFdbCYnaCwqEhLUTk4kEJ2LiowSE+bU7S8rIyuiXBb3KlvBhNA8qmqrjEdFSmSf+nv7JFlSXVklJsZuRoUCFR6RfmpsbsJ0bA4zkVnU1dZLYl0nHk0YW6BCKphlge+XqgGhe6aV0ZFMUNOyGDU1VSLnlEjFhAnCydDqB1otZgmwjEk5GX7KqJhHuKQKjc3t4iEwMdEHhn3FrJqdj4n0U5ReANF5FJeXC1Bx5dJFSUJ0tnWitKQcHR2LUF5fK1UdTAYxYcmJrCjEiogoUiLDoIbWNAfVa9EkuRuoEBkNkyhSM+tp0U4XPUePV4AKJn7YtpRoYq0Hr5PJ1eGhIXx66LAkWZcuXYK6DiYAWdENAZ+YSGLgqxUaKaE4qryHJugt84QBAoNV9jPRXR8akt9ZOUqvBUuhLvIHEY8xuTSLd9/Zh6raGmzcvAnzUTUFZ2KDYIXq8GcWGxKE+P0oK1WZMWpul4Y9YuyciGmSjAAa247JxNdee0uqeR997DEBt1jdwEDTS+ZNIoax8RFhExSLdFQfWpoasXXLFmVtpFKYmJrE8Mgobt++jU8+/ESkn1avWQNvkJIgWvmh7B2T+GdwKl4n2lVYrfIOPSoCAWFU1NXXSbKR12SrlTS4o+4GaaqseCcAsB/trS3Y8cD9CAS1Gmbe6N4yJqOJHQELPocXzp/H/Owsdu3cmSX9pCfhQdJDRsUF9PX2Yveu3QJUWCZH2oAlly5elP3s3rlLPCrEA4SLCL9XQLZjx46ipblJgAqpwDGvffv2CVBBXX07J+R6VIghXgLoutUjgNKaNStE01yAihOnsGUTjaeplx/FjVvdYthLVgXPgdJPBCr4N1k4KpeXJ+GT85b7O6JxmjO724Wajv6uT201jRj1ZSqzc4MDbuGeIexMQXozz5WAYyI6j97u6zh/7jOsXr0EDY2tCAQqxdOGCypdV+g1KcOdXj/T6Oq6ipu3rqO2phKdHSoPR0mUtDeIBL0t5HnjnENPlBgmJ8cwNTGG+dgk/IEkystKUVlag+JgEdJxJqlnEPXU4LMjn6L79mU8sme3nEsqFUYgWCF9KBqdQTw+hatXz4uvRnQ+gYrqOowOjODGtUv41jNPY3R4Eteu9uB29w34AjF0Ll6CpSs3o7KmGQc//hijfbexbtUKLFu1HvNJvwAV1FKjR0xJMIxXX/wnpKK38Rc//TOkg4vx4QfvIBoZwto1y1Db1IqUtwxzcQWikaL+cj+uXDyDdDIu/W5qagavvXEA13v6UVVXhx3bHkR7XYN44CDkx/DIIEaGe9HcUoeVq9ajfyCC+fkAGltbJKk/OxPBxGAPum+dxiOPbEMcQQxP+JHylKK4JIiqyirQDDtX+knXNRzvKHGk1e9kVExMjgujgtgRgQjV51eggl2UQAX3RwNnyo9wXKLXCKWaEkkFKjiG5wIVfJZkgUP5GzOWcoyVqj0uigl+G+k78agw8n8i/RQKYmh4SBgRpWQMUFpqgn0gjkiEcwElrEIy/3KM4zPGOYUJfF4bxyIWBfC4PIYAFTzHySnxqODcwe+IcaXxcSguVonAmzdvSn9k1RrnKqkA5Hzk88u5U1aLrBL+TaYfE9YWtLVMDVttaYEAjutctLuBCgI+PIeS0hD8AZ0HGYtEZqIir6TvaVGGlY5SyUDOl/RtGBKggvOCBYQ0eaKLZ84vCsLoP77X0zeoZtrFJZqMkSSLju8TEUo/0Ti9WMDV3u4ekVak9xKBCrJfeP1ZjAqlRshcxIU7YyVyNByPCpf0k00QZBIFxoMjy9DTeliYSlFjLsn5X/w4yst1cSwLbB3NtBrUeN+IHIHqOiujQv2btABBPSpszGGBEhsXSf8zQIXjjWLabmJiHDORaQHHOP9zEc+mZqKB36X0ExMHodTvU/rp7iWTCiWqC0vf3gGQKJhQv1ugwllw5U4/Bf7+HxCoKAQYFWo+E19ngRXOkrLQRncHVEjfzzG0/u8FVBS6kRmfRdfazqwrZSWd59Lz1RVqj1lo1i17tf3SXSV8h55VCKuSU8nXx/+/ABVWztJU8//oP/x4IVBhijPkmTRJWXmiXECFgjsOSqGV9QWAClnRG2DCKdx0ARWKXXgdkWkWS2k7uhrNZb688MPM95wiR/OWc045fbvQvXb2ZC/NAht57oONwzn/WqAiA2QruC5yNYz9aYhsYgyZkkQaUBPSFiSXudHV2Wz7SmLdpHk4l7A4zCaqc7uVrbG0ILkkzA0Dg8fXKnmur1VCiMfOVO6TUJ+RPGURleauMjfCnpOYLRtfUDmGSBTpOtmy7UV+2JF60s9kHnaZetu5zgIVGg9FVQLKMEEYU7GtrCE2YyllTOq6wWG10/zZr+oH/JzFeVzviVeCqcwX2SxhTapHBwu6WFzI+VLXWwqASGI8txBXSEWa/JfzFjknFofRj8HkkUxBrG0n7scySOx5StsndC3KdbRVTBAww4Aw7ljExg42B6ESTbxvjFu9+MU/ZGSV/vSHMSdPoLJRumJioaswMiX+MACKyWMwdo7Os8BR4zYhT1kmqDBXVKpJASUDUFEulusjP9fl+rzyOvieqG2I5wTb3RqhZ0ATPXdlysp2RhbKFtY6MblZM2cBbk7ekL40WghkxyjeZ2FUCAioqVo9J4JgcQN66DHvMSq+ZKhz72t/OC3w14ZRkZ2wt5RBtyxTJgmvk7xBnE01Qk5o5J6FDVBh38rIROm4YBc9dv82fePehf3MeZKzGjizEMgE8Yopu46Zs4Ub88h4QLgXAdkJe2cS06HA/HPGEedvB0AxVWduVN6egsRHWSdgjvUvACoyrBYTbLnOREt9M9chVOLcdY5hpujb+RZBuYCPHdB1MZthVBQCKmY1GS+MCgUqGpcsksU/JQ+8XpqFFknFJZMz/iK/VCF+GaDC+lRwQCdQ4Q1o1fzYyAioD8oKbVbd38gHVFAeo7kVdfX1GJudkqRfQ32DU9mZD6hQhD7jUUGggtdEAN8CFQE/z4EAx7zIWTFRYyc5t/QTVw3qUcFqyRhKy2vQ0NQmCSRKP9EmN0wTtei8ABXxKI1U51BcVo7BYTIqzksioLN9kQNUVDXWS4UlE5wEd3g8Jj8YsCwEKjISEFrFQTPOqPojGKCCIML09AxGR9RMm8khJn2o2U1GApNlXtGmtEDFMD795JAkWRcvXYKGjnZUUQKIAU2AbBgCFUykMrFCaqsalLrZAfw8KECQAmJsv4H+fgWkYjH4HTqsV3S4Y9GoBG0fvPc+qmtqsHX7NgEnCIQRsKBESoDm54YeqkGYjg38nQFOSQk9LkKSeKLkF5OJTAiqhFYUL7/yupi9Pvb442huaYPPTzOrBHwMDFMJjBKouHIFAZ9XfChKikO4b/UaLFq8WAJ4ym/09g/g0oVLOHLoCP7NT/8CK1euhDfEytAcoMIYtTk4ppHW2vf2Pgk+d+1ymWkboMIyKhSo0ERhOuHBu+++j6aGegeo4BhmgQr2b2JvBP8YAFH6SYCKXRmgwgaRzAqlXEDFrp27BKiQvsJA3hjIEaw5c/o0Hnpgh0jPMKCbZ+BsgIrjxz8XRsXiRYskoLeBoQUqaKZtF0O50k9iMh5Po+tWtwBva9auFIP76GwMJ47RLHu9tHs8MY9rN7qkL7Afsk+7gYqQBKtmtMtZRZvpKO/krTUs2S9nP7oEcD601yUjqgTBmQpo9x7yAxU6MxCMLasqgTdZhPR8GufPfoah4ctYs3YFKsrr4AvRa4dBPPfNZ4VmbhasoHTZPPoHbuPC2RMoLw9jxfLlKCsth88fRkqAjTTm5+fEQHtmZlKeldISeiyEUFpeIjJ78Tng0rkLoIR3Q0MpUkUNGBsZxxuvvYKa6krseOghVNXW0kkPyRSNHueBdBSXLp1FW1sLZmZjmJ6eR0VJGY4f/xSdnS3o7e3H1HhUvIhWre5Ee+dyBIubkfYV49AnH2FmpB/r1ixH26LliMQoFzQrJoLVNXUo8gfw8vP/gNR8F/7yL59DNN2GE8cOY3ToJlYsb0dzx2J4/GRU+OClLNjsOC6cO47I1CiWLFkMf7AEn31+CocOnUTC40NjWzO2b9qMZvptsF8UBdA/2Iex0X40t9Vh2bK16B8k+FKEppYW8QKYi8xirP+2ABWPP/4A5lM+jEwGkYR6VFRUViIYIFBBth/BRwVmaf7Ll3oxKFAhRpZTEwiEqTNkgYoQioJhp1rKAhWUfiKQQQAvlVZDQvWoUEYFwWPORX19fTJWN7e0OPJCViqIzzMBBo4XMfo4GaCCQLMFKopCQZSGQxgcHEBJOCwADsfqaTEvjWMuOoVgkV/ej8WVUcFnjPN5MEA9YWVKWDNtAfLNyooeHARiKAvFsdcuyrmA5PhqgQqbvOb8Q3ZcWmT4KA+lIA7HaI7pBM09XtV/5jNHoMICMzZJwH2Kl4Uxf+Y+VQebsUtSpImCQU2+z0boRzKPkhICFbp45XbiR5RKCSijuS1NxEciMzJX2HndMgfcQIWwBjm/ej3o7hnIABWsMuQYaBIhEzOUflKggvFMd9dtASq45J2bj2IuqpWYAqIIq0HPj0mVOWHFsOgjKsCG20ybDDsLJjjjkqgg5mdU2HnXjl3c1gIVZJtaRoUNFd37lgSELKKtRwXNtGlenu1p4QaS8gEVbDP2UwvyjE+MI2KACj5HTGBYjwoCFVXVFfeAikKzlmaE72JBWvi7hQCXQh56BQ9qdVG+9Fnlm33vcFn/nYAKS6j/0tBRofVd3ibX9Lib1S7P5B1vpWXs56zGTZHFF3layFZmiZi93nWvxZ0sdybeucN9lLbJ00DuGCl7c/VyyPcqtI2U0RmAQ2IyE9f98N//KANUvLTPOQ2yFxd830oIGdaF++KcivYC1+kAFRxTbbe0YIXEgPo+/0kyVQzo83hSupPmC5pA38hqA1dy1eZkssCf3H24/nbvp1C78n0LLmtFucouyXkQIJBCtwydWMEJ875ZE9jvL1B8MOfCYjunMpwm7vQsJEPDmBXndp9MW6sfHEEELUhXGWrrV6FSUwpmc30q1yhsfD0/K/2TNTra9ufa02XurQliFr/o2kqln7QzCJAj7IeMcbQmvSnrY9bGwSInzyUeBlLFTyYJi+nIpmDRGddiHiQZy4gXhko/8YsSV7Ag0MhM8bhWMlHPQX0l+H2b6LdABXsdYydpR7knRvopZ7HDsUykuLm+NqbZTJZbwEJiFdP/NOfEAgs1IRcGhgFuNNbVpLqssY1/hUh9Gp8IG7tkkvSZtRPbU/Msqobwq59lzLS/+2P6Oei6kX3NmnXrfjwSTypTQ9mWWjSjklxamKUm3NIHLJhlmAn2wbX3TsEpja8suEHQgs+ZZbRmgA1tW+2ber/4N9tAABp7XANi2OeYn9kiIit1ZYEkslcIpkk8Zq7V9ml7L/kdlcBi/9T+KMPfPUbFHWakex/9QbbA3/xwu8vvOTui0AnVbdRsjaFdM55hVOSPWvh9a1xtv+FKnEv1lXm5kkbptE4ymZdNLJlzsYOsYQfYAUJ3kQlUFA7IH0bKkOJRDb0sw+usyd0yEgyE6QT8rjYxXktybLcclRzW7qwQAJI7Dd9lF3JknOx+bIWt+XtBZs1Guq7zyXu9uW1vgyrdziLyYqBEkyTq9dFnQqSfYlJZQEaFSj3NilG1ghQKVFQ1N2M6MqPSP0xucJAXwN+DYIgG0GRU6CRfkFFhpHKI3gtQUVMpjAoO/r09PRIELFm8VH7euHYNUy6PCpZhipl2UwtqamsxNDUmOo/19Y0O9TIbqLALcC6SWSWglSTUjeR1xeZZqVqM6uoqBANEudkW85JAmZubdXQi7QTGvse5lQtubaMEyqtqUd/YLkZR4lGRSEiFPkGKJM1P4zFEZ2cRKi3D4FC/AhWJODo7FKho71iEmqYGB6ggqMFzJGghlFWpblTpJ1a/2iQrz8kmPphwsiZUVnpjZjoibAAm8pg4GJ+YEFkHJoEpXcWQi4EWP6dExKeffILamhosWrIEjZ2d0r62EoGJJD4TyoQhRdQjyR83o4LfJbWTgRZfTBIRqBATbga1DBJNRQQTlwRkxscn8NGHB0aqMFoAACAASURBVFBdW4P7H9iO2ppqASMGB/oxMNiPUknmGTqtqXS1QRKPURQMoKwkIMkP9idtMwUsWAHz0kuvSILxK1/9KppbWuERSm5KJcp8EEbF1StX4EklpRJW/EVKSrB61Sq0drSLHNfE5BTOnj6LD979AH/xk59g3X33wVPEwFDpp8qo4DXSCJyLGSNRxECUhtP79kvAs5NshYY6ed54jVLRZAIi0Rn1qJltKg68996HaG5sEKDCbxkVMa0gEanTXOmnSAS7jJm2W/qJSbZ4OimyTjTTJmOiuqpaqb0MGg3wQ+mekydO4IH7t6O1pVUCqJm5eUnSseqKQEVba4sAFc7igYaChlFBoMIGYQT5jolHRQeamuplAcRn8tbNbkSjc7jvvlVg48/PxXHs82Mi/VRawiRsDFdv3EJVdTXq6uokeD1x4oTDqAgFaKZtZoZcoCJnqnAv4IT5kKc8UIJZWfga/VOziODzx/GxlOAAAQW7byv5JwtVCABkZxl+ReWYaPIbRlV9KXzpMvhixZidGcaZM+8hkZrA8hWrEC6rhS9QLJJOHg+p0KR9M6hlwKzsGSCK8bE+nDzxKVgAtGrlKlSUVyOZ9mF0ZBiTk/QbgBiB1tRUozgU4BJJWF3JFHX0Qvjko08wNd6HrVuWoaiyDumEF4c/OYLRoWGEy0LY/fADKC4PYz7mQzKehM+TwMXzZ9VTI1SGs2cvI+jz4cbNS4jMjkvF9bIla0VjfsnSFjQ1L0UiVYWUrwiHD32EuakhbFi7Ao1tnZiYjiESUS1hSq/5PV68+sLPgdht/OQn38XodDX6em/hysVjWLqkBUtWroIvWIlo3C9yQWdOHsHI4G20tTaiqaUdZy/cxOGjp3DrRi8q6+rQsawTa5cvR11ZhUjswO9Hb+9tTE4OClCxeMlqDAzNIpEIqURgNCrJ/dHeW+i5dRpf/eoOAUXGZooQT4dQUV4i0oIEKjjGcfy3zAomWHm/i41pNP0QKCs3OTkBf1j7B+WTRJ8/GBJAnEmA4rAaDcfjBCpmhfFFHxouwBm9WDNtAhVSid/TI+MSvZckaW8Yc5aOLjJSnDuTKv2kwDS9KVjRnpaq9eKQHyPDQzKGEQzmeEQgQubjeQIVNL+mYXhcZQzm6LUx6QAVvHYmtXksy6gggM4xUKR6xHC8SM5Xk9Y+GWu5yCSjgsfj/MOkvCziE2q4zGPSv4OMCs4RBM09HjXJ5vWRIecGKuyCksB6LlBBRgUXxQQqyBDhOEqPEAUqQjIX8MXtrM8G2QwqOZAWsJ5zuwUqbPKdc78bqLBeC+zD3T39SCWSso3KFyh7kdc7OTvpmGkTOKIXEAs4LFBBk0jOlQQhJEFkxn7OHwTQOHfQ4JT3mwCHlX6iPCVjIo7FNhy1VX3sj5JAM+O3nVczIbnGU6Nj45ibnUVFZYVqSLtAWQtmO1WSknPwipk2Y6DSMgIVTBpkklyWgcJv2oSLalN7xAPLMioYH3JbN6NC4iayJI2ZNp+XiiqOsV6Ef++MCtsStqVsTO8M5k4WNotRlxPG3ynBWijiL5zI/dJpcVsmfneLisK0kCwz3uwVwt2c0x2Y4wWT8IU+yCOZJAFEAWBDFy8F2uNu33fVgOVTHs53lN8XUFGQppAPETB9Nl/VfA7Wk7W16/vu9zP90p31/qIudkd0JXtjzTrn3SHnp4UvZX5I7JtHUkb9IzRJnUmWG519+/RacML6VtjH3DBL9M/855TZ1LDRXECFZTyIY51NZNp2dXaXXWapby9sW8umcLe/JGDlq0blIochoe3iajGXv0n+7pl9jZrM1VyM+CQYNoh6NarkDtcmNEy2HgV2HrByx0yMM1GeuezsZ1ZAIEkiq4wQXyIpJB6Dej5Z/c9IOfE4FlTXwk8j8cQZ03j+cVtlGWh8oI9/Wj0FVDc109KuhqI3AD8RA2TxCiCAoqx8rgdZLMG20AJE3Q/XHZSv5ncEfKcUltcnRVUsxLDH5rwtxtiUuGLFvvVK4H5M0a+VNZJ2NetBr98j6zV+RqktzpGifkBfMZHtzPg6aHtyLRtXcEH8JCipZaWk3H0ik+HOSInrepTrFhabSRzleoaUUalrOgGwDFDCY9rCBcsksICPAy4YQMf6ZQnQZeIA7keKVs3f/Pn8z/Vvvr774/+XvTftkuu6rgR3zEPGlHMmkAASiZEjwEGkiIkQKVll9fLXtkslWbZ6ddnVvVz+F3b/g/7gVdXLbZelLrfktlQ2xVmcBwAEAQIEMWdiyHmKeY7otc+5970XkREgwXLbVi+kFgUg8sV79913373nnn323jUjM84EfkDYNwpOqISSgmks5DGyT5TjEvaD5hLU64UZC6p1qPSSMoE0hyXjXAohdZwoMKAeFApa8Hw1ZdYY0IjnU2aPPgfxEDE/MkbN81bwRQFLAUuMZLY1ndexyuIVAlLK4uC5BOChnJbpJysVpedW9pC+l26u8QFQ4RnfD/76/48e+N/+4FnPSuCRCupYs9zAfEulRUfQZOsGbN/Ia+mWaThd5ia8NXiwAIiRxelnXGUrQ5z6BDZS2+xuJQxQIb/qbo8zhRgzV6PrZihkbjmEPc72B6s8mATUzy2irBf2ACNdvhltx2XOZTZ0Jrs8JuRm2XS78ysG/71iU1l0TWDW8zS2v3mUG+x478X7xJ3+FWiZJm96372ACoIUIpFhTLQ7zLSNZ0WYckB+H2IDCfGLkIdH3T0u3uGgmE2hpV4G9Kdg0o8V8v5AEKnBDOLJpCRny+WqJK+ozTyUScnmlRr81Olmsnn37j1iejx34zpyq8tS7WrNtDnB00ybMknr5TyGh0cwNDhsFjVWhWoQQHaEDSZkITOJH0W6W5IcYAKVsheUtKCuNxe+Wl2TQNZkVKiEBmnnRl9NmAIi+1QsVjE0PomhsQkxxcptLnCVEumnZrWOdr2OUiEv0k/hZAIb66u4/PlFYUns3LEL8YEkdu/Zi6GxcVMlOiB9xuuJDFSNlMmG6EUzmcM2edF/Loa8HyaO2JeWGslqWUpiLa+sIELd52BQKkkL+QLGxkbVOM2nxl+RUBDrq+v44J13pS9n9pBRMSXm05rMaCOdoXSEXxgVqvcYELCKPxbM4LEMQBgw8HrUNV+Ynzc65E2t0GBf+vyawKtVsbqyhjdffwMjoyN49shzwpKhZAmD5LWVFdy5e1dpsGSpxGNS4cqgTRZ6QgIS5LBSgpXCEWFSsB0En5ik+vnP/w6RWAzf/a3fEpaEDbpI1+U7ns1vYnZ2TkC1xYVF9SYpVTA8nMGTTx3GuPRBG5cvXcZP/+an+NHv/whPPf00ghFlVFhzN0sDZiW2JKIMK4xB6OuvvS4J6GPHjmFyctSzafBJMGkrtej9IRJPlSbefOMtbB+fwHNHnhGPCh5DfXc1+dIgh8l+BmQXL15EpZQXoMJrpm0mPPEJ+OLSF5JAe/755zGSUfkWBmwNE8TN3riBUx+fwtHnjgibiQEt2S5knTCZ+enZT7B9ajv2zOzRucNUN/3qpZfEXHyaAAYriRjc1Rs4feoUZmZ2Y2JywgFEb964KdXFjz3+MHztgEg/fXLmEzz15GHEYqSN13Dtxi1JhtKTgolSC1SMjY3pOyhLg6lItpObgAb9a08l4DfAtgStHu8J6ruyspvJquzGGm7P3USpkBONeZpiDw6Oi6cLAdiWABTcWITg91G7nsCR6snSr0HjUd20TGwbQyQ0gEArhFajJqDDqVM0q89gemZKjIADwSiCgTSqNbLSKEFE8EgBCx/qQKuMWiWLjz96B/VaSQyp69Um/OEWBkeTGB0bRiQaF9PsWoU229ycKUuDwAdl1X75y19gMB3D44cnZN69e3cTA7ExnP30PIbHEzjx/BNAKyAMMiaOL1y8iH37DmBkZBIffHAKN69+jkJhVfx1vvnNb2FoeApnPvkYhw/vw9j4LjRbnBeA11/5BwR9bTz22OMYHp3E+kZeWASJdEokjoLtEP7ub/8KbQNUfPbFJpKDQ7h583OE2hU8efhxBMJp1NoR3Lj6KS5/cQHj46PYd+Ah3Lqzgs+/uIUzZy6gXChg29QE9u47IKBZKkmmSVAS/3dnryFfWMX2XRPYMX0QC4sV+P0JjE+MoVgpolSuYfn2dSzOn8Zvf/d55ApJrOUDQCiATCqNdCojawHnG2VVELCowx/ihqKNmPGoqAijoirvhy+sJoIEgVOJhMxrOjcB8QST8xF5xyn9pP4+SrnnmEwkkjIfMXHO69yam5P5a3xiUtZLm7i31ZFims13tl2XtUtYiWRUkMVGL6FIFMlIQEBerqFMeKsHRUGS3eVKQdYRSolxvVDPiJrch5UH5H1xvLPd1veIyLx4VMTjSCYTsnln3+h3OC/H4fcFcfPGHBoNTRJE46TzUwNZTRpV+ikiYD5lB8n0U0YFBeZ88q4xia0+Bn7hGvFdpccE51/eJwFnbghFOo8m8fG4gDHciJfr6uGTSMQFhOf8wuQ5ASSABt8sUmBsQJbBugCmXCO84AgT8jZG8Eo/cUN85/Zdmd/YZ1z3uH5K/7eaKBTyiA7EMeBhVMRp3k2fj2oJuUJB7p9Aha20tKyRaqMmY6JCRgUoQxlFlOdnRSE35aYS1mFhOFIH3XsYjYe1OFljFGGorq3KWE2mkgiHtIrPSfpxQ8+iA7MuC6nPHxRpLBtzWKDCShdYUIdXt0CF9AeBitU1Ac2UPRORDTpBskJBQS5b4EGgk/0rQEUmLQmHWHNEQD5K3InpuQB1CkJJ3O7Zq/QCnbfu6Oyuwk0CuDuN7s+0zzr3IuaMlsG3Jdd5j6Ts/W4v7zsB3+8C95FUdrdT99va3sf3TeQbg17TNNlmuRu+3ue6B+DS8zm3tWJY93eeHztmurul3/asl0SkJyndq7Hur03SXQYR38UtaWsvhV/balRcvCbb3WO945odOXDDRPDern0GJsbZ0t4+/aoGzj161iTSO7r0y0aL0LK2jkN9vVxJKne4mByD8/TsQOm+kA4ar+yTc4RMepqgZGzoDG3PmHQqqB0LT3ce3HIlc9/eYWqBFMbomrDwecx2zVxgaDru3VsQQu/dDA0ZG1QB4FrOeVE8mJiUDQU8JJxOUMB6mklhlEmQb3kU3ndQGAgu89leW56B12/T7S35G32K2A7xyiuXkeB+XZKtusdk7MK5WWN9TQJbHwnZK0oFucoyWYDBFtPx31xvtFjSnXPVn0F9qNTfkIwGlfdSCUd9tnbe5zl4nLA9ZT+gFfy2ot+V/uqEqHhv1iSZe2vu+SRpXyeTIKgMekr2iIk0k8w12cepkbQmyLkPsNcne0Rkpfg9Mg7ED0T7hPE0Yw5hJ4jisVbFuuNQY0ph15Ihb+SKOEq4L6avJPeSUjghAIFP5EYZI3H9Frkq+lpxPmU8aZ+FgDCa3Of92XiK9811WhP4ambNflVlgghKxaJblGkMrO2+1OAcAjSorBNBHOYBjOyoiSg06a7yjuVSET/7acoZXd//AzK22wY84f5dvREJEEmBYzgkQJK018TPClCqxDb362L2LYV9lLiifpKybBSoMHtCkw+0cRPba2Mtto9MdMYnyvJXVonkTOw1O9RSlFFVp2+muabrw+HMMp7X0Err32sd9njdWs8Q+q3FYyiWSg8YFV+2vjz4/W9eDwhQ4fy46KoLxXdHZN7g2nO8u46as7mpbid+6Nk9XqDCJND7mqd5X15vu7xeDPbzrrZ5GyGLsWucozO1Ob5j/2GZEwpUeOgfXXfiAUecIKfrGh3hb1cb3aioO0q+94Dqi2V4wqPOqFvPRyaL53PVNuV3vLW9nTxjPaM1I9PDewIV9ap6VLA60TAoHOknA1REMsPwBfyIMcnCwJHgB4GKFhCKBKQilAZp1LVnAMAFix4VDAIEqEilZJHkNUI+VlVXMUigIgCsrq1jaWkZYxMTmJragWyOQMU1ZFcWFajIZIxkCrBtaqdUbhabVUxMbkNiQKUj2A9cgGShQlMTTZ7Nrk3sW6BCF9uIyCFFwzEJhKu1kiSrCApwcRcKoKnQ0CSAykiVSjUUilWMbptCmhXglbJUMHO8xSJhNCoVtGsNFPOUyqoimk6JXMvlixfRqtexc6cFKvZheHxMAi/6LrAC0gtUsLoiGo8ilUq6QIWRDrL3w+fGpJOwHcTrIi7SVGRKEDwga2JldVVkQAhUSFBKSmqjKdr/GwQq3n0Xw0PDAlRMTu8U0IAJKXafAhVK0eTrxOt6KZrWjJWBt03+MEHGKmF+x1bDCGWSvibUbq/VRKv89Vdexcj4GJ47ckRYHOIPQdAjHJZk2a1bc1henJfghBUSNDRlMofBhQYhSt3k31lVzKoZVhSTffKzn/8MsYEBfO+3fxs7d+1yaKNMGtETIpfPYW5uTjw0NjezMnbI8mg0qti/bwaHDx2WBMqli5fwN3/9E/zgB/8OzzzzDAIRrQIRVgQTVoaiLIk3E6zbCt433vi1TMnHjx/H+PiwAhUm4eSyH5h6Y0U8350W3nj919g+MYHnnnOBiho17o1Eh1YksXqGHhUXUC7l8fzJ553xyv6ToJibEl8bly5dwq25Wzj5/EmMGJ15vocNU3FCRsWpjz7GsaNHsXPHTrmvQlFlUxhAkW2xfft2zMzMaBUK336/Hy+99BIOHDggn/OaUsnVaOD0x6ewe/du+Q7bwftkxTU9Kh5+9KAkEin9dObMJ45HBfvcC1Rw3Jw5cwaHDh0ShkWAcmUmIHVmO7OfE9PwHjOurngK0NrveoGKBhmAfoINDUm0f/bpWXz0wbuY2b1LALN4LCreO+mhNEZGxhCNpYQB0Wj4EfBFzMZEAVu3Ys6HkYmkGvuSMUEqcruJW7eu4fSpD3Do8H4kUhEMj4wDbbKSYmgLUMHgnyeiJitd/KrY3FjAyspdrK8tYmgwjdGRYaQHEwIK1xsEGsNAi14trF5SnV+uCba4kUnZv/iL/x0nj+7F5LYR1Js+jIzOYG2thFde+UfsOzCFF54/IhuVXG4TV65fx+S2HdjYKOCz8xdR2FzBjh0TOPL8cYyN7UYu38Dbb7+FZ559GKPjO9FGCuVCFm+98TLSyQE8fugJDCSGZO7OZTeQGhpENJaEvxnA3/3tX6NVmcP//O+/j4tXs/CHY7h95zpQy+IZsmoyY7g2t4zPPnlb5HuePXIU6xtFXL02j9t31oThEfK3sG/vbszs3YfJyW2IxOJONdudG5dRKKxjamYbJncewNISZQgIVIygUC6gXGlgYe4qlhdP4bf/zUlsZtPYKAbhC/nEfDyVSkuSlOOO7zPlDeljw4o47pstUEHAkJt2Ju/5HFg9x4Q6gWQyxVQX2CcsuFAkLEzFfLYgLAytxtONJMFkB6io1WQe4gZ6bHxCZQqZuCf7giwZrlPhkEoSEKgol8VA3XoM8XysaEuG/FhYmJexx+Q4v8d1TIGKogNUcFNIjwZudglUcK7lO897J6OC/SDSiEwsgIBBVu6Hv7PVgEw081ZlLkUAN6/flvHLzXeUwGOrhkZLNaDZFh7PdvPcBM1DAhxoJWa39BOhHM7vFqjgcbGoMdNu1BSoiMVBryPZlNeryBXzSAzEEZLEApPyfgFpxMA8qs+J8lu8NoEKgg52E6vzqVZadntU8He3b9+VeU9NuV15APZPLp8X6Sey/9h/lH5iO7juliplZIs5A9TQUFqrO/W6AQhQQRC65PGooB8NEyMEA/oCFb03w7YqlufnedcEqKggmUqIcWi70QlU8BhJNomMFdvlAhVkhrEvCFrwffD2lVSrsvo0GFR2YhsKVIRcUIrHqP8KPSo4V6pJKRkvbAvHQyqdlH6ItUb/iYGK+9nP2aRaZ59KmP0AqOjoyF6jTncg+pstOWq7EN3P47hPoELX3S7jas+z2xIY3AdQYZvt6wPEeIEKZyvocGp7gBX9+sEkb7XZX6HQTeIeI51jd+1fAlSIfPDW3a8WLXWDPE5Ff493ou+ztPmFHkCFYxvjJuxNZNbJQjDt6DeetpzZLffX8eftOifB3RmbabCmN6GHd/a3TbDrEe4VJXFrmQImftckfWeHuHFgl9xTF5Cg1ex2P2k8F7w36Dleir3Nnk/ibLOn9V6rm4Jh1wI7nvTYzh50L2EkeWw+xUj0WMYFP3Yq9E23qKyNyg3ZNcSeX+NQY+ZtrmpjcSnDtNJP5lnYPZFdH5kUt4wHrhnSatN0/VzfE6l0N0A79752LvAeL9c1beX6ZPMD/FPYrVKgoGCArfAXo2n6boSV/cDiOLvHoz+gHRq2gIDtEA+MekOS6vKMCC7UqvAxoe5IBxkPKTNoFIRROS6u9dIeua7KLVnAxxoyE4QQ/wPzI/djis44bq0MqC0etGwDScpTxpFAFMEOw0xR6VAFRRzJLJPXsX0sBtTyDIyviFFikUI9aBwg7AYjc8Q2lMtF/OT/ZFyoP//298tmjGhRochYGaN3YY0yDxFxzbdNxkqAJTmexwhgpmboCnrVJe3l+haqTKU+R1ciTIoTOUblhiizpV4cmhcycujOa+EBOg0LxgImdl5gLMo+03nDfZ/cd7F3bOadJewRWjip/i5SDPJA+qnv6vLgF7+hPfDnP3rGabkb3LjGMu47ZBP/XFC6b9ab9fb+zhN+2q97F3V96z2MCvPdvkCF+b1zOc+EICkk74+HDbEFJOhebHsBFR4wQSpejbntFgaJvWan5JRarXVPNh4pqg4zI3stz/FfIc7so2rlBk1b+snbHhNe2coIiTbce3YCE1vFYcMxG5+ZiVuln5qoNzShz82+mmnTe4GyRvyThtGu9FNsaEz0/SPxATGVEpYGtbdZHRBRA2guaaxGYCKaCbBN6lEboGKAiQ6RZFCggtXaQ2nKCjWxsLAk19q+Y6dU9mdzeczeuIacB6jwi8wAsH1qpxoKR0OYmJgUsEHBhMB9AxXBYFikn6LhuBpG1wlUULrEC1SwIpOyLLoQMnAol+sCVEzumMbA4CAqrJ5cd4GKOiVkqnUU81lJesUHM1hfW8EXFz5Dm4yKndOGUbEPIxNkVLSkgoVAhYINmvhoNmqIxKJIp1OOlIUk/k1Shceyvdb0yX6X0lQrK6uyCFpdcAIVIyPDzqsrZlaUN1rbFKCCskC7Z3Zjx54ZAYwokcGFnVW2XNeZoGMi1AUqlGapVZWUH9HnYCtw5mZnpc2S5LAGZgaoYEKbSaPXCFSMjeKbzz0ngBHvW6t+tAqEz2RteRHzC/NyfVbRklnB+2JSUGigBjDgG802MKHE8/8/v/h7GZO/8zu/I0wB/jAwYDDJeCtfzEklc7lCJkVZkomUxypKFWwYDx04iN27Z3Dj6k389Cc/wb/9ve/j2W8SqNA+4DOwldc8twQbtqpI9EpbePXV12XMUPppYkKBCvuOWkaFbjsZrDbEN+W1V9/A1OSkA1SwLyhppUG3VsL0AyrYBmdT1QuoGFLpJy9Qcf3aNQEqThw7jqkdO6RfmVRUZkVOmA3btm0T8EGCRlahBPx45ZVXhFHBvrVABSVSyKjoBiqYiK3Wyjj4yAH420FQQufM6U/w9BOHNLHZrOHq9bkORgWBiieffFIYFgRINTT2mOv9dwIVUoouGG5LJNY219fwxiu/wvLSImLRIIaGo8hkkkgPJkUKJZlKI5MZxkBiEL42K4ZYXa0+E742A21NQieHaCJNuZWIVEz5fQzMa/j07Bncmr2Eo8eeEuAlMTDGo0E+RAtVh41G5tXSwm0066wmCmB8ZAiDw0m0A5rs5twTDqcQDg4DrSToG9cKaoWVVUzQIBy4dvUyfvm3/xknv/UUxieHMTi0DcmBCXx24SreeP1VfOMb+/Hss0+K58Lps2exvLKGYr4q97Jrajs2syt45PFH8cgj38DmZhVvv/Umjh4/jMzQFOBL4dbNKzh75kNsGx/DI48dRhtBYf8QeGKleTyRFq+On/3XvxKg4o/++AfIVuJYyxZx4eKn8NfzePbJxxBNDOKlNz9Au5HDE4cfRyyexoUL15DN1nH58hxu3V5EJhXFww/vx9SOnRgZGUWYfgt859rAretfoFrNYde+nRibnMHSMtlNTPwPo1ApoFJpYv7mFawun8F3v/s8NjaTyFVi8IXayKQGpaq/F1ARCHHeV6CC7y3vjXMrgYpQVE0H+Y4wcU7Q11aCDyQJVESUfbGZd4AKO1cSTLBABY+ZvXlT5KdGx8b7AhXCqGgZoIKbaeNRwfsnC2gg7Be5Pc5/nAd5fpU/aqJc5ViKIB5LSPstUEH/CS9QYT0qLFDBDRqln3hOa6bNOYaJZs6hBPM4F924fkvYQF6gglJlsh4Z4ITnFKBiZUWkFu2mm+e28ymPpy0ImXcq/QTZSFN6i+2sNapSaBGPxhAOqG+NA1QQHCKQ0CZQ4ROfJviaYhAfCrN6sS2AfcVIP7nJDs4qyhS0bEHLqmB75ucXpA0EVPgdW4nHZALBlEg86gAVlBC00lvFagkb2Q0BeUQOidWjxkhTpJ9qFZmra5Uay0ilsi4WjjpEVTLa7LzqZVV0ROqeuNbO+5o4aWJ9fc0BKmRz7VEacBJZTDa0GkJLI1BBVivnQ7JTmKjqBVTY9Zb9IOMMhlFhmBIKTOjaUSqpVCgLHaTYwAtUpJICSEXbD4CKrdvQL094dH7nfo/fkrf80p1wryvcE6iQbUmfdvX8eGsy1WnUPY+/x71v3cr1vs8+YIQcfI/fOad3jjFgoFIl9Otf1rNfE6jwNs277extvr21FfLsupL9blN7sDbueR/22W29jtTMuB1lkwXG6Lrz+HsNme7nIN+0slLi39OZz/BW13vHkfeeu7frUvTS0ST9h7LLNUFu/5NEcC8GiQcMcdugI8Ge2+4dZM3xq0+YSvXYlrqN4C1yjy17UALKkvx2R5Zn6JlrWDktbauOEwNsdaQsPIlWjzyXMD8p41S3JsBqdmyNr8XrwSnIojG0rwXZdAAAIABJREFUGjjrmsKKd2MU7ZGBUqxFtZ4ssGFBDnvHDuBhwA/bd16jZtlHWhaQh3iie0bD0PGyo8gcIAtEwHZlg2ifsNhMk9viKmO9DXxklJDNoMUEjFmiUa5n/C73YG5OiQG3MC1CmpdgO1kox+IAGSPcNBODMvJQ4ksghtXqS+H6KejfuUarRBFLNXQeqVTp76jeGnbd1bhFxw3BkECYEl2a9LbghIhoSFGhsgbkHpmnMYxYeXXkmlRBMAUUJqek/W28MYyqAveCmvRXI3BhbZpCCrKaeS7+8FwEen76Vx6g4kdls3NTSTLui+W6BJpYIFOpSiGOV6KMz1IKt0QNQ5+X/eH3uWO2vhwOI0UMqnX/S4CDLAy2Wd9da9Cu+S6qf/BdknHjjP1uoEJ9UaSvWpYNrf3sBfncN/Ze65DnXTNf4NUoVyYqDAR+HgAVX7ZSPvj9b1oP/PmPnnbBAl1CnQSfrkxddyTvoEuT0t/2AyocsqI5zCTH7XccoKLrHP2kn7xN6YgMrEKsF6ywC2v3uW1Tum/sHsCGSUJ1XN7oCTr3b4MbJ8ixQEVH6Gd7uMPk2pmgPJUW3d3ac1z1BTM8v9hyjL3vre1yn3f3923/WmNtDbpV99oCFcajok5Ji0oPoEL9KghcDIxMIBAOIRyLqxZlC2jVmeRrIxjxi3SF9T5QoKKAzfUNrjTCiCBQwd4tFcsI+oNSSZhJJ9GoV3B3fkEWr7GJSTFvZlXu7PWryK8tS/IylRkUjwH2AoEKGrXG0pRAoSxMSKr0lFFhpJ/ausm3P1wUezEqCFTw/GRUcBFW6ScFKizVzyZyVD+eCxarBhoolmvYvnM3oqm0ABXZ9XnRWI+GQ7BABaVk6McQHxx0gApKP03vnBZmyu4ZBSp4X2RUkHLLAIjJHQEf6lVEYqoPzqDJVsvbxI4NeC0dkwsvEz9kCSwvr0hgImba6+uSgB8dGVHqbpAAR10SO5trG/jwvfcwmBkUoGLn3r0Yn5yQPmCCITOYliQoK1G9QIWtrLQyUGyTyjxQN7wEAhWszBfdTxMYSXKDkh2tlkhTEagYHh3Bc0ePiNwUq2+trIRWdLKCqC3snJWlZQE3+MZT6kSCfPqjUJqH1caGSWCTTb9+69fSr9/73vckcW6DOV7DFwQKxbxIIlHORf0i2nL+nOjGl4S98c1nnpPr/u3/9bf43d/9PTz73DMIhplw0eoO6w+impR1FuiLxAnZSAw03333fanMIVAxMpKWINgGaFZSQ4AKn1bVtBo+vPrya9g2MYkjR55FOKwVRdWaBmCkOmtQrmyOzz//HJVSDieef76n9BPfty+++EIqfSn9NDw4JDReC1Tw/SBQ8fFHH4mHxY6pHSYgZjV5EOtra8JssECFBLFi5u0Xjwqai+/atauDUXHm1GlhWdCY2wazZMZQ+umhRx+Cn4yKch1nTp/BN5487AAVV67NOkAF+5XXPXz4MCj9FAyH1DZJpLVM8sBMifeSfpLZvA+jgusfhZ8YB/vF1K8hnjJrK0u4cf0ybt36ApVyQUBYMpGGRgaRSsRlnktlJhCPpRENJ+D3kdHAMc35yY9I0qeJ9DDld2iux2mXmvY1vPvmq2jU83js8EOIRtOIR4fQaPH5FrC5sSKSZ+xjGgOPDg0hnYzJnEkK8vLqiiQSaWA8NbULA/FhhIIJNNs+1AnKG3CC3cOpjxsKvj8fvfEarlz7CE8+vQc7p3ZhMLUTrVYC77z7IT755GUcP/EMnnjyMObu3MaZ0+cQCESxb+9BrK2s4caNyzj8jSdw+PAzyGVreP/dd3D8+NNIpEfRQhLnzp7C7PXLmJnegYMPP45KtSmV+rFoGOF4FMFQFK0a8Hf/9a9RL9/EH/3xv0O+OoBSrY3PPz+Han4Fjz+8B+mRMbzx3mlMjA7hwIGDuHDhClZX81iY3xDAggy26Z1jAlSMjI2L6TpNyaukyAO4feMyGvUiZg7uxuDoDgUq/AMYHR0S6Se2686NL7Cxehbf+c4JrG8kUGwMAIG2MCooxcR3uJtREaB3UVuln7g545xJRgLlnoIRBWUF2IxGhbkm0nR+PwhUBMOqxZsjo6JG9oA7V3UDFWQ1pQcHZQ600k86/+m85kg/teqoiGwhgQrK7YVkTef6l4ywIn5J5n/OTfzhPMyqwVJFgYpoJG6kn5RRQbYE50++V9ajgv/m+0c5BsowZHM5WY+sKbOrH9zGQILyY35cvzYnsZEAFUb6iYwKnlc9GmICfvKe6IMQDWtfc3JT42btN6m6N2aOllHBvhuIkxUQRtUCFZGoA1SI9FMxjyTPY4GKth/5XF6ACgKhrNhjwR2ljbjGUrLKm3Rixb+NETqkn/x+LC4uS9u9zA+uJVwz1jfWpZDAMirm79xVoCIcQbFSwNqGAhVk+3EtlqhWNqYKVPDZEqggwG2BCg7oBhMfsqnfmiBzC5Ns7aHWJ9skhTIqmrKWkR0qkl2UFukCKmxBgFxD2LoBmV8Y2NHXg0AF/26ZqZZVIeu+VGmqBOSXARW8dybXmNDySj9Rco2fhVrDDxgVWzYKX5re7vrG/R7/VTLonZfodYUvByp67YD6eFRoKUbPLVPvj63JRI/v9EvA99t7eRK/Wx/Fl/etm19mRGE1rjpBjr5nuV+gwgEY9Iwm/+s0+18bUOHsTzuS8NYxx2XDOI+mX0fZZyp7eJPGtntvyX/YnIF3fHkAF/M9hwHbw6PEW4foBSwYG/K52kpsBR0kba0FIl1glg6nrTfiAMQMOsX4WbSBJB53gJYuoESS5C2tAndZcFsLT50hb7TvGa+4OQqPEoX7qVmP1PyZSWSR2GmyyENlpjSW1OQ+40nxQJD9nOabZC9p2sVjNUlsgAqyAgzzQTT5jR+JPY7X1AJATSbLemyq3JkY596TQADXWel7MYw2ca3x2bQm21xHpMq+A6Sw6X4D2BjGN2MNxjpUZaBigZVsUlNv631AhgIr3dUrQX09GvIcuO4R+JDf0xCZ+whiVpSdFLmisqz39DhkEpxFaDonKNNE+ssk4WXtFSkxfbb8PfuETFzudPh7FoVY/wv2IWML2YcxMU8vkqD2m/UV4bmEDczCGlFFCEh8yvNT4puxotwrwQeeg4AUixtYVEXzOxm7LrtLxh6rR3ifBHSEEaNFilooqAVazljrMtP+wR+SOWq8YMx3OUYsIMT4IkwVClbpsRDUSDKxbfw7n7+acKuKgvYZZa9Urkx8R1ioCn12wkK25vEyXvzSfr2eMnkJVDTqqpZhQRZvPlT2jHwHWBwkwA3BFS/roxeg2Xvi6p4LnEyeYTCxZ6Xw9gFQ0Xvtf/Dpb24P/NnvP23oTHZ514mkaw1y/+0YlRmVWqPn1vd4S+n1VCk4cEUHUNE5RfXqUdcfw7TPQfVNIt0sqF44RM/THVX2C5U9wVoXbURRfH7PPZfV6XWu0cUZVZpsJyDgtK2DUWHmdE9A4t1E3mt09TiNeZ72W97r24BoK0hhkW/3OTqdq9Iv9j4kdtMArxdQUatXjZl2L0aFMiwIVISiEQSpf80ghLEP97is9gj6JIHH1B8ToepRURLpJzFVTaUQTyVFT56yL0wwV0tVZETSKIfFpSVkMoNIDw5JYqNYquDmtSvIri5JJWdmcEi0GAWo2L4DtWYT6bEhpNMZEGwQSqNUPahROCsv7Y8keA1QIQtToyFVpfycbAyePxxkBaoyKrgwUTbCBlyqx62BFnsx4KdESAOVeguT26cRS6eE7rhJoKLdQpQyE5UqGuUqysWCJLIGhgaR3VzD5YsX0Ko3ML1rGtF4AtMzezE8Pi4LaTQW1+QNNc7jcQFMmCyKREKSwLW64baq01aAircCAQ7zI0aplSqWllZUniEYwtr6Ogq5PMbHx1Ryg9IbwqgIIrexiQ/eex+D6YwkmHfu2yssBya5+FzJqOB9sz1M5vO6oiUtZtIqAcE28TNbyctrsEqYxqkMkmTcGX8LAhUMhxYXl/DqK69gbHwcR44dURkvY9Jt6bISNLMwxa96nQQNmEwh84QSUhHzbKwkh/f928xl5dinn3oKe/ftc4AK9g9jq0KpgFu3b0uwxsCTSWUxHV9dE2CE7T2w/wCK+aKYYn//+9/H4ScOAUENqnkegjn8j+CaBG5tNRKfnZ2VQOjT859hdGQMR48eo+cvKtWyMaPXamxhkDB4I1vH75N34/XXfo3xkVGcOHFEDGP59gujQuYZ4+3TViYNPSqqZUo/nZSA1pWTUkyVY/aSBSpOPI+x4WGVb2Elr9m4MUn64Qcf4FsnTjrME5GdabexuLgogIGVfpKKFcM5e/XVV7F//35MT09vYVQIULFtmzDayBxRQKgkjIqALyRAxSdnCFQ8IYnERqOGK9duyjifmFCQ7PTp03jqqafk32RUiGyT0QeWTY3Zj/Ieeykt23eWc04v6SelU7grjWwC5QM12S7kN3B7bha3bt3Cxsaq6O6nMwMYHhkU+SaO1WQijUR8ENFoAgE/q4RC8IdDGB/fhkhkQAr+dDPLjW0T9UIBr7zyC2SGIziw/yBarbAAtxvZZZlM06lBDJNZFB9Ay+jXCt3dF0GzHcbly5/j7t1ZMSqfnp5CmlXJwTBqoJSQpTPzdVMdXB9BjEIFL73012i3lnDo0YcxPjoD+NI4d+ESzp1/E4X8Or73P/wb8ctZ38ghEmYFeBy35+5idW0Z0UQQzzx7BGvLBZz68EO8+OJziMRHUGtG8c5bryGfXcW+md3Yu/8htNoBbGzmEI9FMJCmRGAQ7Rrwi5/9BNXiNfz7P/oBbi1UEUkMYmlpHguzl7F39zi27dqJa3cWMTO9D+ureVy7yj4v4PKVm7h29ab0x749O7B//x4k6CmRzghw7QIVV9BulbHvkT2IJkaxmWVfxDAyMogCgYpKA7euXUQh+zleeOEINrMp5KpRkXHLJDLCMLCMCr5DwlKr1yBABcHnaNwAeJQuLMs84Q/pxonzJD0hKEmnQIVPgAoyADmfF/IlkeYTTWMxKGZSmgbPLWEN8Fo3rl9XI/kxAhUhWc+4kSYbTxh0sr6pprIYXTdIh1dzas450WgYsbAfq6srMi7tnMz3iBu5UqXoABW8Hu+HbbKMCr4FbCvXQtsPwhajvFEuj2QqJQCIbb9W9XGdion007Wrsy6joguo4PcIVPB8nPPIWvNKP3kllYQpqNlPqcinjxSfB701mDivN+uyTpNREfIHRVpB2J/lkoAm9L6iZwZZTt1ABWXVCFRwPZaiCiN9p3/qRtor/WSLAQhUsO18ZnbNZX9xXlvfWEM46gEqbt8VOSwybMjk2chl5d6Z+Le63pKU4JzepI9HUzwq2G5+TxgVBAJMdaTMbR5WsLSVUZapbHSSAzZpZn7HeXJpeVH6zgtUOJWPTqWgMahlosUXkPmenR+Lq18E+4X3rs/bmFMa6aduRgX7S3w2olpEwOIIxkUEM8T4PMDxr31MqTIWRohpfHPoXxio2Lp66BbHRP1bth39E+pfntLu2hX0rda/3zPd7/H/kkBFv52R6KD0/mW/2+tnwH2/QAWv2u9Z9PvcJr5Niw1sYHZcngZ/GbPCA1RYqZEvy0x0JsY7gZ+vA1Rs2WmbCnlvO/phPGYXbAbUlwBNHrBC8wKdx98L+FJgwOzMvX1vY7jOLbPzVJy+6gIqOvMA9i4622MfvWVCS/LfxptS+e9JFZhYr/vZeZ+V9cmUvYLNO0jCXqv9tzAqhBGg8jc2nlWAwMpOmcXS3q15btIsOb9W0ut01vkEbbvkvC2V4BF2ANce4/khFekSF2txFtst8pZGhprf8QIVkmWQhDz3eywyUykePjn1RvB4VHi8PtgyrguWpcBYWaAskygRFofIyBL88OSGTD5DjKiDWvCqlzDPsa1ytOKf2YaoNsh1jGE3Yx5JgBuPCge0oEyxMDaVyaBFZSofRCCBahDc64q0MSMgI6ek7A0jXVyhTxqBGC0QtuuJMDtMv6lvhK6JwpgVvxJ93sLAZL6BShEiBUXipZ5bZJl9ygBtcl/RoCSRMgjYR2wri1gEACPA1LQsEfUb4Y6JxX6MrzQPoubPypYwrBXzsgkYJJ4Qup9UTwcXpHIYCX7ta37/bzxm2j/8sfFiNAWyEgeJKoCybxT4aIi6hwUjJE7huDR/KktHGSk6xtSzhufh99k3BC3cXKPKv1uWqb76LWMgr+wanlvN5nuBeOqV64wlvqNBjgOvr45OX86M0Ve2sJOdZo+Xd8H48cre8wFQ8WXL3oPf/6b1wJ//PhkVJsliJm5NWnt9H5wjjMmeZxGWGd0c27WAdeuvuX2zNVHe0W9fRV+0Y63sdT6vFJPn7I4TmzcAdO9vK6ixNfBwKy48C523E2Vi7hFoyUc92uWgDTqpdj2Q/kOqF0rR62h7Sm8w7lynW5jdObjj8blABQcHzVq52LhGjVwAJTHTIFChjAomYliRXygV5e9F41GRGJ1ALMEEDLW3afiq1FvxUPOrsSYT9Zr0rTpABaWfmOiIpZi40oqDcCCIcqGM5EAMmxtryOUKUsUfjQ9IQqRQLOPm9aviUWGBCpYms+3btu+Q+GV0apsYXNGUiQu2UjsVqKjWK06P2ioPm3ggUMGqWC9QEQqwMlA9Koi8M8FjkzK22pPJZL5jDCCq1Saq9TYmtu9CNJVUoGLtriQ6o9RRJBuiXBVz3kI+j4Ghoa1AhZhp78PQ6OgWoIJ9wOfCfmQ1KPuACSqXxqhBiq0CVlkmHbv8rgUqLIOBgEExX8Do6IgADj4yKqrKqMhtZvHhu+8hnUqLR8WufXsxNjEuCfdgyC+yUxx2IunV0IoZC1RIQOUJ/Kw2Oj8nULG2voZ4jFW3BLCMEXcoJOahC4uLeOXlVwQ8OXL8GLZt2y4Jf2+ynQAaKyeY/GNyisFvuVgSFgATWSEfNa/pTaH+GDaZIuwKHyQptmNqCjt27FAPFQMw8JyUQ7lz+44mk+WdaMs5N9Y3JJlF6TKyZwq5Aq5evorf+73fw0OPPIxmuyxJFwtUsJ9sFbMkDU0SjDIxr7/2hszJx44dx+jooCSrbX+JCZs8s7YEm2xvrdLAq6+8gcmxcRw/fsRhVBCo0IDKBSoYWF688BlKpTxOnnxeEmLsO4dJJNJPwKUvLimj4sQJjA0ro4b/1Y3GLJOkH77/AU4+/zx27VQvDwmc2y2pfqaUE0EHgg9iaMaqFQBeoMIGe1b6yQtU8D4JVAij4pED4lFRqzYFqHj6CWVU/FMDFZZWfm9GBad7d753/mqmUj4rIqtqtr6AhYU72Fhfwvr6EqIDLQwNDiKVTkkikOOWVflMqMciaYyObkMqPYxmy4DF9MJot9AoVbG+ehevvvkLHDy4jzX2kmxOZ+IyR0YjCfh83KjweL+AooEAtfjDqDdZ/VPD9eufY272MkbHU9i9exLpzDBa/iFJGPPHyj/J9qjlR6sRwq0bp/Hay3+DvdNTePSRJ5EamsDpc2dx8/rnWFtdFmmcYyeOY+++hxAOxZHLlbG8tIZytYCN/LKYwS/cWcOFT8/j2y8cRTg+hFwZeOO1lxFAHXv3TGPnzhlsZkuIxRJSIRVPJtBqBdCqtfGLn/8EpewV/If/8EMsb4bQ8nOsVnHx7PvYPpHE/ocPohpghVsMd2YXsTC/go2NPM6fv4DFxXmMjY/iwL692L5tQoAKAlot+FGuVmXJnrt2CT7UcOCxfYgkRrC5yY1QVBgV+VJeGBVzVy+gVPgCL75wVKSfsuUIgrEAMslBDMQ1Cc+Np867dQEqyDyzQIWY69UbMrcSqPAFtfpLgAomaEMEKgKykYsnB6TKixVsFqiwG1IHqGi3ZK7hNTmfjYyO9gQqbIKBc456P5XEo4JzIUFovowEKuIRggCrUvlv1yyuY6yUZHU/E+FkVBCgoKmgA1REaEqt0n4C2hsmiIA1DfVh0DGedjZ+mrAnWMuEfwhXrxCogBolx1ixR7NpTW5b6aduoMJKOligQosJAjqKDVBB8JhgTSKRknPXmgRuXKCCfUIviEK5KN4QQW58KcFGoCKfR6tdR3yARs1cG0JYWlpCPpdTE3BToafMCheo0MQ6wSJleVCWUsAS41HBe9eEAIGKdYQNMMHnON8FVGzm1aOC5t9ajasJGc6tVfobNRtbgAoutg2pCiSgTL1uV8vcVp3aClNvIsqu/xbEUKCihkSSIJyatZL96k1QWZZhJ6NCgQpWhfL8NpljwQregySsrPQTzbQJPnmkn3iP/IzgtMheBZUtw4IMJkWUoZOSdyXUGLwHUOHKl0gUvmWv0itwvr+kvSaSOn8eABVb+7VXr94rsdxf4rbf1uhrABV9GRh9xoA82PsYH5Kp6ncuJ1DQddf8v37a9Z0eZt1OL3jP/5XGt0fyyF7LsAP6bmH7eVQ4jITOZ2Ir/72f/ksDFaITb42VjdmuJgp1TpM0tSdvb5OWqodvgEfuV805eg0FF0fxxIVecETiK+NX4Vyu/3jyghROgtLIB7Fi3mVjeDSnvDGpkdNhItcCAOIxIJ4M7tPplquW/KcBra0fgO2bbpDL/bcCFtbgWkaxSbJzDVIZIXNRwyBgwl0llLSPtfLdTfASjOFnKj1lq+qZh9A518umcAAPtddz/PwcpqApVJSkNK/HO7ReA1wnTSGh9IXzvrFftfxIZKOsp4K5hgMYGblhvWftV636p6+iX5LoEiMI+YSAQlP2nIyZCMwz5yDMADGt1j6xptXqbanJfbuWKwBj5bL0WTFm5lqrxtHq36USVMrkFUaLYXCwjdw3ULZROBvmGlqkrz4gLERknxOkobSxFDgGjUeESCqZHIAwJ1UqysYTjsSwtLErvyVgmL5PPIcwLn3q28h2kr35V//ZZR/88Mc1AWbEc8ICIQbEEhaHYdLKvYkxOOML9QyjNJK02wBVChhpHEFwxu5VFcDQfpS5wBRVKFBBNg5BD/UBsSx/FmbIHq/b49WcqdEiWKR7KgV8XE8W77zYAYR2TqM6O3uYRN6VQcYw22XemQdARY/Oe/DRb3YP/PkPnzLvpRs+CMroJMG7wwrJKncF+jyGyGPvEMS7oXF7SyeCntUInMi90ak9rQfh7r3R6AYsPEn37sdky2h1TvLCmc5EZWZ4Z5LQg7xG1Fbj0bPxMdUWbpVHZ79q3NkFBjj/Nqted1v7BLjuM+rceHVUXthnYqKpts94bXja4J7eu5lzw2S3e7rNtJXOyUncelQwsa/ST9ZMW+VrLEhBACM5NolkJk2MXxJEsrnlxpdNC1IeI6ZABZOgNZdRQaAikUqKmTZHCM8bDYZRzBYQjYSwvr4ii+T45CSCobAHqLiCTS9QQemndhvDI2NyvuHJCUGkLVDBAEsomqQ41lyggt+xSX0GENT2JlDBHzIqMjQQFUZFG5VaUYIEq6ctshuGPdANVNQabYxv34VIIinJYgIVDBBjlCISoKKCfDYriZHU6DCyG+vKqGg0sGvXbgxQ+mnvPmSGRyTxzQS3ZVSwKpbt4DOJRMOSQGJQZJM7trJTg4Oa/E4XxbYCFdUaFheW5L7JPGBijQl3GvLaSmEm3IIBPwqbefGoSCVT2LN3rwAVBI2Y6KGxV5JV235Kg9BoVgMI1ZjUyh5rLiUJiBiZIHUJnGZvzmJtfVWSgExgW8CIlR4MGhfnF/Dyr14WRsWxE8dEe54JXzs2eT/1Bk1ZWZHRRDKZkr5j0EKd89XlZWzSU6JYQjqVMgkRa/St1QqsoN22bVLosmQv0AeDfcky5EqtjLt374p2uWpw+lDM55HLF0QeJJfNYXNjExtrm1hbWcXv/u7vYtfuXQiEWlqhw6pa0/d8LsIuoezLQALDw8MSKL722huSdD558iQmJ0fNRkC0gKRKRiplODP7lOXQqLXwCqWfxidw/PhRhCj91CZI5AIVOk9oddOFC5+hWMjhW9866ciFORUiDMzbLZV+unVLpJ1E+ousCPpeGKo2gYoP3v8ALzx/UmSctMJIKbaUfTn18cfiE2GBCgZwXqDCeldIJY4x07ZAhdwnGRW3bytQ8fABqXiuVho4c/r0VwcqpJL4qzEqtmwOrema9bhw5mkyDtxqGtlMSKWOMZsn3b9NE+8gOP3SdyGfW8fy0l0szt/C6toSarUyUqkYMoNJ+Y/GtemBEYyP78DIyATiAyn4AiEBwJeWl7GysIJWs4y1jTnxwRgbm8TI8LDIiTGxC0SlfwL+mMyzBC2UHcEqaratCV+bwM91XLp0Dul0FHv37UciPYZwJKabWbklHTciEVYLYX35Kt5/+xeoFjdw8MBB7JyZxicXzmL+9jx27ZwW09s7Cwv45nNHsX/fwygWK9hYL8AfauPzy2fx7W+/gMW7K5i7PodvPvOEABULqwW89evXMRAL4OCBvajX2iiU6jiw/2HEYurR0Gr7Rfrplz//KXLrn+NP/uOP0fJPYmWjjLW1FZw//S5mpkfw6BOPohmMIJeL4NrVOWQ381hZWsW5c5+iViti9+4d2Ltnj7DuUqmM+PnQspAya0QaZ69+jmCgiX2P7FUQJc8KtQjGxkeQK1LKrYnZy5+hWr6KF188irX1ODZLUYTjQQymB8UDQebSqrLYuOHiuCUYoUCF9i0BQ87R2WxW6jxYZUgAOR6NiqSd16OC0mn8HYEKK/1kNzuco3leyhtZoGJ8YgLDI6Pw+QlA87+QVs4ZurskCpq6NrGdnFPJiOOPeFTEVOKPc6gFbQWoaDVRLOdFa5lABc8ZicQcM23LgmNfDmYyTsUej2MynUAF1yPOmwroKtjK5LNIHPjDuH51VtZwL1DRbOsm21bZsz+l0p5JbalOU6BWmBqUbJINayejgkAFARXO/SJJVSMgbzwqyCYho4VARamovgoOUEEz7SLq9TISqbhW8wfCAlSIVJeRfrIbWhsbCwPRABV23Z+fX5R5mpJObJ9dZzlONrObsm5z3eMlXjfjAAAgAElEQVRzvHvrjsOoKFaLIFDB++d37bOnjjWlRNi3PEeZUpiGURENR7Wi0Uo/ca41CR7LppC32zBEOYZs1aBtF2NYjkMCFSL9ZMy0yX5lsYCT+DEbb/l3W41JrUcFgQq2m/3C2MIyFu09WKCCsoacZ8jYZL8RlKG0BOODNTEuJ1ChDCE+AypLsGKU44kxHGOIcO0eQIVJiNgp+6sBFfe5t7tHJWTvM91HovvLmtIvCX4/yXQdkV92pR6/75N67puY73OJfpc2RRg9v9Xr0vc6vt/d9e2/vl+4v5vowSxwxmLPM5kS254Fb7076us8OcebwT77HjJG3uZt9V002+d7ABXdt9fxyLpxGKlau8ed9AB8tNxlq/RTr9yCjPBu42/LqrUsAgMcdEi4mKS1J+Rz/npPoKKj87r296bPJM70POdOAMA9QS+wgr/1pEdcrw3ThZYNId1mJLsFVHYq2r1yUwYic1GWDhks+4poAr+HTJVlhkiSV5PqbpuVkaEgtSZVtXxd70+6wNRMKhbkk6SuSkMxPqI3FCWTVELHqZi34Du9DiQhzL27MbEOhbWYziTdrQQVz69yTWpcrWbLWpym5t2utqF7zyrho8VbCpLzd5YlKB4VbSBC+Uvj90hgh/+zHgfSNjIfK/Rs1LmWfSSFE7WaFMCx6I9t5noofh1GxUET+gqsWMBIGRpM/mvbLDuB98JiUYL4jHlYYKLrq0p1c01XeSplqbCvKcvNIiOCKSIfZEaVSFTRw6JclvYJi9PkZpgi1H17SPaolBW1UlJaj0tWql+YnQzqyKplvMI1nc+ATFJhdVQ1ntMCHgVW9N/AX/4nVw5KgQr1WKS/px1jEruQ5RBQJg2BCgt4WLlJ9p/GN940pUrriWKA7VeRsdJ9PJkm3u/o1GNzn945ymMGT3aFGUu8j2qNEln0TlQAxI41yW3V6xLjCbvHxGL2XoQhYkAvy4CyoJk3jlN5Lu0zDXF8DxgVXyOCefCVf+U98Oc/fNJd6rxAQ0+gwi6o3Ql7u1zqZNn5szW0sZOgLtCyLMlX3AXXrrJ6Jm/AYRdJoWlt+en+zD331mMVzfVuWOwEoC3xnEsy9ZzQOFN5gQqVxnABDKWJWZS/WyrKbYOe37nCV61+6b4Jg/Dbj+29dAc6zj3KpNxV9WXZMLanpVHu/Wt/O5GbS1ET0yVSCHXDqoyKhhjdsvpTGBXyn2FUlCuGYVFGZmpaqn6pW12ulB02hfS/3yeVe23R+idQUUapWMLmxoaYaVP6aSCZ5komFfGRYBCFbFYqmjc216VKdmhoWBaL6EAC5VIF169+gezyIgaHh0S/mxRYxkmZoWGMjI0hPTIiLBECFAQgbEAh12eC2wRGdjGxyX0GADw/+9cCFZSPkurBWhmNes0DVGgliVZEcEOvhlHlahO1Jtkd0whLe+nHMS9GoJQAabAyl32YyyGX28TI2Ag21tZw6eIlQfaZHKQHwsyevciMjfKkiA8wQFHAgZWqClQw0KDh91CHcbNUGRjDqLox/7YLpAQ69RoWFhckMKBROJNNNHWdGBtBuVaUBJsYuPl9AlS8/867wqigRNKufaoDn8/nRHaKlY8cWryOJiiCWxgVkjihlJG5NqV6bl6/iaWlRaSTKQl4yBpgskLkSuDD0sICXnnpZfEgOHGSRs47zfhS6rEYajHAbdYkwSJsDVZO+ICN9XUJsprVqshLMUFH0IVVtZJgYrAVDIgUytS27ZoobLdFZ53eCcl0QgKjhYV5CbjYxwx0yI7ge8BAj9dYWlzGytIK1lfXBajYOb0T0QTBtLgkCwl68f0hayaXz8Lna0o7x8fUn+Htt99Do9HGkSNHsGPHpATTTAzy/AR9lNKtiXGehwUeL730MqYmt+HY0aOS5CFAxoSWBtBMWDNQDqDebOLC+fMoFvJ44YVvSWLJmonpHE0xoTYuX7mC23NzOEGgYoiG3lr90zZVKlevXsH7772PF771ggAVStfWWY6J1o8//lieEQEJJuOs1iwZFfv27xPpJ6XoQpKnPH569zS2b9subWWb7ty+jWKpgMcee1iqnUX66ZNP8CTNtKNhtNoNXLs2i2Q6hYlxlX6i5NRTTz0p0k/WxUgCYTNx2hn8Xht9iy97Z253hRBXB888aT19tEqPfSeVywTzWyK4osf72igVCpJwXV5awPz8LWSzKwgEm0gPDmCc89PwGBKJNDKDw0ilB4WBtrSygma1iUwmhUSKuvkm4G6r4W8wnEA4lIEP3JyYINnHzanSw1tNDYKlKgttkU767PynnFLx6KN7kBnMIBKJi9xSq01zOpoKB9Cq+7G2eg3XLn+E3OYKshtrOPLcN9BEFflCGTt2zAgQ8st/eEne0RPHj2NqajuKBd3UvvHOP+C3vntCQL8gwti+bReisSFcvHQDZz89hYGBkCRiN9bzmJk5gJnd+zE4OCzjq9nyo1lt4e//7/+CwsZl/Mc//TEQnkA2V8THH7+Hm9cv4cD+3Xji6cPwh+OYX/Tj2jUCFTlcu3oNN65fxeBgEgcO0F9jB2LCuEsgmcqIt0e5UkO72cLc9QsIBGo4+PhDaPno0cMkawRjwqjIoVpr4erFs2g3ZvHtbx/F8koMm6UIQvEABlMZxGJxBQaqdfNet+RPAvBcRyNRAkik4DdRprdDdhMtX0M2gZL4jsXUD4iG2gE/BhIxBIL0sKmhkC0LOMxXkvRxji0m5zkHrK+tSyL4xo3rMi/Re0OMEgMBhLlhN0AF3yuVh6BsYRH1WlU2f5Lg90Eq9uNxesqsGy8JNXgkiMv3tVDOC6gQp+RTuSb3QzCbQGQ4GpbnzDVxUMYQDSFrut40GsiSUZFQ1pDKDtRljiCjguCH3xcSM23OZ2yzelSQeaWmnJQYYCKA/cn2rq9vIBjyyfzFRrLtXLvFw4Agqdks0z+DSQkCKMlESsDmKoEKXwvxWEz+Le2uUK6yqL4KTIhz/DcJVBTQaDJRPyBrN9u5srKqsoEe6ScBqX1aMSf9Hg6b5HpI1vo7dxelrxNJtpMMJZWkaNRbYkLP+ZxjkqAAAVnKGhG4IDiUK+SN9NOA+HJx+hAAr9UU0IVJAFY7CgsnHpP+k8pPAwhxrFhgQZJFBky1wIEFKWzsKBtyox9O2TbO16k0GTYBAVvFN9tQrlSWQqtPGRPyuowZeC4CFWwPz0dgjGPSJpk4/drYSs20/QJUkN1KZpGAPZGIFBPUReqQgBJZegQr9E+Of44nJofC9UxfRkV3rP8AqOi3Mf066e5/QaCi522YJOj97L3/yYAKmzLq3gbfg1HRq50i8Sh1vT22rv8MQIXNGsvV3ev9fw9UdIIOW3IJqoHZkUC/b6CiB9hhb1MjY7M79wzrjj21Zv3dn14eFfcae1Z6ysTGmi9wT9IPqJAn8RXGqbDdTMzpsh9UaJXFCyI5JQl+ry/nVq18Xsuex9RfeqSQbFtciSat7O994zbBy/mf8YDI57A4oo8qBPdn9hh5D6Syv6aSTpRTkjWWjGFNXPNRcY/Hc/I4rkcsZOM+WEyUjdmxxr2MJ5TVoSwNkweyJs9iMm7P6o5/x3tb1BA02a/H6bNTAIEsFWt0bfwGDZAvnhxS5V/TXYHZW4mHhAEE5ETGaN0WtbIfVIZJ26V9bAp9zXuqey31VpA9K3MLBES4LoYj0mfWQ4LnEWBEEuhqYq4giLbJ8fnweGHYwgJe2bI/GDPze9wncx0nACG91WoLCEH5KbaJoI6AN/TpCAVECYPrO2/DMlMcU+2myiox9uCz+8lfxZ0B9f0fUWa7KbkBMlF4DWm7iVO4D5e9q/ie6kAkUGCT/to474zKe22IiTiLuhQ48sl5GWNqHMf4VwEOLUbxMht0f6vPxY4TRdukbQawEDkwAybwKH7O9499xrjHgl0CzjEvQi+TJr0ItXiT44bfF4k3Gcdq8q1jQZU/mDCycnAPGBX3s/A/OPY3ogf+7AdPeogQ3akbnRCdH0lY24oHAy44iW1Diew+3hPmuPl4/a4kpr2ggLmUNxjakszvWuSdtm2Jlb2SRt5fumkpR4dOZh8z8RtafQfrQaZUzwrsNsp8bJNURtbJLPDeAaD37jIw5F9Oh9gT9lnl+wEZHSCDuZqNKLpHn0xyvYLePqwQ96Hrs9IGK6igD0/WAqlal6puRYiZAOCmVhkVClZ0MyqGp/fL5lINhKtOJR8nby4GrHpsN7WyvFYti84/K0YpZj2QZHIug0AwjFKhiHDAj+z6Gmq1CsrVCsYnJpFMJKWSMJZIoFyu4vrlS8guKVCRGRoS81RWDQyOjGJsfALJIRqqms2vP+hoaAqroq2SVnZB0sS+JoBEs9tQIcmkoISLNYRihTQDEt67t4pQgiZTkSJyE9Um6k0oUBGj1BI9KhaERBhhhUKtinqF0k8F5HObGB4exPrqKi59/oUsZLt2TEtyY2ZmNzLjE3IfMSa/awRQYBD7mjwXJpgIVPD5cHG0Y5CJNbJJ+BkTuzYoET3wpgIVlMGIRRLI5wsi8TQxPoJSpSDVsAwG6BVSyObxwdvviLQHq7On9x8U1kqhkBfZKQEqxKOi7nhSOHJYrIYxla1kE1D6htrbnG3m5uYwf+cOhlIZGcMtlnQaWSEu3ivzS3j1Vy9jfHQUx58/gR27dkqltOhzG1osx5ZN5jNw0zbURVaC7yUraDmm2f8Ld+elMjxlNNppwExWCNkJTHZJBXIoJAHT8MiQAGsE0mg4ZquKCTiQMUBKJqum5+8u4M6t21icX8IPf/AD7N2/HwPpqDwfBuUEKhq1hvT/xuYaGk01SKWmOgOtjz48DTp3P/vMM9i+Y0LGHpO6nEMZmDkyTWR4VKoyTf/qV6+KmfaxI8ekXRzLHBf8YVU9+4aBJPvp/LnzKBOoePEFx0xbAyH2tybbr1y9gluzc8qoMNJPUqltgiYCGe+/9x5eeEGBCitRwj855j766CMBKvbs2WPkx1Qn9jXjUbFj504nSOb9nPr4FKZ37xIpLwuczN+9K+bljz36qFTvVioKVBw+/DhiMd5jHdeuz4lsjfWoIFDx9NNPC5sjYKZAK8d2r0X6fpJZ3YC3Pa935eCbr8rw9oeggVZD1SqU4ilgbW0es3NXcPvWFQRQwsjIsBheDw4NIxyhrFNakuFhMWduID6QkPFLj4IrV67iqaeeRjyRQDSWhM/PgJ4ccz9aPtK3uUHkNWkCqHqvymoKCVvrk08+Qqu2iscOPSrASDicQAtMPkfRbgfRrtexMH8ZZ868iXJpE0u37uLhh/bjyaceFuA4PpBG2xfCe++fwvLKkhh/v/CtExgb3YWNXA5//8uf4ujRp7G8sozDh57CQCxDFXt8/NFZXJ+9glCILLk89u99BKMj2zG1nYB2RvyICFRQ+omMio2Vz/Anf/IH2Cz4ZW64desGisWsgLhPPPkEEslBXLlRxs25eayvbojZOv2LZnbvwP59MxgfJ+OO728CyXQG9XoLpbKCmHPXziEYquHRJw+h2ogIUOH3hTEyOoRCOSdsj0vnTiHgu4MXXziiQEU5jFAsiAxlCaNxnUurdVQrVUlG8x0JRixrLKrrT6OFUqUqQErDR/+gsCTEOedafwNupuMDEZkXK+UmCjkyKhSooJSeJNoJVDSbMo8RDLx58wYmJ7cJE8smzMnQoMQT50qCMayQq7VqAowQTFegQlkLNJKOGkYFWSeUrOP1OO9z5S+UC5IwTsQSImUWicaEFUmggow9gqFlekZlMuJfwXHmABW5nLyXTC5zPrJ6zdxkE2Qko+ImgYq6sg9jAzRubMg8KgwL+ncY0IXJeo55X4hsOa1IS7DvDFAhm3XxJNLjuHetVipIDBAkIVBRVoNs44Ug7MkKiymKklhXbw76UNFIvGyAirj0NX0rBBgyZto28c68DxltUvFvgAprqM05/PadRbkfSkiFgwHU6RvS8qPd8CGfz0pSnv3DufLOnduSSCCAUyoXUCjSaD0msRG1pjmTMKFPQLBUpSyXxiICbsXVBF0ABOtRwfVPGGxtTWSYSkcrH2jXDzvns/DDzmmrayuSNOD6zXGHpiDiJsljdJ7tWmEqXOlRwZWDfUngh/dNoILrTS+ggoAPtRlXPdJP1quKsoG1sjIqCGqp9JNKX4n0E820yaCpE4SiPJf6YjBBYJlJnPe8c/RXmtv7MSTud2fXN7n4dUCBPhf/J7vGP2Wb+rS1D67Rt5DeJgO/cr9/HaDiS07e0S2dFfBbv9k3W9vzIr2T/18PqLifpycJ+a7KeC24MHs952T/PUCFs3vsvVXvarD2RW9/EUnsGpBA3l/ZSmlFtHd/7gyv/lnzLUNNBRa0Md74TBvtlQAyt+EBK7ouf8+B1AtoUFkkc2HTH73GhG10z9+ZZymxvWUrOEGo+kkKQ84YSVvgoLs93i4TTwEXFTJd4T4wAac7Cky1Yrz3j4ICvL70qFlfrBl093cYi7GNUlRhqv8VoFDZIi30Y2yr92ajassa5flE8ocSP2IHon2sRRraRlt5bwEbW9RGIKejjw0wwO/omqr7ItlPmnyRSlMZGSpZc9uyfktOQ1gIWiigSgKaR5PkNwsWrBwQWQYswgiyOIim221Zw6zMkxITDFAnzH0DjJi8iWUAiHyT349ymfKpTPS3RflBAQD1dWBxHuNLMjL4pzxHA1bwvrSQQfM7NkHIdpIRzGIOiY+MLwT3ryqZZKSiBEDQHIm8zfIs2xrHCetCizmUGauymFJIwedifFb4PTJL/stfslBIf374hypLTUBEk/u6m+L4cMaF2e9LMYYwiBW8cuMb70jj6DaFcSZO0jYrq0LHqhcQUqNxO375AHUeUmjTpWsoECTfN/JSBEQ6ACmZvtQfwzKLrWeYWLbasUXFAgN6sPhEZa200ESfjTJFLIghz/GBR8U95+AHv/wN7IE/++ETDqptk+n6Itqb6Ywqqa/nBgVeYKP38fqp68vQeY0+QEWXlp23BbZZnRsN51PPEzBgiK10dX5jE/ZGY9Kgsc6E5AUqHFTdVjtIBLflGlpJ0LkR0oWuu11eQKL3eXoNoX6bKlXT7B31OxUVXSd0Chg8i699Rt1AktDinHoFcyJbTNJhpm2knxoqZyFAhVQnVvRPGgU7DIsyth14zNHl52Jkq/nsgtwNVFgzbSasLFARDEXEKyEaCmBteVmS4aFISHwnpFqz0URsYEAqOm9cvozNpQUHqOAul5WGw6NjAlTE0wQYrEyGLpxcEITGCE00dQAVXIRFc5wBQEkT3YEwhoeGDdLNpEcJzSY9Krg5d8ENfZZagc2FvlQjGOIXM+0wkz5ipr0gDJEwzbRZ8Vqti09HoZBDJpUQKYTeQMWksE4oJ0QNcl5rYED9BpiY4UafCSwLVHDRVwaDASoMA8QuxMJqaFQFqGD1OoEK3o8AFRMjKJXzshh7gYr3334HmXQGe/buw/T+hzA6Ni5JFpF+SlI3n3TZqlZyGMBHgRFWZmjfEzSgpAZ1M1ktSxPiO7duYXRwSL7fNMGFrYpfW1zGay+/grGRURw/cRw7pne5jAqzkNsKBn7HmkUzMbXC6m7qiBtWgPi7NRuit7+0uCQBLlkSDO7oyyB6oax0YFWnaJP7EDOJLa1e0api3jMDM1YZ57M5LC0tY/bGLG5cu4kf//jHePSxRxGK+SRwkyCXkk/GP4IJy2azJgarTPox2Xbm9KeIRgfw7LPPYmQ0I9WslBpj9UWn8TUrh6vwE6h4WYGK40eOK1DRaqBSLepej8kumZYDqLda+EyAihy+9cILHYwKjgUHqLhyBXOzs3j++HGMDo9KoGSBCvbv5cuX8d577+Hb3/62sCMsUMFzMEn14YcfSrU3gQqOQQ26gNdfe03MtOn/waBTrtlq4bQAFdNiwM0+tR4V+UIOhx5/TGSrqhX1qDh0+HHRtGfy/roHqOB16Y3xjWeeEZAkbEzPLBj3lRJWX2Fd7z9Hm+XVLCFCt/asrX6EBaQiI0mZVmQblbCxsYRrlz5AKBLE5OR2AVgJHnAMEPz94vKnMh8cOXIcE2O7UC628P67p6RPDj11ENFECOFwEs0GK5W1+oZJVAbgZD1wTub8xsSopZ7XayVcOPeeSOg98uijGB2bRDyeUUZF249Cdg1nzryNK9fOIewPYWJ4O1ZWFjEzsw0z+7ZjkAbrdT/Onb+IiYkpnD13XuaG508eFU+bt95+C1NTU/I+75mZwY6du0Dlv/fe/RiLy3clCXrw4AFM79yH1ZW8MCo4l3Fr0GgSKg3h5f/2M9y++QH+1//lB/jo9AUsLq1i98y0jC+yvQ49ru0+/dkyFpbWsLS4KuMoFgvjoYP7sGvnNmGpcJ4kUBEbYGK4IUAFy8FvXD2LWKyFx596AqVqCMUS/WjC6lFRzqJWa+HSp6cQDizg5MlvYmVVgYrwQBCDqTSiYTIigqhVCbJznqPkUBXBiEpABUNMpHJOZmVaA9lcAbWmGipaoMImtxWo4PEhlEsN5LM00+a8DqHpM0lN9hyvQSYY+4Dv57bt2x2gQuYkyhxUVf+Xm03OgdUGJRkLaLD6sNlQBoffh1QygUg0KJ4Xg4NDUlHGuZryRxxD+XJBK/8pUVRWj4pSpYJNMgLIqKDET7kqJuXWaFu8Osio8AAVtqpMNsm+tgAVQBCzN+7IhpXtIVBBqQBuDruBChpg09fBR0ZFN1Bh9Ji9QAX3l4wFBuJkG9EbqwxOkrwX/scfAj1cz5lcJ1NQGRU+AX7pOUUmBBMIzJNsbGwKuBjlsZbqz72qvz9QMXd7XpIvHIvREMcIWTwEj8jayAlQQSkjjpvbd27LPXPtIXhOaQZWIaZTgybhrgAj59BitSDzJZMR3UCFTahoQYnOrdaMm0iOF6iwiRaJC2y4126jG6igX41MVZJ80cnMAhw2AeUCFVEBpqjhTCCFi05/oCKI1bVVZc9Eddzzz9XVVVRLNNMm+EKAgvJe+ifPTblGYQ/V6M3zAKjoXK7uJ3UtT/IrrHbdm4r7+0qvK/TDLszgus92/XMAFffqq/7J2l491St5LSmsr8GouJ+nZ4EK2yYtHPT83AdQ4XyrF/DQlbzufQ09w1cBKmTPaxUVpJP6PG/rg9Dd6T18PpyYrGfNYCcbRrIAFlDoI1/dj1rQG6gw7b9HvaKTOPf0bzdgYduk7DY3U2G17Vm2Zfda7BKb+HZjV/fkig3KJN8p6e35t5XQsmbeFgzpNcYl5rBV6iI9yeQ2JW5daR/v92QPbgyPpaCGfkyyZ1SpRzUwNgoWIpHkeibZNcgyEOh7KVXnxteJ51XQi3lkZVbLnZsH2zaAfsd92MQJ959ihKx7FE1Su2A9E+b8sQwIlUM01fhGEor7XMoQ85vKRtCYgffEZLaCPZprstJX3HdaDw8XuNAEuRq0k0VqKvW5RxVQyqfseil6VPY9Yw7GGbJecy8gZue6hxfwwRSi2r4TMEc2xTwfZVBVrle+wyp/ggEGKDB0A5E1FY8wY97Ovuc+mTE3JalEucIYqrOoh3Erny/34FTZ0OenfpL/x19of/Ln9/+nmjAoqFTARpCxyz/VjyOo7RJZMfWLYJ+S1dE5/bizj4lcVP7JDH2XHWHkx+r6bBQ8agnAo94pzhcM4GBYPR7pJ16pwn41pubsMws0iMeGXxkUXlBIPDSkxlqBWJsbk3fUFIMow4LPhUoelN1i8RLlh02q9QFQcX8ByYOj//X3wJ/94AnTSH2B7aLVG6iwC6rXQ8KgiSbM6Ezkyxnd5L7JhLvsgnsAFbbr7HfMv3VB8SCZNujYEumaD7Yk5O2KZFPwFmAwx9tsfUfAZUMCRbDdH3sN91x24dIUvy48+mP7wZ54a2h+v0kzu53sBivcypCt19Crd39unn335yIVpbOfmQMtGcDR+eQi5Eo/MSGuYAWTF8VSyQAV9KgoOXJQ0489JQsLEwMVSj+ZRd9O/luBCur8ZwVciCeTSKYHEQpH1Vw6Esbq0iJyuax4IIxPbpNFp95sSWUxK1uvX/lCgQom+4aHpHKP56IsEYGKWCojG12l2RGE0EoML1ChtD9l6UhiQuihmoDlD4EK6vYzqazVmWo+yuQTf5jAtoltfVW0WqJUbaCFgAAVoUhUgIrsOoEBBSrq9JOgGSn7s5hHOjlwD6BiGwIh9VagzJEAFYk4mo26ajw70k+qg2mBClZiqPGWVj3aKkwCFfVWTTTx/QghHIyhUCwKUDE5MYpSJS+LpQUq8htZvP/OOxgaHMK+/Qexc+8BASqYEAtHtPrRelSo8ZNWntqEtmVXsAKYbRWmANpaNT07izFhvlBeQ8ne8kwArC2uKFAxOopjx49h5/S0mBPzGXsZFVrloLJSVrZofn5egxwT+Eq1i2inE3wK4tOzZzG/MI/tNNLePoVqpayVLgZ7VQBLK4nU2DMtj5fPndcOx8JSuby5kcPs9Rv47PxF/OEf/iEOHT6EUFyrQiXUbbYk8WXZB4zfs5tZrCyvSSD74QeUxkmJGXE8wcRaW5KRlEIR42tDQybbhIEi6U7/+I+/kjYfe+6YGrW1qEtfUKqqTwMlC1ScP3cO5bzLqJDElnNOVgq3BYigsTkZFQSFuoEKelgIUPGd72B3F1DBd51ABVkO+/bvl3ef1dxswxuvv46DBw5IH1uzMV771EcfYXr37i1AhWVU+EAaeUs8Kh4/9JgkANtoKKMikcDE5KSM51OnTuGZb3xDDIYjEmwrSGYD/n6rdK9NZb9j+1XrcpyKGbX5rxOogEjcMbHtl2CZMkElbG6uIru5imiojJHRQQzSe8YfQKFYxcrKGs6ePYcLFz6S5Plz3zyGocEx7NyxB75WWFgoI5Mp7DkwjXA4g1AogybNs9tkYGgFEROWluZt2y008HoVzXoe586dwcrqooBHY6MTSCUHcffOAj744E0sLs+KHNGTjz2DA/sO4caNG/L5c0cfwsTkGHQ/LI0AACAASURBVNp14IsvruPgQ4fQ9EXw8quvIxyp4be+exKxSBLZzTLu3L6L+cU7OH7iWZTLDbz7zmnkihsYHx/Fc88dwdpyDmNjO+W6rDzjDNlo+JGIJvDqP/4cly+8gT/90x/h9TffRSSaxMOPHsby8ipu3pjFww/txfbtUzhzaRXzi2u4euUarl65ionxUWFTTIwPI5MekpV5YCCJSIxV/00USzWZc29c+QSpZBCPPvk48iVq91LrPyIG9rniJmq1Nj7/9GNEQ0s4ceIZASqylSiiBCoymigNUGuXjApuqJotSYqv5W/h4oXP0WwHcejQUxgcmkC12kYuW0KlrkaKZG1xDvECFexrzs3lUh3ZjYJh91mgoiHSQxynXqCC75FlVHA+CXHM13TDSTYYjb2rdRYQdAIVlDNIpxIIhQPCYKTslmw2Gy3DqICYTZP9MRBLoFquSMUeixA2sllEYjQ+bHkYFfRKUkYFq8I2s1lhWhAcsyxFrczj3EnWTgBzN+46usexeFSAR5dRERHT73qlJvdEoMIfVrNJPjuCJ7wHqeYTENnDqGjQzLkmHiKyuWtUZYPK5DeBCvYN5yTOF+JRIfMy5wqfSCoR4CVQIUb29bYAFaoxTBNwjQ04l7X8mlCwoLV9lpxvZufm5ZqUQYxHw6qPTVJZKyDSTzyWfcP+un37lrKdwiGUykXUquzrKFLJjF4LAQHYCeaT2ch5hu3ndcXfQbyfVDuZ87StKLQFF/I7w0rknOad7/lvF6hoYWW1k1ERaAdMDssw7kxywYIVPHc3UMECJ5EPk0pFd813pJ9i+vx5LQtUKKMkKsbutXLZxGc08lQDdmumTQatxBIPgIoey9P9pK7t3qjfKtfn8/u8RK/DHwAVnX37zwZU2Mvah9JRUt/9S5d14G3tvYCHvsCXvU7XYLgXUCHncoIpc1XRmuszbu8BVHzpCO/a/zvHd7VbwZ0eo7cvs8CVb3JzLTYx7enfHi9JN1jRD6jQ7aW2S7askpDWuM/mJxQwtiwAb/s9YIVhZnT/1ib2LUvB3se9gAobS9sqd/5b2B2G3bDleVAGp67JWFvoR8a6gCJGqslel2uI7MGNwbP9vawt4mdkKuFFMpPxjPpJCNDeBXJIitib4jFDywIZwsxvsVCNfnHat5TlYdwhChOmLYzXbVzBQgc1YA4a1j2ZkKyw1zaT1SDeGFpBZnw1NIYQmaqAXxLeVFiQz5q23cqcsAbTGofo90SiMugTXzPGCYxzxCPKFORxvQ9HoirPJECEwUaMjwX7nfkJHUvq5UFggAVOUfoqEKTgPYuhu5sjYkzEGJjPSgpzjLyzSISTIcO8T6UqRRf8d71GIMV6npApoIUMKgvcwl/+J9dM+wd/UHaen+ThBGhSEEWkwSjZJJ4kPEdAnpGVF+Z9CIOh672WwkMDNDk5HhBAUJ8SSl7LMcIUNb4bxvRdz6n/70yf4m+hJu/sH/2cstNaICTeXuwHgkqUbWo0BcjQog9lf4g3C2MkIwXFe+GPMoD0uQhgEtDCSCpuWGBJWvMAqPjS6f3BAb9hPeACFfZVthTEXslsU2FvoPvOBbp7EnC/rwtKFxBg+qmn9JNjTGpgf2+fWrqhpVz1BSochR39tlcLUcy6NSjQjZv11pD0pzm+46Km0sPS4TvBCrsIq0acPbMFKngeL1hhz2uBIXe6u9+hY9U0PU9Ob9VTFdXp79HvWorcd9XTaIqNz9pR0WI1sOGKWPqjoTmqR4UFKmqGUVHuYlQoWHHg6SOyGdfKfk3OejfKrJJjdSsnbko/MTlMQ+JKrSYeFKnBIQUqcnmpTFxeuCtJ/NHxcQwPj8ozoJY7pZ+YKLlhgYqRIZFQIVDBoGDH9G6kWPmZoFEtN79qbMUFjgueJoAVsHAYFUwRGKCCn7OKkc8/HIpKotzqRFJqqdmoOZWoNmgxw0MT3QE/yrUWGm0fpqZmECBQUSpiY21eEpc0OK2zKpd6/iLvsYLBdNIDVLQxTTPtWBwze2aQHptUoIIVGw2VdmLShYCJ9ajwMipkZBqtT7IqeD9MltnnIcltNCVRT4mKeDQpCSsyBLZtG0exnBNmQaValmFC6ad333oLQ5khPPzII5jctUekuOhRQeknSkAwACJIolUWnUCFlasgUMG/M4SgRwarhO/cvoPx4WEFBTxABRfujZU1vP6rVwQoeu7YEWyf2oHhkWH1NaBmpxlfFqhgIscyLKiXzx8mwKhRTnPWNo3Pg5RBSeD23C28/us35fm/+K0XNMFO4zCjIa9Uasq4qKRSkhWemYz0JR8yGRUE2ajbTq38c2fP4/vf/z6e/sbTCEa1AoRBruiqmgBaE+gMbhooFgjmVfH6628hHIrhO9/5NqJxPqu6VtyGVRdUEnQMhHzUAq9Idcrf//0vsWPbFI4fPa56pK06stkNqVL3+TXQ5txUqddw4fxnKOVzeOHFF9XDwyS3hAZMw9p2C59/fgm35lzpJ/aJJMdMhce1a9fw7jvvyDloWOwNntgf77//vlTUHzhwQL6XL+Sl7955+2089NBDAkiwWoZJRs4npz8+LdJP/NwCMbduzYk8y2OPPmIMntsOUEGZHDJRbs7ekUrbyYkJAYzodUFGBUESMiq8P16AoRuYuNfvnDnf6sn2mby5r1Zquulu6u2byicm74L+ClqtGuq1CrKb68jnsmCCltJamQyNc6nVyioePq8ALl64hLOfnsPa2hKi0RD27t2D7dvG0KpXkErEUTYyMY88/jjSgxOIxUbpVINmKySyTNKPXuNJR/dWdyp+H6uuijh//hTWV5ewc8cUSoUSCGRV6zkMjwwK2+LA3icQDKTRaLbxj7/6OZYXPseLJ4+IXw6BiN17H0VmdAeuz87jpZd+iqmpMXznxe+h1Qjg4sXPcP7CWTx/8hjq9TZOnT4nUi579u7C4489ifk7K5iZViPtVruGGqvYW36MZMbwy5/9Da5eegt//Ef/Iz49fwnj23ZjZGwnlpbWcf7cWeyZnsRDD+/H2S/WcfX6bZz95FMB/GZ278LBg3uQSg4gFk2oRF5sAPFECqVyFaUiZXiauHntU6RTQTxy+HFkS2R/DQhQMTycFumnUqmOi2c/QiqxiePHnsbiUhilRkLe5cFkUoBDO8dRro+STFcvf4Hrdy4Kc2Nm70E8/fQRxGIZZVRs5lFrqu5uLpeTinq+19ajgslxxidkDuU2i7LZFOPgCJPUdWGeWaCCY31hfl4AOkr8cfyysi0UYHK/qpVb3FT6W6jWq7Kuch4RRoVUjQWQSSUlOb62to7BzKDI6LAqj9XwHMfZAs20o4hHY6hVlFFRLFeQpQ9RNCRAoZV+osQSN+HCsqzVkC8U5P4IVrDNqpOsBsnRGN9d4NbsvEg/ib9DlFVsDQndBGCOxRENhVApVRyggowK+36xTZQglOp6WVu4aaeXxTqaDV6vjsRAUpL4tUZFQBDxBAnpZpggBeclMv/4XTGgb/pkDadHBf0W2NZ6jeblNFannKKCHMLuI4ge0KpPK6nWIf10e1ESFARUY5GwrOmthk+Aio3NDUm8E6jgXGmBCp6rXGW7SkglkwK0cL4lUMENMaW26BvCZ8328E++gypdpYkobpobrNY0pqK6kRcUxyRDVJrBAtPSGUbCiZ+vra/Is6KZNqUeu4EKbuptfCQyBH410+ZGPJmkFwzHaFP6UeQaxD9E419rdklWIvz0/lhxigks+3FjYx3lgkqOCaNCCkp8KkGWSMi4eABU9EML7hNF+DqMin4blz6X7itd04cdrtml+7mP+z3+K5y+O3Etw/d++rzL18DTZ736Q3aREjf0ylj3vu793rVnV+7ueZ1Te9vrSV73aM+Xg0w9BsjXAipsn3uuyPnt/2XvzZ/kus4rwZNrZWbtO2oDCihsVVi5iKJEkZQtiaY87WVsy0sv0TGSe4vp/jfa88PE/DAT4+4OqXuieyJs2Q61ZEuURImiSYq7uC8AsaMA1IJas9as3CfO+e7NfJmVCaBkedyKQCooAFX53rvvvvvu/e53vnNOnURb5bfNwII7gAhuA+0a3GwAB36+104PXjtQJR0cS7tlh6r9F/xdMF6t6YLKNaq7fwMRTNLIMw64Nnq2RX0C1/rBMUmqUgsVqQ3dtmM/+2SxXaPxp1L17ySTeWolZen512h4OPBcEoUO1FCy16EIHhTnoVx7yBbgn/JhcAoG3MNzTWXfaq11rADvwcD7F4DvGA9sE9dTu12XPA+2jT+SLyeTyy6BLu+8oiksFC0hbYUEPi6x6nuui0z0c71j7GZeY9ZbvBzjJC8R7U3Ig93OYkN7JFbgx/8ot+3nCa8IYr8ngECTcK7FJmnMQhEvhch7ZjuMZc9kvOVfimIPmKS1l+mqyGLRy8FJKKmiP2+yzLyeCj/yth/1DEuT6jVmrNpKaWP2QbJFIAcLeBmPcS0nmMHfm7SXxWzMDzD38t/+i+1v+fnnX2PewGJDnluMHPmc2LD0e1Ur0CAIwH53nmyO2WJnqjIi9NycN4nmQwf0GAPH4me1jX0d8FyssJZEdKiyHXQ85cVczkgQThjy52BeSWNBsZjJPvEeyHiW0TzP72SSmRtiTkYMXgdyyGy8YL4c3hBdY8JLPzn/kvtARZNJ6P6Pf3l74N//k7Pu1W0ATAR+5Jc8Ta6eYxQ4UgtXDXXUDjYfZhcSueM8Il9lG/jp2mbtygJc/WJlQjdk2xla1/2+4YK3a+X0gIln19WaY9evtJXDd4Ez1c4Jsk+qhIxqBFMBaqon8/Ola/IdQj0XzFTvre67/p8GatvHGQZVvhlY8exr7tkEEOHAwwp0owFT/HZJi28A/GGVhtPX4yRLM0cz02YlaTOgwjwrJh95rAJU+M21T4yyr4JABRN41JamhjqTwZR+6uzpFVDByv5kPIb5GcpFFDA0MiQgg8+DutnJ1gBQMT+HbgIVvQZU8K7GJyZkqmqMCksuSB+cVZtFk+rwQIVGqNMGtO9aJScTGxwzTOj09fZJP5HAAJP3pWJem3N+uLjaZt66V9CYAyqKoYgBFTHSIAlUzAjIaCHLIZcVm4IA0eLi7YZARVuqFRMTh9DRvw/hWFQbeDNvotkqk85mcs42NAIquCB6RgWBimpg1YJyuGzGmAGgggDR4GAfMjsbqm4kK4avx9baOl5+6SUluKamTmDk4BEBFesEKuJRJSyMusu+tQpfL//kg0tVhLIqmfRgR51kFf/szKxjVJhhtNjfrppifSWN53/0Y3mEfPaxxzCyf0yJOo51Jth9woYJM8+o8JWmt29TS9+SxwQqmLCj9BPZLKlEQhXjlKxh8PGFz/+Kvktzdw4yBnqxGBPfZYFoFuiElKyMxuNItaWQSCUE7JDlcPXSZbz+2pv4wz/4A5x54AFs56xCmuOGfis0VR4WI4hBEQNDJnRiAsN+8P0fKVn9pS99CV3d7SgU89je2qqYmDLRqcAzRKmygkThvv3tv8b+kTF5VDAhR5ZNOr2sKugQfSXU3giy+Tw+/OADbKTT+MIXv6CkKRNTfCcZSDG5HYqF5YFw7epVPPKpR+TXwXdFldEu4CdQ8dJLL8mjgvJOPnnF8c5zEaigD8Xx48clb8IqYp7/pRdfxNTJk2Jh+PHHn7/z1lvYf+CAwA1VtZTLuHnjhirBT5yYlBwZ/QXeefsdnDl7SjI5hUIWl2im3d6O4aEhMYB+9vcEVATvr1kEwD4W/8dR8QkosQKJlUz0sQljDZnMOnaym4hFQ+jv61fFf6gcRmaHCXoG+y3o6x9AMtlmhrPLK3jnrXdw+fIlbG0sIxzOob+vDZ3tLUjECbaG5dGyb2g/Eq29SKYGEI62ooQYQg6sCLLqgps+Le/IIZ9dwztvv4orl84hn9lWwE7QaGhkADu5Mo4fewSxWA/mb9/GufPv4NyHL6O7PY4vfP4JJdJTHX1o7RrFYjqL8+fexofvvSFZp8ce+4w8W1577TXNvRzTl69ckwfE1IljaIm3orO9H309Y/J6yJe2BVhSvqqrrRvf+uZ/xc2rr0v6afZ2Gl19BxCKdSKd3sSrr7yAw+O9mJw8hIs3svjpyz/DuY8/UWL62NHDOHJkHC3xKFpIZQpTAi6FVFu7ZJ+2t3nPOdy49gF6ehKYOnMS6Y0SdrIEClrQ19cliZ2trRw+evs1dLal8bnPPYS5+Tiy5Q7EWyPoSNHPgjrDO5i9dRPXrl6RfBwT/5193RjcN4z9Bw6htbUTxDEzGbIMNvT+NQMqyKjgBiWXLYlRYdJPBCoo/VQQUMFNMAERvjvzc3MYGjaPCgMquBGMIJ/JWoUln2+krEQ9PRYoT8jdN78TjYQqUmBkDFC+iWshN9EEPzlO1rZo6pxCMp6QB0dLS1K/S2+sCUClR8xOJidmGUEMD1QQgKQ0F99Lb6bt52NO4x6ouHl9TmsD16qWpJlp8/2pABXxOLIOiCWjItJiGtacjwVUOCNt00hmQj5aA1RUpJ/yGTnveKCCfcVqQXoxeECdcy/XPTIBiuWcPHCMal8Uo4JrvwcqlDyIhjT/NgMqbs3cFlhMwCPhNtiUlqL0EwFkPqsgUCGwSuvrVgVASSZatZklUKHKQ5jBOZ+NdKijEQEVPunh2ZE+OeNBCv0ZADP4+5rkTyBzRaCCz4pAhe4NkYr0k62jVU15qwqMYHZ2TomxtrZW/eeBCkWfDqiwBIbJR3AcMy5bcEAFY0CtpS0tYstu0ay9xqOiClTQq0nSF3dgVGi+C8TBQRC66e7tbgnN4IGWMbqHjHf91faSgP85Tr8rdXin6/kNVZMe2WNTm6+JzU/UcCd0t+vW7H0Y1Niq2/Czl2caPEF9G5rJDdlGavelbeNqv73b/fhawUqZc4M7qZyjerJ7OG3NiRSvBtpV+WX9zwIn3lXF3/TlcVvRO70TdR3hd6WuFK7uzG5s+mft2mS5gto7rxlDDTu7OWhkz8fOV30bPGvCX7TatBqwwKcUdj2b4HvFJCn5nIGiRg8IBO645o4aAQDOm8PvyYOd5ZPFth/xe3ZXZOrzNG4v6pkFKm8MtNviwEbDuNoXVUayJV2DfdFoWAjYCIAzukZlTg6+xH7sOKNgAQmWQ5KHgCti9LJEKsAQpGffV9wjLwoDHXRbKtBh2y2J7U2Jdf/Ou4LnNRkjggwG3jNW98wCM8m2JLfken1cr6SzXZtJd0kOKVFv/hRM8Pu+EZhBpgd/RokitZUG4Hl5TjHXQWkmkxgyRoUq+6Mh8zIsmb+D/Y5xj/Ni4M8dqCOGaZgV+HkVlajdTuKc67iADBl/e1UCay/3wFSKYF+q79jfZIHsMK4gK7usNvDjvTPkh8Edg3wUGJdQjsueE4EID4Z5+a48C098p8Oki/g9xabsdwcQsA/5vL7xn6pFwX/8rwxg8WwKnobXUfGVS/QLBHH3ZaBSyYr0ClaoIUDDmddLiqlEDxMDuky2y95P89GIuHNRHoztcN4kAoBcEQhzP/SQUx8ZEKEYx7187BcWNRpQx343AMezSr0sVvCd5SbCwCLHGHFzEcc175/n9/4nzO3wRRWjp2T79ftAxV0Wpfu//uXrgT/5xwZU1CxLgXU1iOoGKU52RG3Svyme7k5SXfiqptPV6waWxdqLNujUxkvovfW+b7NNyPW33qwkwFdt1Cb/A1p1QcaGmBoKeVwy0N9voGOF4NTfh4sUggwUO03gU9/mXRG0D5caP9ddNxhsQz3nMRCQ+b/WeFRUJQPoJWCMCv7nzbTJoKAE1Ba2tg2koGfF5COspKUckRlv8+MZFfx7FagoSh6GiZ+N9Q1sbm9L+qm7p18ySWuracQjIczduqkkwvDoqOiMnPxrgIoLTvrJMSpoZloOh3D4yDFLKHea7rOSOkrskH5nTAoCFUr6u272CwwXZbZZJqPlsqpz6VFBoMKkn+hRQcNS86iwygJbjEVVZJAWNUZFORLFyMhBhKXXuImVpRkFSzQOLeSzyG1nFBjdXphDd0eQUVHCwQOHlJiYODyB9t4BROJWZZ8Xo6KkpIsHTrxHhaQ4nJm2wIIw75ta5Kx69PIithiGoiFVRxpQ0Ya1jQ1sb2yiv68XO7ktRGMRsUDYP1vrGwZUdHarQn7/xDEMEKhYp1GoMSrYb2RU1AMVlapUVoTSAIzBXxgynL1+7SrmZucw2NsHVqFThsjifAuI1paW8dwPf4Te7p4qUNFLeRcLShSIOD8Ffp/JKQ9eSKJCmtxWkUrJJ8q1UDOdbBGyIF548UVVfnz5qV9DT28vVpaWNSZz1P8sk9JrDB0GC6rqoZyPzGBTaOto03kZ4F29dAWvvvI6vvJ7v4e+gQGspFf1XUqSra+uqZ/H9+9HV3cXUm1Qsi8atSDrxz96XhXHBCr6B3sUhHL8892i7igTPd1dXWLAUFc+Ggrjm3/xV5J+euzRx/ROMUm2urqsv4cYVDmggiDjB++9j7WVFXzxS1/U7/l+MnHHD6ulO7q7lBhnf5ycOoH9o2NKrmoP4KpZCFS8+OKL8qg4dOiQq06x+YXBM422R8fGMDU5qeeRTq+KUfXiSy/h9OnTOHL4iIA6vm+s4CZQMTI2JqBCmxMHVGxvbWJyalJwH82N330nCFTkcPnKdVXa0g+D8nBvUvrpkUf073pGxb2tGQHwPDgTB9gUzTZp2ma4aV/bKVGCyqrefv75H6O7I4KTJ48oEd7amjCqca6sxHShTBYEwbwoBgaH0ZJgUprBa9TOsbWJmZvXcP7j9zE3O418fgupeBQ9XVHQm7Yl1Yp4sgN9+w6gu3sEqdZuhCNJhMK+SslYkJagtCmO58/trGNu5jI+/OANpJdn0dWaxMjQPkyePInl1RWsbmTwwNnPIxLtQqFcxvSNC9hOz+LZ734Lp08ewdmzJ9HeM4h4+xBml7ZRyuaxvjKH51/4HqZOHsEjjzwoyaP33zuP6Rszet4Hxvdj6sRxRMItaG/tw9DgQY37QimDAljBlpSs1Df/23/G2tLH+Hf/7p9jp5hCpKUXpVA7trM5PP/c9zA8GMfZ00cwuxzHn//5tzE3exuDAwM4duwwDowNqyI7TqAiRGp+Qh4VmUxWoAHH++z0OQwMtmLy9Cksr5FJ0IJIJCEJrq2dTWxt7uDDt19FT+cmPvMZSk4lsFPuQChWRCmbwcrKEm7euI7FhdtItMQxNLQP4+MH0do5KP8QSk3xnS4UylobV9Np5AqFpkAFwTcBFTslrKU3nV8SEI1z40hj5qqZNoGK2/PzklAjUMGPgGBqI2d2NMeF+f8RFhZk5XtkQEVZDDLOwWSRMTlMA+r29k6jz5fMUJqbqfWtLc2fBJPpURGPJ7Sup8moSHFDTqAii86ubhkbc8PHNd4DFWaybf4DnAOMzVAyI+5SCDen5yQHINmfJP1VipJ+8kBFikbYO1lVVi6vLCOWpE+DUfMJVJj0k1WcEajg5lBm2oWy1hxJP0Wj2MkZUME5zBcRcO3jukgZKluP4gJDGXsUSlmB/lxDuTckWMh3OAhUBKWfTLYprmo5YwpGQKCC83Yb5bzCIZNhKIRQpJRUmkBFxLyVCgWZaYuNEYkiQ4BMklStSLSklDygXKMqLymplNlUvBIEKjyjQnGVqyblePBJDgEVriqUv68HKoIeFcsrS1qzW9uM4RWlv5HzqLCiBtvA+zmwAlSUS5KeJKuCs4vkEN3mWxJ4bq0UcyLFeSkGMhzZRq5B/DPR0oL0WhrbGxsVRgXBG8YBnlFRlX4io6mxR0UleeCj4l2xd20yUWH3XjK/5kq8RyRhLxdwDd/rIbotf5D9Gbyv+v3dHZkLe732vS6ulVtrfAHDBBpCGI2voAOYBKzJsNt3fyH3UNufuxvR4CK6h+rPg99ouJv1+0dn8uwZSPWDck9jtK6h4tA3G7O1mfIGG8H6k7ksYN2PrY7fQKOm3vQ1SXEmPhs/qKaPLqjAELx+08fU5D31sZCldQNIxW6tAf8iNWtTyLEN6sdGDbBRYQeYj0GjT1UWx+15nAGvikIl4eqZutWjfdJTfV75cfWe62NV/28bS7sb0ii2lYyU+6ra4eZ/7W8bfQIeEjVTUqAw1YMWwetxf+RBd5/gVlKdhVZOSkgV6mHmEBy44FgHbIaMql376pvl5RBVqBYAE7i2CPBwbGiuQyYF5OL3ui7iM/CST6rwJ4jhzJArlfVM8pdKWs/kXyHAxDJEjAOY0Ja3ZjZnfhxOdld9Iplohvyuzz34RN8+Si0RjHD7XPYF2egschPowv22q+6XaoJ8ASlNVB3jKmYgQOCAI+51mcRXPkfm3vQvI3BgU5h/3qrudzKOigPEgjAmgrErDEAQ08HJSHkJMoEM8ifxcYMDR1xcwDHM478RkH76439hEl8CaFzxs/wiCEj4/iYQwMKbWAyRkPWrf740USc4xMI6AT3MWZUKLvY0wIV9pfxJzo7TG1EB1AyAENhCWWdn6q2CPXlNmN+JAXgWTyv/4Bg9/BnHLdtnKh3exNzNeE4O2+SqDVgx4MS/l/Z3+YrYYBTAorEWoYCDM/6+L/3UeA66/9Nf3h4woCIAIbi/Ngtma5fsWvGnuwEV1YWzGopUzxBYUhuudYEf1gWtZvC9l09V5qiC6PvTNwsYKowKfx0DGiqL6t2ACh1mqKzNfkHApHGA4GBZF+AGO8WtVM1id17CTXK1AFSjm/MPnMf8HYAKSj/RTPsegIrjj3yuKv3EClFHPdTkTaESehmIrVGQJE4+l8UmJYe2NtHa1o6enj4kUimsLK+gkKUh8m309PVhaHhElQqkfzI5wiQOPSouf/IJVhfmlGSuMCrCYRw9Pqlrt3f3SKaHiwgXdv5ZlH5iTkkQr4FpSL0tcsaoKEgCgp+2tg709vQoCaUK+51tq3rf3LaqCUkF2eZc74kqNaLYpp9AJIbR0XGEIwQqNrC0dEuBQdIDFTTJDIUwPz+Lrq5OVd6f/+hjhuX3MgAAIABJREFUmfBOHJpQn0xMHEZ7b7+Al1jc6JVclCn9VC7lxfDg4s0EFpMxhsz7xAWraatAhU9aMABiZQN9HCjxwuuk0+vIbG2jv6cHlLdiQMR7ZaKIAMYrNNPu6MDxySmM06NCjIo1VRWzLZL1IUukjlFhVagmV0EpK/VTGNI/v3rlCpYWF9HX1WPvD9msru3s1/TiEn70zLPo6+3BZx93jIpeY1R43VQGD6yW5TU4vgRUFEsyuVZgQfaGgIoIQqWiZHXo83rlyiW89OLLiEXi+LWnv4yR4VEHsmWUQKGsldGFQ0qe8U/2H5OUShY5Iy4mtC5duIgXX3gJX/nK72EnV0CuXJJshRLzm9uSiLKKkTK6OqM4e/YMDhw4qMTdsz/8MYqlkECAgX29CmTY73wvaCTPMdrZ0amkXhel0cJR/Pk3/wKj+4bwqYcfURUz9f5X08ugBwyDNb7vrBrmsfTioPTQl556qgJUsC2c35hkbEkm5VFx9cplPP65z0lWiePfqpDoCVPA5YuX8NJLP8VT9Kg4eFDviZJ3DNQKRflX0DD7xBRlmyzRvrG9hZ/87fN44MwZHDt8VMwospnWN7fw6suvYXRsBCMjZJlYQHvzJmXetjA1dZzOtdpAvPXW23jggbPSfmdVydXr02hNpQyocNJPHqiISb/VfdzGtBIQ+k1fcCmpyXXsnj8rm6vAMdpEukAysFpUfsYgeHVlBS/87U8QDm3jH/2jp9FHqTIG+gUG0yY7Q14M5wgG7e0dnejs7BagaBqoRmfnbJLnHHh7Hjemr2P6+lWsrFxHsUjPnhQ6umiITBPeDgz09aGjowvtHYNIpDoRitK3hJU4tgoTdFtJz+HyxXO4cuk88tkNjI3sw4njRzV2Ozp70d5Nk/sSJo6cRTTaLbmW1fQStjfmcO7dt3Dp3Ht46KGHcPzEabT1DmF2ZQOlQgnDA/14/vkf4c03X8RnP/sQHn7oLOZmF/DKa+8imy3iwIH9OD45iWikBQMDo0glaeLNZ55X1RMZa1cuXMGPnvk2UJzF//pv/zkKkX1ApA3FUBL5AvDCT55BW2IbDz1wGJv5Xvxf/+c3kN0p4MCBMRw9NoGB/j71LZkaGvvRGNo6upSEZ/J7c30Nt26cw9BQN46feADL6SIyO3FEIwn09lH6aUtyZR+99xL6u/P47KOfwq1bOSylC7i9PIeFxRn5GXS2d2HfviGMjewXK4FV/bky16UiWlvb9G96KG1mtrG8uqoxT5YCgQYmaLlRomQB359UqkWbxhz9LCj9lDNvBW1EywUlr7kZWllaxdraOhYX5jEmRlm3AACftKefBDcyTHwzdZQvWgGAfJhYBR/jGhDV+ehBQcYAzcYJvDNWYR9xXPO9pHRcsiWJnQy9NVICKtY2zKOCyf/trQy6urrhpZ84r9JEkX3X3d2te/QawJboJ+MwJuPqmVu35e/BqkKC2/Qj4jzDebs1lUSqJSlvDPbJ8tKSPICsys8YblrDA5KC7EMyeDiHmqdEq8ADrofsH5qRe6CC0lv8DhPyBDxMGzgs6TAWLBDA4DVoLL+0uKR5yHtPeeknSi6wKpFxCIGKFg9UhMKYnVnQ2tDaRvAJkuRiUSXHxcrqstrFeZrrwczMLWk9cw0heMt5jEn/VDKJaIzsTGNV0Gdie2cLuUIOme1tPV8v/eSrRq0IxFVCSnvaNtGhOCsATTpAsoN63/zO3Ipt+MzpG8Fx0tZuQIXALief4BMqwXwn+1+MCgEVSbFE2Ne+qMODJZwb2d8qHkglFf8QqOCa0ZpqVQInkTDQLLO96QCfqpk2xwzHUofWszDCO20GVMRbBLB5qQsxL11hQ2U+vmsx1M+RHN8jUHGnfUvTBPSetjreCLe+gjxoHhpc7IJgTYP91J6uvZf9mNsSNcnW7nl7Z6Ikf89ARZNk951uu77/7oAy2PbQPycvOezBDp+p/LvhLr9QoKLhfVtGgEBF8BkGt9q7n+0/IFDh2AYWvwX2avWm5k0Ap5o36RcEVLhR4NQqquBJc5ElJkobASsGFnngoybEbTAOm4EZOoeTMrIQt1HQXD07n7UlbysVjtXw2+Up/LWCQEUFiHGgg0+OGyPBywxZQthYee55uZjeGBiWNDYnw93FRn5P4aV1Ktd0cjtaU5w0st8vW+NrEy+qPfIyWJJb9Ilma5MkGhnbO2Nqk3ayvbfWP5fQZlxKSSif6GcOgybYJvfDfZQBMTXqJs7noqZ9LscgiSrnxefbLbaFuwetwyEm063QQ74bMHNqtttLOXlApwqAGZtAPpIs4gyFxJDX3kQ5Ma7rOfl2Mu7Q+suiMhZPOoaLxoXWYNszqyi0aOwH3iPBHH73G9+oelR87Y+NZSKJTQdksJhJElchKwxhTkLMmTDzOMaQsPYbeMS4X3t8shOYe5ExdlExppgtTpaKQ1Oyys6sm9eMhLn3gvYjZMQzZmdOQeck08fJbvFPFc/IS6TKvmA8wudphazmF2LvkIFAlocIoVC2eFaFj041gn3POF8FHjA1D+tXA+MiMTKIjMVzn1Gx99jj/hH/g/fAn/xjb6ZdW+Bvi0cjAMMn2P10FwAY7liuUl3QgtJDHsUNLm2Ni2cCCfVdpMQmPMVdS4pdJejtUFlsfQOaJP9rfR+qi1Ul9mwAVPhjqkmrYNVJIGHm+Zm7xko9OBFsZPN7rj6GYBDBvzcBKio/bsTy8H3mrl3DqLDKA06OFY8Kh8IzecEkMxkUlE7Q392/jzmgwlf2+wVbAYcDKlhxyH8zqU3AgDI36+sbqpTu6+tHKpUEZXu4iWXCYHhsv5LiXAxoPk26Ije7lPO4eP48Vhdvo6enF919fXr+5XAYxyanDKjo7VGg4ys3rIqUJqg7yOcNqNAC6dB+v0Cwmp3a25KpiCclN8TkDBdneVSU8mJU8OM1x3msJQTKCEcj2MrkEYrEMHaAid0Ytrc2sLB0UxJEZFQUszu6B1bozM/PoaunF+mVZZz74H0UczkcPnJUprCUseru7ZfPRSyeVJUuq2W72lmFbUAFF3K2kYFIFXzhAkwQJaoFnX3paausnGWfzM/NYof63p1dWFldRXY7i/7uXjFnmOCi9BNBke31DZlpd7S3YXLqBA4eOY7egUFV5NOgVdrfTOSLeUMjZQYNlpDzbBYl5xIJt8EhULGNy5cuYXNjHZ2pdgt0rDTdnhdCWF9ZwY+e+SH6envx2JOfk/QTWQr8rlVwmFYlE/u8DpOFFuAWsHB7UWM4ErYAjcEWKM+RoARYGVeuXMSLP3kJLfEUnv7138BA/7BMusngyRWyYLXp6vKSqlkVMMiUPYZUC81BTRuUCSgyHsjeeO655/Dbv/1bYhiFEy1qC68rQ9qVFZMfyWQQCe3gwP4xnDnzgAKTl195VUnBRx99FOMT+wWUUVqM19zYXEd6ZUVBTDZfxPDImBJW3/zmNzE0sE+ABxNgLS1RyS1Rp52AmlW1tEgq6r333sFaehVP/ZoBFRwDFjxakMcq/gufnMfVq1fw5JNPoK/fwJJcnolTqyhhMpseFU998Us4dPCgnlEoymQaUMzlDagYHcOpkycFvvLcK+tr+N6zP8SnHjqLqYNHEGLQGKJpbxZ/+5MXMTY2jKHhQdMcLQIzt+YlpzY5eVzvFdv41ltv4cEHH1QAys+161VGBZO/ZFR8Wh4VQ4ip8rU60frNicZKIHlVcRWqw5X9kX5j4iLNmsUzuGkRgFV3PRoVky3z/vvvyhT76aefRn//ICJkOpQ5z/A+KH1WreIiaNjXR2k5Ayok7+c2jDJo42aDieT1dczMXMf1659gZu4qlpcXkIonMdDTjn29lK4Jo6tnCG1dg2jrHkJrW5/GNhOVt25exUfnXhezhwm/iUOHcfTIcfR09+H27UWc//g8Yok8Dk4Mo6uHUlQDCIeSWE2vYHN7Huc+fA/rt5c1Fj/z2ccwdOAAVre3lEwe7BvD+2+fx4+ffQaxeAaPfvoUTp88gevTC/jk4k10tHdiauoUwpEWjV9DI7mh4xjMYm5uFm+//iauXvwIHR05fO2r/xih1ASKoShKISZ8o3j95RdQ2JnBgw+MI5Laj//jf/9PiERacPjwIRyaGJM5dyFPMJSn5+Ygis7eXtBLgl5I66tLuHXzY4yODuLwkYewnAZ2ctxcJGSUzfVrY3sVH77/HHo6yvj0w5/Gcz96E/OLa9jY2UbfYDcOHz6G0ZFxtLdTvosygNwQFVGMljSPt6XaNfewNoxAxdLqCsoFAqNmVMh3j/OaT4C3JZl8J42+jLX0FrazO6qi5x6sgJzJ6pRCWFlMY2VlFctLCxgfH0NXF5PDtlHlBowyT5wrWdFHIL9YNgakf8c5L/KaPB9BEo5RyjoRqOD8Q6CCnw0m5xMJJdG3M9tqNyWQOO4o1cShzvugfBmT+pR+4u8pq7e5ZUAFWRUCSJz2NNdeGkUSqJifW0J2J2egQ4xzhwEVYqglCFQktClm8mF5aVkye359Zvt9hV+QOcD2cGMoEKLVzLRzbkPLeZnzM7/Pe+Z3OFdW9aJDujeBzwkDKggQMPbwjArP7JMcAJ8sY4mWmCojKd/I/5gQmL1lMoMER/gxGQvTKSaAzPZzXmBcRKCCIDbXbMYQlM0i44qJf67VVr0XU0o2k8vIc4TygXECFamqR4VVOhYFaklCwplkUqYK7HMmkBiPsNqQxqaS7Kbuu69SLWJxaUn3b94dbkOuZIhVMgY/IcqylkMOqCgi1Zo0kFxAhUlUBZ8N75Vjj+BXOBLwqEhaUQOfDYGmrW16VND/xYAKgkGeUUFg5q5AhepwgvsZv5+4U/a9eeHO7lB974yK/1+Aiib7z2pysObp3Zly8A8KVHCk+0IvlakE2hoEWJQWdXudmiqDuo3M32Vj7kGKvXZIY9ZBM+oO53lfTVspqKvblzdjadzL3f19AxU2xsrmIRHoqv/RgQqjGptihCX2g4n/uvixSUeHmhl5BySSvP6/pIjuMpTUl4E21QMJwWY0AiqU5tY1dl+o2bnuBFY0um0l/uvOXwNUVC5fbYP/WyUOdycmE0FmxG698KACz8eELNdASzzDGAQV3yOTbdLeg8+vDrTZfa8mZyQwwRWsMf7xkrdsh6SbxAQ04KG+Cw3b974Dljj2wIqYBI6xzFtj21kwyPOy4ICKESxckZeCK7JUNb5T1WB/ipFgntFOvqoKvNh1uDeydZjnUB0k9wOWXAswuewezdPLckMGfDg2tZNwtOdo41/MSwe0+OS4/u2ACvNMC6tAJyGlAidJxXNKXsr2KQJI3PV0Tfe8lICXXyX38yad5OM5FlT86Z9WR9rX/phG2QYeWf7C+sE/ExaX6pmH7BzsL4EtPGfe/CwkFVVgvsqMvkMRvuNklBpLw/e79z2TF4UDubw8le9XjT/5WEQryiC2V656cPF+9PwcY8cfY/JVXnHFvm9sFP+S+DfDWBz8vn/G3B8SKLFYN6KCWO0JCKqxOPI+o+Jelr/73/ll6oF//0dnAjqBeu0DL4u/k/rsfS1Ysaf7rSSD/ATql7Jqrqfxmt0saW8vdqMKg6oOZKMWVq9bmewaoO7VIwPAQEXKKmB11gyocBTNWnYEz9pgE6TAdDdSYjhGoL2Vr9T3lFvAqsuMNd9/vyEIYwtvYGlyx9R+uQrIuDbKgMgmYf65F6Di+KcfrzAqvEYx/+SmlVRkVrzHJBFkQAUXcy6EZC/wd/v2DWrTymQBK/C4loweOICuvgFN3pzEs9sZfbcKVCygp7cHPb39klNhMuHY1AkZSnb0dlc2z1wEPVDB5AorP62NpleoJ8eFOZOxxU7GjpSLiotRwcWWFfZmGF2QNA8/2ly7Sk8DKkryCSBQwcre0f3jSlSSUXF78QailD2gtmJ2R0neciGv++3o7sXa6hLOf/iBgIqJw0fQ2tohoKKLHhmJJGLxlCrcCVTQYLdczEo6Ip5oQX9/vzMxN7NtJVkC0k9M6ug5OH1oAyrm5MHQ2tEpqZLM1g729fYr+RNriQqoKBUK0pF+7eWX0dnRLqBifOIYegYGsLG1IakSJcEYZOTyqhzxQIX3BvFyFZTwUJVHKITN7S1cvHBBwFNHqk39Ruknf6yAiuUVPPvMDwRUPP4rj2NodLQCVDB4sYQuJUgySvCzUpjPjNqY83MLVmmbiFd0JsHq2STlsEq4dvWygIpYNIH/6Td+G709g2KDtLYzicQqhjwWFhckB8WElupcafzawqpZmrrnTP5DBmAlnD9/HseOHpXfSjyZQFtHhxJvHCesiGbya2tzEyjT3JdmpJ2qkL1x45YYAvR3ODCxHwgV0d/bK5YOq8FXV5Z1XK5QxNDQiMbwn/3Zn+Hg/gM4c+aMEmw0cd3cXNf9e/34ZkAF32sPWNmoj+CTT85LhusJB1SwT1klU0ZE78mlCxcERnzpC180oILjKxY1L5t8Aa++bIyK0ydPVkxe01ub+OvvP4NHHn4AUwcPI0RabKiM7WweLzz/U+zbN4DhkQE9Q1J3b94woIKMClXF5PN4++23cfbsWZORCUG+IkyO0Ty7HqiIB/MbgWVBEgV7ACqCGx7NjYFjg7/jlEEZruDHJzipS7+yOo8DYwSeYpKaYRAqo1yEUYT5zPDD+Y5ABcFDA02tKstL5vmNHMcYf0b/mOWVGXx87iN88M77KGU30NqSQ1dXAj29fejo6UNrey9a2zrR2d6BzOYW3n33HSytLWGwfwSTU2cwOjKBVIqAX4ue/1r6Nl559fuIJ4o4ffoMerqGJUVze2EW28UtvPf22+hra8Pl8xf0bB569BGEW2Lo7O3DQN8BnP/wGp778Q/R3RPF/Nwl/MqTj+P45FncnFmQx8ToyEF0dvWjo9OYD7zBUjGDmfmreO/9n+HqhctYmL2Jg/v78NWv/TMgOQ76+5SZsC1Fcf6DdzB74z088qkJtPcdwde//k2US1FMTIxjZHQfUqkOFHKm5QrSzsNsW6/kwfLZbawszmF25mMcODiEQxMPYMUBFQQfe7o75RW0uHATH3/0AkaG2mT8/V//61+jo2cIYwcPYXRsFEP7RhCPk+FRAovNuCkiEFiKlmU+TfBcVV5M6PN8K8tgUoPvJ8F4sgD5fC3pHkZ7KiWwIUuPivQmtrIZW6sikG9Cqi2pBP/ywqq8GFaWF3Dw4P4AUEHANQBU0OCalVdONoDvj5dg4vvDRD4NkzkXsWLMquQi8uVhAmBzi+tIQuPQezRwPFPej0aJzYAKMio8UMEKe16rApajLKk9PvPbc8tOwihqvhWlvNiNXBuSvG48ocIFPhPOuZxb/cbWm5D7RLgvLiCTg3MkvyepJwIV+axiHt6HZ1SIeZHPiwEQBCo4h/DnPJb9QZCAa3GGZtrOe8o2jdxRlgSkh+NRJSQIUsSjlCEIYebmbc173n9BkauLodJrq2Ky8Npcf2dnZzRWyCwhULG2vo7W1hYVaDDm4PzAubtQKiNbzAoIItMxHq4yKsQadGbaGvMCuMioiCAcDaMcM61qxiNg9V+hRLRWiV4CGwQDeDyBCvZdRwcBbkvi+KKNeqBCbAsCFTP0qDCgwjMqTPqJbbBkAz/sV0lcsR/DUSwtOTNtjj3KZ0WimsM3tyn9FAQqbE7kucnAlDG4GBUtjRkVXjfaTcSVxO8dNy97BSqa+CI0vUZTIfjmrdpTbtwb59afrsoE/6WQfvIMiZq9aU26uwFoUddRlYzoHR/4Pf6SJ2uSXG5S6FbZiDViUTRhVvgEvyqE/YNyQEUQmvGJdA+f3ONNKA3PeKvhp6b7GgA+d7hIbWy0u1XNgAr7eTBZV3uRpkP/bvew68DmPVUTu7mktCVzPRBpbaqmEZt0RFOgInC0e6bybrgbUOG+4MGTvQAVVp+oevxKY2uekRt/jebEO13Hr18CBpp8gkBF5bkHpr36zE2FOSHZIq5PVY9B9pMknpwclNYSmVhX2X+qnJe+oCXa9W4EcipBYERgiJM0smS8AQzesFgJ8SKlfVncEtZ1G2E9kupxng/GYnTS3/K0NLYAP/JtyDNBbvflAQsVajo5K7FHnYcE1zfv4SmJozoZOKkFsNjDGVCz4E3/dowBDi8m6G3EGcBmLFHLJ0k2SJ4cZgCtPTIT+k7CmPeqIhcWhojBWQX7ud/TnoksCDErrN00+OZ5WFSys8NCRgNlvKSSYk8yA1yRoVdvsHbZfs7iA54rj69/vcqo8NJPnlGhUS0zcEovs2jOmDW8f3r7sW16vgG5Ki97VelnEKTi9i2ifTjjLT+cTTGAsSnlxKusCxb5+HFq74w9Y0lG0WSc/czYSx4nJaX6qGCgvI+T+vJm3EGZKL1rFQlN5i0a5QLNj4VMFstJ2XO06xnD6D5Qca8r4P3v/dL0wJ/84ZlKDOUb7RfDGmEnv6hW7syjmXe+1crEHnjn7LyuWsFw2+pJmgZ6zYEKX7mxqyUOVa//uWmGV88XDNYbxox1baou6M3a5FFYp81pkGhdhNNoE+Tpma7FLp6STEvNp4EwpX5fdw2Hmtc8sl396ysEOEnWIRp6TB78cGfRZGsBQAWooJm2FqO8jEG5YFYZFTuqsKwyKnYw+egTDqigBBErCsL6N/8rUxqB8hdRJj/zJk+RL6gilHIUTOgMjwypopOSRNTkptb48P4DMtlWVUIup027ByoufUJGxYIYFT19/WJTcHU6NmWMCgIVqkQgCBGyJJEl+2g2SskgM2H2ixP/zd8rMVO2qm6aXNLM2QyTuKjlZZy0ITPtsqpUfbWnX4wqQAWlnwhUSPppHbcXHFBBf4J8FqVcAYXcDhYWbqO9uxfr6WWc//BDB1QcRmuqA+OHPVCRQjzRqufBivv2tgSKhSxWlimTkcTIyIj0F+VR4eQQgmbaZiiaVfLAAwjsY3p+pNo7lDDZ2tjGcP+g+ofyHJSmCAIVXZ0dmDpxEmPjh9E/NIT1zQ1EYtQ/b0XcAUkMKtj30lB3Jua+j5l4EM0xGsZKOo0Ln3yiYKcj2WrBkQcqWAmLkDwqfvi970s+58lffVJARZekT5h/qQIVrKLlWGMCjpXCZFTcnl+UrEZbKwOrHZM6KRXQ1hpHJFrE9LWreOEnL4n2+Zu/9bvo6R4QGEBpKFYQM/lD+SeCY5Qi21yncXa+Ql5i1SdNyvgesXqXCT1en682GTU0PWZww2QfEzJsA//Oem+CS0wQMiCZn7+No0eP4fCRw4jGyurPhx605HyxkMeOkoXrAuFoUkxg4K/+8i8xNTmFhx58UMEhjb8zO5ti4LBKnIHQ3RgVXg+U45pABeWFHn/icTEqOM49o4LvwMULF+VD8aVf/YI8Kjg/RKilz+dAoOKVV5SUp0eFr+RZy2zh29/9Lj798IMOqCgiH6KGPvDTl15FTy9ldPpcpQ2Billsbm7j5MmpCmX4nXfewcmTJzU38HPl6hXNIcPDw3q2b7z5ZoVREWdVVN1s6iuIigEC2t0YFcFT1G97LTh2SaI6oCJYIUYgM0TzXUmGmRSXGBWODl0KsSrIZCz4bpANxcScJWKrtGbP4LCgnwXSIRTLDJizMh6fvjqNF3/8I4yNdmJ29hOsry2jo7MTvX0DmrMIZjKRqmRzWwqTU2fR0zuKUKgd5VAriuUWIBRHqLSN119/FhcuvIOhfYM4c+oBySml1xaRQREff/ghkpEINlfSWJifR2dXBx54+EHsGx1HMtGP69du43t/8x10dUUxv3BFSdfPfvZzOHT4KFZXN9ES70BP9xAiMTI8WGUErK7exM/efQEbm0tYX93A9OWrGBsawD/7p/8UkfaxClABxDE3fRXvvfVjPPzwOAb2T+Hb3/4J8rkQ9o+NobevWwyBQp5ANuX2IghFWtDV04eNjTXsbG1ieWEW87c/xqGJYYyPn8bqOhlKVr0dCwPXLl3G1YsfY3PzGh56cBJnzj6C9z+cQWf/AaQ6usWWoLSQqv3IMszlKwB+MVxGLpNTUlUAEyV7slksLC85T5yE3nuB9DHzGeKmq52SOKGw5LHSq5vIcL3URo6pBxozJ8U0Wl5YNqBi5TYOCajo0NiJU4KIifkd84KitwQ3YJxfvQSgByq4Ief1KaHGc1HOUAwzhLG1uVUDVPB7BCq4ifNARZw+E+VyhVHB35FRoTktsy2ggowBvpt+82cSDWUkKPNUimDh9goy2zt6t5nkzheyCktUdR9vQYpABWUFCFQsr+wCKvx64ll6fNnpMcE2eKBC/UEmWBCooESUY1T4d8wn4zmHcE0km1PgByKSQ6L0FSUNZZjpgAq+lkwwhmIRRGIxsSIFVCCEWzfnFTfwPB5E0BpVLGJ9w2Ib/o7X8kBFC/t3yxgryVRc8lPcTLNTYlEDxHIsRNjZxs7WtiT/CHCY94fJCWizrOpKyk2abCXX1hL/c0CFMSoo9mzyMoVyXuOe8xWBCmOaGMDkCxl8PBRMZhGo4P8aARVBRgX7ix+eV2weSoBFojLT5qab0n3UgGYSRfKG2xsuJmEhgAF17C8+KzJPuL7+ooGK3SvF3fY6ewQq7pDg2+1f5/cEe0Iq3PpR3dlplxAosv2HAyoa3EczKaSQG7/1e6CadHF96nivQMXe+rUpUBHYhu0aLY0ucUf5p6pcjt9zWtwUiGAq52xcrHfnEcsp4RcFVPg9b21k5H66K+bStxridP+wQIUv2gt6VKjPA/0UfIxN0xXNnmsw0x0AnyxJ2fhpBeWaKnOuvtzYO0PJz0av112Aisos0aToxv/ez/dBUMEOMZnXhvCuXuHdjaoIUgWMtX3sLENsV2WuGJeJWAEVlEKyfbYZQzNxXJX3s6p1J6mjbqo+pWALFIs7qV7vK6FiQsfM5jmUkxBDwZLejRgVvHffTi/VE+xLS/Bbop+eD3w4XkTD7wfMo6JF+1yLO6wXBQCIWVKVrgoCSv7++V2TLo5qXZRpNmUCSua/QUlgFsrw3kw2icX+wrmBAAAgAElEQVR+ZEtE1AcsbKRfIAs3xBCQkoVriyRouTcxhQKxHmgcTm9GzwJQwaM3/6bxN2XAc5XCKoIWAhgCY9AYLF76yQrjmIeR/FOpjFwhj298w/vpAf/yXxlwwA+fP/ucBSjsWMpmsY2URlWM44q5NM0QK6APSI5ADlkWJqfLWJWFlsyVKJ8lyWcyhXeseJfjht9hkSFZqc7zg0CFlwuzYjljazDet3FCVYWowAn+PJOlHxqZNiX1PwtDVfzqZbmcDJjfhzIHprHuc2+OkWNynw6Ic0WmnAHYLu3v6a9Kxv19RsXdlr37v/9l64FGQEXwHipB0S6gohqR1bDL7tQBlfWiNsFfD1Q4lmNQecqAjQrtdVeq6c6U5UCbtLjaMhagjlW/0LSCoDaiN2Jczc+CbWoEVLhrVlbKRjJLu4EK3rKvPqvtkCZSTjUobF0/NYwg/HcaABWBoDsQD7uqAk70ATNtxzzIEqy4C1BBRgUXJSY4fEUd/1T1gGR1kmJUcPIt5HfkM8GKeiYmuHEfHBxQsuPKlSuSa+jo6MS+kVF5Tag6IZsVUMHzUM/66qWLSC8tOqCiD2Wi26EQHnjoYVULdPX3ucoKBi4mQ8RxwCp3/sngwict2Ga2XUbHlD3K5owGGUugr5fniRiqTh1DelRktq1qgcl4Ji+UyXCBDz0qdkjbi+DAwQkZvG5vUWf8FuKxKFp4LgI1DG5KBczPzaOjj0DFqpN+yuLw4aNItbbj4OHD6OjuQaK1DZFoQoFJoZBDZ3sK2cwW5uZmJBs1TL1/VmHSxNwbUoeZzIorKGPySfqJznSaQ2BudlbeI62dBCo2ZPg12N2vJHAiGdcxZBZsptfwKhkV7e04dfoURg8cxr7RUQEVlJKQGWg0JpYMz8dFmwu6p2jKiIzSXwnqVdMoFNJw/+TceSUt21vbFaTmS0UliETJLRSxvrJaASo+/4XPY0SG1N0KikQHFR2VZqNbeo6UW7L7zWN+3tgQnZ3tCj7iMQaLWQMqIkVMX7+Cn77wimQ2fvO3fkeyLjT4DkfKAmlicVZ8risRT3COCamlpSVVXzM447NPphIKeAgQMHFMw1TOeZFYVOAFgzr2PY/XcbmcjLxZ1by8vKyg6tq1aYEO1PHPZNc1lh566EFp0ecpM+YqoxnJr66tafw/88wzePDMWXz6059W8JfJbCK9tiJDWUuoxgRU0Ez4gw/ew8Z6Wh4VfG/YF77aRQFaOCagYvr6NTEqevt6FNip4rkUVtDH50Tpp1/70lOYOHTI3ikGuOGQZEne+tlbGB0elvSTBakhZMtF/NV3voUHTp/CyYmjjOZQpA5oOYyXX3pFye7BQQIVZAoQqJgTUHHihIEdbOO7775bYY3wZ1evXdX8UPGooJn2pz6lf3OE3StQEYTQ75QG8EBFbZWNrSm8llms2acCYAhEN3q0Z0jYmmIVMyaZYHItOk8opKQcZXMsCWnrF88nOrcz37N/m+5sKZQzun8+jLffeA3LS9fxwNkjuHL5Y3z04fuSLGtNJjWf9vcPoKOzFeGWPNo6etA/OI6e3jGEo9TM57uWQH5nBx988CqyOytm5r2ZwdTUEYQiOYSTLbh86Qp2NreQirUgEY3quUxNTeLI8RPo7BpGNhPCN77+dZw8NY7MzopkyCgl99SXn8bw8AEUcmF0dw+hHIqjVIggn6Ph9ou4MXMBI6ODGB0+iDde/hmW5m/iN37zNzA0flZARUlPNY7ttRU898M/x6mT+zB27CQ+eP8q5mc3MDoyhu5uVskzycoqMxqVQ5r4ZHyRiUSgYu7WdSwtn8eRo/sxMjaJ9c0wVlYzuHL1Mm7dvIaNlTUkI0yar+GRR07hoYcfw9xiEVuFOBKpLqQS7UoSc+7yjCST2cuD+l/ZTBatyVZbN8vAdi4rRoUkoVpbNZ96toEZMBtQwZGys1MUo4JABTd88XhEvgRkYHADtLK0gsXFRaTTizh4aAzdHe2a/1gRJwNHsuQo/cTNsID0qvST9wkw6SfKBoVVFEAvG9MpDlUYFWsbnPOT2gz7tZtr4tpaGh6o4HrQ2dFthQJ5Su7tILOzLY8KeiTx574q35gjTLpHxAxZXFhVYp7rjxgVlP6i1rIYFUkl/gm6sF2eUeFjNp7Ls/J8UoFrDJkSXLM8K0KmlWRU0CNIwIwBnEHmhE+k2/qf1X+cFy02Ddsc72T9qgwOshWMLBtmYQLX8HiLWBWcAwiyci73PiQWJ9jGnyAON/7qM0o/zc6AJtHs6411yl6uoa2d/U4PKvonUZIrpnU+W8ypjwlWE6hg4t5LKvq5wXbrnEcscRFPxFCOccNckPSF2BRO/kmeFWGCnpacmb99uyL9VDHJDCSdfNUr5yjPqLh1a8Z5gCQdg8QArGDCp1pJSo+KlEB2MmSZZGAhCtkqZFTw+W1sres5cawQqCCb0TOA+M5VpZ/2zqjYKyDRbItDyaw9ffYKVNwhqd20TbuuUbv63TNQsdc8/h074l6S45UVc7eM05462S+8dX/uOkezG2yWPW7w86ZZ6wbXvodnaUm93QBMZbwGk94WXdytMH/XXe8dqLjzQKjeVvV7rrRt91OrByp4iEApu5f6T9Mr3w1sqTkw2KcNBlI9CuF9zJoBFbvyAu6cjTwqgptoi+oq93onoMLHjUFCkR8bjTIhaMLQCI6OYJ6jPudRz6xo9t0gUO2P0X7LW+MEu9ebN9epVlBG1/JHFgd7ljAPlbytAljH+lMczPjWJ+/tGAMxXCK/zi+Cm0ixkx0zQ4bDgThcMbTYhpaUNtYDwYlq3G2Sssa48GbRVsPpclINDMEDWRXFZ54VpTWSwIb2VyZfxHiR32Fuw5s4M+HMv/viPTEYXJuqwIW9K9w7Gss2osINnptJecZ+jD0lFRmmVwMLJmMuP2GFVJ4hyRZSbppAhMkgGZtCJtGSq4ZiRnaTP5/kmx1rk+exWIPPhLGcsVo8aCTvUOdnoep/Sl46nwV/HX9N7evc+/Mf/1O1SPdf/su84hWeX0U4MZMalZk6zynk0xL53JuyTbwXk3am+oEBWpUxo2LpojwRqUDAc/F3xbxJgUmyibmDStFZSFJR3KKZZwSlnr3fiMvreEaEk3WSHCi9TVmgqeJRA9f09lPCybFt5OUoA3dXiOHGSBWsIKhEJoUVnoiR4uYeHkOgSYCq5Jb3PfILXa5/nvX2/jH3e+AX2QN/8keOUXGHk9YzKzyr0YgCQVf6ZidpFMG5nwUWen+d6oJq3/FofXXBbLg8NwiEvAbc7ut7nwp/7mpxQ+NXvCZ+qbTZn7fR/VUDonoGRhVwqTbZMcgCEkwWqhmN0Cevqn3hg7na1ta1o546ptW1riInyPTg92tO4RNm1hajUroQUgkxB1TQeJqMCrIpPKNiZ8d5VNQxKjIZTH7mSS0CTHBwkfWLJzfbPClRbTIqlOzJm/QTEw1M2rLCk5IuTKh89NFH+g6NO3sHB9He2a0FJsio4Ob9ysVaoILZBMq8PPjwpyTf0DXQpwWJo8UDFVzsCFTw2akKwlX/sY2q4kvRB4LgitEtCVT09/VpEdfmv5hHoWjJZ6tmDzIqrDKB2pQEKihDIqACHqi4iZZYVDIOBGpK2QLLSFRl2dbbh421FQEVhWxWHhUCKo4cQUdnNxJtDqiQGXgWHW1JbG+uYWl5Ef0DA9g3NKTqfybpdb+uOpsVCXx+0hNnwp3yRSnT0p6dmdFzpfTTBuWFdnIY6OmXbwRZJWS7MAjZWltT1XxnWxtOniJQMYHh/WMCKkg8bmtNyVxUHiIMrpwWewXIcUAFq45VreGAivPnzilhwZ9zLNBsilUODOZK+QLWnPRTf38fPFDR2dVl7AtHm2dQuLNjz5PSR2b0WsTc3G0szN82o29KTURZPZGrSD/RnJjSTyFE8du/8xUBFRmN2YgqjxlzrK2vKXnG8dze2qbEz8baOja3WIlLhoTJtdDQmCwJ6rRbAGqJMqs8LihRyQ+TYonWJFZXVlVhysqWixcv4dix45iamsJOnoZhJXR3dqKnpwvJRIv61jTSQ6Ypni/g2WefxcmpE/jsZz7jtOQ3MTN7S8AfTX7ZD8lEu95jelSk0yt46qmn1CaBhE5HXoFexICKa9euVjwq2Kc0maVHBccTn9Nrr76Kp5/6NQEVnDOK3FhwrsgXxGwYHRrGyRMn3OaijFIkjG999zuYOnYUJw4dkZF5MUJpnAhefulVdHd3YmCwV2sAg7Qb07PyvDlxYqoCVJBRQXkrb8TmgQoyKrz0k8y09+27I1Ah1RP38TNucE26U/AnhVO3cQlu9BoBFbamuYuVTAO20bHlkJmq+e/zuTDR66noHqjwYIUHQZhYLpULqrin8W+oFEcxR8+Pv0FPdwyTxw7g4/ffw4VPLmBleRnrmxkg3ILB4UEMDSfR3tmOSLQFiWQ79g2NYnBwBMlUB8qFFrzx5kuIRMs4dfIs3vnZe1hYmMPxE+No70givbaGG9dvoKOtA4cPHsaVS5dx4cJFnDg9ifHxo+jtGsPXv/F1PPTgUczevq7E9Y2b0+jt78ev//pvIJnsREu8HYlUByKhGM6f+wAfvPcShghSjB3E0YnT+O5//xvMz13FH/3RVxBJDstwvBSKIxJqQWZjFc8+8/9i4lA7Jh96CDdvbmDmxjr6egfR1k6wkGMoZH4yAFqSbZLL21hfx872Jm5ev4yN9WkcOz6OROsg3n3/Kj746CK2qY8fC2PyyBQO7R/F9PS7mJgYwomTD2F+qYT1nTDa2ruRbEnJ/0WbHQcECKgg0yVcQp7ST0m+WwTiStiiCfqKeVRw7DKRKwDcsSD4Pne0phoAFawKIzW+IONnGrDTWHppeUFsmYmJ/fIJsiqrmAMq8qqcY3U/f86EgmdU+Kq9WqBiVbJzYmwV4YCKMgyoMK+GWqCC0k/GqOA86IGKeo8Kypd5eSOOV2PuhQTMC6ggoyJDryD6FsTFDJIsAtkeyZSS/h6oWCWjQt4WtrH2QIV/n2zzHsb62rrm1KBHhSTrHFAh00R6hnBto8Sh8wnhz9hG3g+Pb21NabPP5AdjEfabJc9N1pEMBFVaU17JMyriBO1iSt7QKJznI+Dhqx6VQOG1t9Yray7bSY8KAhVMXmysb2oea2tPqU8YS1SBihKyhazMymmmzZhB3hasrHPVotzYSmpSRFLzduCzKsgHLABUMN9TELzv/HFs4+uBCs+o8AC2nysFVDhdZu9R4YEKGoCb1FVZ/euBCj0jJk8KZgpJZhBrcQm2CaSimXqsClRsZTadWboldqIxKyhhHCg5tb8HRkXz3UzjjDRNOff2+ftPJzQrvGqWX22UP7e7dXupRk1udrKGnaEqnb11U1jpqD0dUy+bcXdD7mbgyT08owZ7pl2Ntezo3u6h0T03ybOrCXe4yYaPTT/c2337iuZ7v5EmDW7aH+77dwV9gnfUrF8ddSjY73d7BrblrXw8m6EpoNO0IwIMCX/OiqxLk4PuMDx8TsSrXdhY8oLNliSpSAo3OI+aUO/PFmhGs3kiWFjj18NGrbfjrVLfx6tKmnpgwhXkaMS5NU9tll9BSBX6JkFEdQUveRpM91dWGyuR9x93r6rWl9RO9fr2FfYL99uOfRJgsVT8Byq+DcZ8EFPDfY97VK7HvBOBB+7vnvXAddWYAFaO5AERxfdurFnuxJ6RT6Kzr3yBA6/HKZHrns4fYFRw7eb+i56CPIZrL3MgKhJzUlU2O1uuSJdR0rugCnvuce1azKcYM83228aM9OoR7Hd5HThfB8vL2L6OOQ3PKgkmx2kqbbEuZaz8tVhTWTS2ABPvAjnIJIg6uWcr//I+Gdq7uOcWIXtXIIXFBPzdf/iPVaDi3/5bxu4ZM7l2vB2em/G1JL+Z9LekpBmuO2YGzxcqG+gloIj9w+tIysvUCUqsXPJjlaCZ2A4cM7V7M8UsZTJNzLzaH2OAj8VyPldmxW1l5ORLYn2o8c/nJrNvky0VU8JJhMkUXidlzGZjwu/FPWhC6VGBLU5aSmNW74TJXt0HKu59dbr/zV+SHvjfmgAV/qWqxqDVpLzeN5WWBVgFTQIAy5XfAajwCXDfX0K8qyttECSpXuIegYpd1SgOOK9MJu6ibkG1xM/uwM2kojiZVBrpDww85WCbfPsdxc8tmMEKivo+8fdsqKhDZ2oCjiCDo7npdc2wC2be7BZ24xA1NGJ3Dw0el1sCa4GKIKOi6IGKnBL71OCXdE2WQEXATDuTwfFHn9Dky0XHDIxN91hV/qWSbUi12HIBz1tiPZuTHAXHABOQPObixYsVA+v2ri60OaCCFYnUXOcGeWc7g8sXPqlhVNwNqPCLA9vPZ8EFS1WhGfO9IEhhJkZWRc9FhkCF96iwalomqMioyGjBrQAV0pbn4lwFKmimvX/8kCQlxKhYvCWgoiUcRWZ7CzuUJkomMTszi1RPV4VRUciRUXHEMSqOoLOrpw6ooKF4i6SiqH/ev28QA4MDkj7xepa+woCJe89qYWLGMyp4b/VART6brwAVZBWwb8h02CRQIUYFgYrTAiqGxghUrMu8ldJPCadZmdnJOkaFJc4ITDAg4oeMCv6bEl2ra2lcunhR8jgtNB8r5MEAiQkcBo5km8hM+/vPyn/jyS88iZGxMUnbKGBzBm88jh4VvB8yKkSzLZZwe34BC7cXRFpOkY1CKiyKaGkJIxYr4+b0NbzwkxclS/K7X/lDjAyPy6icpsSJFCVxSjJ0Z5KIEhVdHZ3qOzIaGEwwwcREKE3lbToKYWRkWMmvWJTBihnnmpZnUQENPT+6ejuU+F1cWBJr57333sfB8UM4+8ADYlzw3mgAvLh4W34mk8ePYf/YfrFQsqy6LgPf+c53sH90DJ96+GGBI3yXbt26gdXVNY1fSrt0tPeIXUFGxcrKMp5++tdqgAoFVgps4zh//lzFTNszKiRxVrbNxccffYQ3X38DX376aewbHBRbKZFKgiwrSs68/tprag+BCmmbKyqO4K9/8AyOHDqIqUNHEOamIRpGoRzCKz99Fd09XRgY6K1Uk0xfnxGj4tQpAzt4HnpUNAMqmBx784038PCnPiWAM1aZ66szpTY4vM86oEL6to45V90WNl7Y7dG6zUkN+L6bUVEJ9tmWIGOuLtFQXx/JcUKggsCWBbduLnFV2ZVAm4nxUgHFkD2bUsEAvY31Ofzkx9/CialRpOIEAi5g//4J9A4cwCdXbuGDDz5CZpOgXQIDg32S3eLegYAcGRfdPQcwfeOqxujJEw9jJ1PGa6+/hvT6PE6fHFcC9Nq1G+js7MX+0YNIJTrw0xdewkr6Jh5+6GEcGJvEf/5//gtOnDyAa9MXEYpENB+9/c7bGBoew5e++JTYHPGWFNLpdbzy0vPo6Yzg+OQpDO+bRDLej+98+1u4Pv0u/pev/gHC8TEUyxHkiiGsr21jce4m3n7jhzh6pBuTD59BLpvEres0Ie6SETE3FtxMSFKQ7KlEK7huUBoos7mOW9NXsLk5i9OnJzG/kMH3fvBTtCQ6ceaBUzgxeQQtsTYx+N5793kcOzqMqckHsbRaQnq7jI7OHiToMdBG5oZtWvJZkw1UNVwkb8yJJAGEMnKlojwqKP3ELa4o4pmMYzQY/Z3jpLOtHqgwJhxZD9wUt7a1oZAvCqhYWJxHZiuNicMH0NHeqqQ6K+zIROC1+SHgy7WH82IQqOD1feKXIAjnNAIVtimG5iu+b2sbWxWggms2jzFGRWOgosqoyMgQmfJl9I/hK2KbYM77BlRwSli6vSqgwjMqCPazWkzV82Q/RONiSXpGBRPanjVQD1QIQKgDKuRR0YRR4YEKfico9cj7E0uks9OMyItlxSK8rsy1KXuga9UCFfKoCAAVszMLimlk4O31jJXkD4F+NTwHE+9ch6dvTKMjAFRInrA9KXYe+5zyAZEwmZMlbGe3BVSwKIP9w8S9B0/8HGkGw6wYDImVoQKDEmM206kWm4KhbwCoCDIqvEeFT2zoGPfx1bBKAjCGLgK3bs4I8GhrbxPAQ6BCjArGPa6qUYwKl5ghUEFGKZkq/DkZFUy0cM3n2KL0E+c9z6ggUMF75FiilKKSO9utv1iPirtnt2sXg7slQXctHU3kXu6YpN1jsrvJ13+hQMVe97pypt3Dfag/GifUm3d5bSfe/XKN5KUaFvbvvtt73o7u4Z4tpWjXChxmiV/78a5hoptsco1mHdW0SY1/oWTo3TszGFzt6q9Kvrxhm9w93OkdCBxXyUU02on7eEzfd0V4/Ps9vqeV+Eu3vDegzLR6KsRXl0m2Kvamnzv9KlDhb/Gq+Wb4KmobJ9Xz3+kR1cSV7po6Y4AJYd1UHU/+d571wLWheisuyRtI9Cpvw3yDO0VNO323OFNk0+svi6FIHyoe6qv6/X1V+4xoerWjKn9z986ktL0cbi1SP1HNwJLC3s/KwACL173Pmx1m48R7QlTXKDM89gn4WgDHecg4pYT6F9Pfi12Tl7TCAc+k9owLYyXYnsOzE3xsIYlG11afn5AngZgn9NAgY8LAi+CkwZ9X1+rqd1KpVue9aTIbbA+ZBUzeM8EvdgmLQlzcqP248j3GAFXuj7Oyk4KSn0Y2a+oFrg2cK1RMqLbzu+Znyj7geaxIhWCI88t0AAbBB8WdAP7vgJn2v/nXJm0rUKJYUBzB2NoXpviEvW8j43xKSqr/Xd/xeB9/0MeCEqoCB5zfocV0CY1QHk//Ez/mxX7leJIXmQEsJh1mck+eseEZL1boV0KIsbr89sj8MDCM+34pa6jyt8qM99M3VRL4jPgl3mMFiHFMersGwZZqm+QZyXjqPqNirxHJ/e//j94DdwMq3JwfuA1Wnu8GKrQQNbhZl5ur/U2w0t9RCRql+f0JK1WtlVXpniNDd93q97VQ+AU1WNl6lwfllRdrwQqPnzYKG6uL6W6AY/f3LVCoBkOWzHIVB55uUWmvYzY0DOZsMdSnHqgQJ7N6o9avwZM0ACp8IOO/xknVPf9a6SfvUUGgIit5HAEVDrCoeFRkMjj26ceVZGElvvwQSNGjZrakcqy6lDREae9x8WRyIJfH8oqZOo4MD0s6aH5+HhMTh+WVQMmjjs4u6QIyKbO1YTIavMbF8x8jvbyE3p4+9PT3aUNMRgWln3j9TiVCq6ZLpCLyWdA4lAs0gRZvasUkN1FrgStFY1QYUBFHV2e3FlgGS9TRpvQSGRvVylHqQTr9eiYonPQTaZEEKliZvr25jqXFm2bCGY5gfS2N1cVFjAwOYm5uDsnuTqylV3H+gw+UpCdQkWxtq0o/UZ86Th1ya0MyEUN6ZUkBBc3E+/oH1MdMBjmmpBZOSiExUU4AIZNhkj2kyk+OpdnZOVVetrZ3iB1BM+w+x6iIt0SdUWnOpJ/EqGjFqdNnMDI+gWFKP21sCKhgla8SUgWTAzHpJw9UWKKMHyafJL8VDiG9to5rV66orezjPBk2RQIVNBU1oGJjlUDFD0FGxRO/+nkBFZ1dVaDCvFQKSuZwGLPq2SiyJSwtr2gcZTMZyUXxWUbDvBbQkgjj1o1r+MmPngdKEfz+H/4TDI+MG/00GkKqLaEqVSYJqeFOHXHKXlE/ncmt7i4zaTft+GXJ3HCMHz92TIkvJpMVaIbNp4NJr5aEJd66+jt0jpWVVTEyXn3lVYyMjuHTjzwq6Ss+GMpI0eicTIihwX144OwZVR93dnfp/v7yL/4S+wYGMDV1Qka/kWgI6dUl7OzkVGXMhFtbayc6urrxyfnzWEuv4Omnn1aii+8eg1YlNWWAGqsBKvqc9JP07stmOvfxBx/iDQdUELTjxoMV35l8Vuck22J8dEwSVqzo1sYqEsZ3f/gDHHVABTeEBCryJeDln76Kvt7uAFBRxvT0DNbXN3H69EknB1XCW2+9hVOnTiGhvqP0Ez0q2jA0PCTwqAJUDAxKUm7X6lEHVFRmRQdUVKpXmiQBVOWmkwbXA4fl1xlWWlLPEqgyqCM1nfYU7thauYeqVh+P4xjp7mbSnYbLpHNbsGobH1dNxriXFVplMqYIVHCjEkYus4Ppq5/guee/g3gsgy9/6QtoE3MmgmTnIFpa+7C5kcf1y1fx8YfvY3l5Hgjn0dGeQE93K1LJOKKJdkRikFH9oYMnkIj3aB7+8U++h52tBUwdPyKAiSbVw0MH0ds9hMsXr+JHz/0VJsZH8dlPP4E3f/YmwpEczp1/HwODQzhw8BAuX53G3Nw8xkbH8eSvfB7J1iQ+/PADpFcWcGryMMb2T6GtdRyxcDee+/H38f77z+Br/+IPUAoTqIhhK5PHjekZXDj3Pm5eexcnpoZx9tFTaEkMYuYG57IUWNlN8JiU+GxmW4yGlmQC4WgcqytrWF1awuyt62hrLeHkmVNYWilgcSWPwX2j8ntgNftONiSvn4/eew4np8Zw5PBpLK+FsbqRR1dPj8BlyiWFIwQdDajgu0Z2XSlc0KaP8nV8vwmUcE1cXF7SnEMmF8FOguBc/zgfs8JQTCl6VFD6aW1TXkEyRY6aeV5bGz1uclheXMDt27PI7mzi8JFxtLe1SWKKcyYTvNpwEjCPRDUX88O1j2CBVezFDKiQLF4E6fSqzm0bTQ9UAGsbljDmf2JUEKjIZO5B+ikjhllnZ4eSywILJB1APWGyIRyjYoGgr3kJUfqpwEIFbZ4JVBDojksGktVoqyvLFSkrvvec87zkEdcvvh+Uj+C8zPvk9bj5E4OT3hfyqDDPB75/8qLI2VzF43xsJJbh9rbWB95zIVcUYGVMSWMueEaFPKKd9JOACu9REaJHhZlpEyjgdbXxdfHVyuqy5gQCXZRzun7tKtpSbRqjBNLoVUSggr4dAncEVJBxUsbWzpaSBCzKoFwS5cW4trLyTvO3vGssOcxEvySVEnFknBQBh4M8KiQDTpNMbn5NaoL3dnthQffNZ+eBCkuIVILCSqWiBdch3Lx5SxUz8i8AACAASURBVJWUHR0EKoxRQaDCkhzVZIGXPmhJUu6RZtpL2vxzfEm2LE6gYh0bm2sVoEJFDQT5oxG1yYCKMLCV+gUCFU2Mru+0T7jHBGj1FM116RtupiyltKctZbMm/UKBir3ed0XeZw+3omOq4832Rr4/7rQPs2vcObfuE7IN+rZZ3t8zHaubVLvQnR5Pk35qfshuk+XmQIU7S0Nzgp8nOf6LAyqUrw+cTk/RxVy7R4B7Fs2AiiZJ6uB5KocqkxoYI36Y3BPoEEjny6Nib+9dBagIhIWNiiBr7v9OY83/rjLULUFpL0E16e6BkLthSfVgRSOggvtENd/tWTm4vXdCLeBSBSo8WKJ4NqBOre97tMODLlosTZWB6yj3hH598clwe6fqOkbxiz3lCqfEARXWG9VX0dYw+iuYnJDfY/pr1UftFkdbxbsH4Fko6fvA1B+skp5xE5PW9Hfzob9f34LP1WJ0M1jm941RwCIBk3YVpMLzKHltiW8PBDGuYJtVxOnMo/09+OS6Z2b4vYA9tKr/k9Z/STlZboL93Zpq035YUkT0AhE7gPEBQQ9o7+ZljTxowpPy/nkdL+PkxwHjwK3tjMVDDnComJWLoRDVs+J+ke33ShqxWIsK86zJJuPF/TrXfsapf/ofqoyKr311W3GxgS+2j/KFrtofUYVB+1UW8lCW2yRCzZPDZJW8nwPPL8CnbF6kZB774g4+Kw9o8RUw0Io5BIuhrADS5KbUdzRUdICQmBF5Y0kw/uODL4Xd9b3RuopwrQ+91yDv3zxFzKrQy0p530EWVtrzZ6GVmXnzuVdGuhQHzPD7PlCxe1W5/5Nf8h6oeFTU34fbUPhpv8KY4wzodRudQVAgFNjVG3cFKiqBni0vtame6qrDhE4g9V93nWZBRHB1t0N+fqCimtS3nJRbDit7jdrIihuz+o+vpLV1tz4SY+BhG9cK2t8AqLBL+0W6UTR3B6DCdpHVtrset9PVgxa+9bb0V5pcA1TY5M3J05tps9qbySADKDINgYrjn33SZKJ2dpS4ZWKayWv+W1Wa1GCmoTUXrUIBxWxO8hjp1dvSuh4cHMTK6rqSNidOnFYyl1V7lCYIh1kFkMfm5hba21uRy2XwybmPsLK0hL7eXvT1D3JF0GJ4+swDWnDa+5lQZpLcNuZM7vD3GxubkjwiUKHkUdSqJ00/3KiSTBL5qocuJ9thuohWvUGwhtIcZFQQqa8AFVz0wiHsMOkdi2J47ABCUVbib2Jx/pZMUBPhKJaXFrGysIhDB/bj1s0baOvrRHo1jQsfnUN+J29ARaoVBw8fQntPr/qOyRgGAgw0ufhurK8h1sKfJzHQv0+BClkvpMc7pqQzZWZCKquAEeEikkkautLIeUHPmdchcMJFtLu7RywNVvbmaC5eyGM9ncbrr7yC9taUKv+Hxg9ieGTUTJ4BdLRXzTgJOLAPTVrE9CS9vjilRRSwlkrY3NjGtatXVflpRp40WqU/BJMfEY2PzPoqfvC974LJ8yd/9QsYPbAfHV2dtrC7IJeJ9Ex2R5WjXR0dCkz4s5X0KmbmZrCRXsPgviGNgSg102NAW3sLbk1fw/f/+hnEIi34vd//I+w/MIFMNodoPIJEq2lmLy6YIffqygr6enqUvGNyqburS888vZ7G+uYmLl+8hIXZOTz5+BPyUckXDeTy1RE+4KSXx8C+fiUXOY45Dl984SW177HPPqZgqRwuYyuzrYQQjV2pPT959KgCzMNHjogV8c1vfhMD/QMCKcbHx9HZ1YpsdhvRcBRb65vSoS+WzeR7+vp1ZDY38eWnv6xjvca+ycRI0B/nzp3D9PR1ST/193QryKX8GRPT+UIRly5cwMsvv4ynvvglgYkM7pLJFuRQQraYx1uvvYGJkf04fvw4CrwHh6U+88Mf4NihCZw4dFTTUy5KT9cQXn/lNQz09mBosF/vE71cpm/OYWl5GWdPn6ok6AlU0ExbElrFIq5ep0dFG4aHhgRYkslBnw5KszFRG/zUbrhqZ2yfqOMzqmwAG2R4rAorMBe7MWeVYiXp4TPR6SV2Uq2UCDLTZUozBef02kxHdcvlE40cG/SpIHAkoEObMKOfc2xrXmIwq95lhVQemxuruPDJx3jnrZ8hvWZ+LEcnRnD6xBEU2bZsCT0D+9Ha2o9wlGa+BdyauYWLFz/BzM1p7GyuIh4PoWegHa3tYbS3t6C9tQd93aPoaOtGOr2EhYVZXLjwCY5NHUFXbw+6Ovehu2sU09fmcfPmR7h08X1MHj+CsbERzM/N4I3XX8PRo5MYHN6PmbkVdHV044OPPsbw8ACe+PyjyBc2sbWxgYnxSXR07Uex2I1QqQ3PP/fX+Pij7+GrX/ufUQjvR64Qw+raFqavXcNrL/8tlhav4/TJCTz2+El0do9icYmAcwiJZCsKBWrkbyNSYia5gHw5g9W1bVy/PIsb124A5SwmJvpx8uyDCCWHkS+0CpQlUyTV0YXtHLCyeAvn33kGD5wcx8TEg1haj2N5NQNKGkViEbS3kS1gNHMyHTjPSgYK3BBRNrBDcwzfU86zy2QJilER0xzSxiR5NCIGEgHPRMrYM7lsCWvrmwLeKTdHjxyOCZN+ymJxfg6LC/MoZndw5Ohh+zlBUGeuaKaQtlG3sUwQhWwPSgSaFADXN4IT8QiQXltFqjWh9YRg1+YWZRnJEFuXLw8r/3k8+4aJfFa9k2HGOdtLPzGBzH5ggpqbRkopkpXA9zQ47xtQEaG6IZaX1uRR4YEKk1C0za034ebmlHMmZcuS0RYlxDlPmd+Fl2HiBt8o9bx+ZpugDIEKguVx5AhUhKkL3WLG5aGwSfXtZNV3lSo9hOQzRaCgq7tLG8lirijwmTEMweWg1BQZdgK7Y2ZizmuJARGJ4NaNea3JsXgYrW0sAmD1IRMKJaymV2VwTRCHMQnXPAHX8RZsba0rNmLSn+sJz+XXSnptbap/d7Rp5zFk0PC5a7PPxIQq+1h5aBtrgkIM90qhCEIFyvLZxpnjg4BaKVSsSMVzrHgz7fZ2glj0x7EqVHLFGEPw3JQxZJ5FmuOI4OatW9qkkxUiaSZnsl5hdjhWhZeRMoZkHIuLSw5AMlNPVtiuptPYWidQwfXW5EGiUUpYxQVUsE+MUdF2H6io3xk12Rr9UgEV2mPVpyB37RRr77xua/T3BVT4i9b6nDTNODfMFjRNgTdIqDcFKir79T1U/uvCe0vA/1yMirpL/NxARUOQokEiu2Z37cAeZ07skhd3yNoEAYrqHrgZUNGs90LOW8FlHfTH3wWosELQQEKcC5FjNQTZAc2ACsNs6hP+9l55OSmPI1hbrb0+IcrzGrC+CzFxKguBcwe+IvaMl9JxRtGKPqiz7+JmLyHpGZoVVkAlx1Lf7upcYKwjF597jX49awMm/HX8PlCV7E7G2cf30vt3e0VLaFsyWrLblDZiYphJYXcfBBgiSl67e2OFfSBd4hPIFSaDm6rUh96Tw/Ul4wTGAfSjYA5FuQenMMD74rV0D7qGMSJsv2j37dkJHlTxskb8eZ6J8FDEmFllVNgN8ttKpJy5tMkcGZ3SMUPcvSiGVVLc8kPGZnCG4s7oW+wCQgzhMDLblGVq0XVtb+MYBw4g4t6M8Yjt441FQUkrPn9+GIP5PbuYCqUS/jQg/fRv/jW9SUxiSqAOQjpPxctEPhwGEogRUeRzsliJBSjsW6IABJ7sfXLeEUUzZ7dxbzkt38+MZXj+yriXcTolj+kTwSIbSk6Z74Tt76iIwBwFiy2oUkEJXhuHjOVMGoxsYgOGeJxn7WufKWkuK9ZlfG3f4X7CS4OZubv5hFSBCh7He1csep9RcYf5/f6vfil74I5ARSUKC0zELtOvF90BFbvhgJp5u0EoVD1fvf+FhU6eneG+p4k+GHnWJ+j3BlTsPTwz3DsYdGjqron2G7WpvmfudA8GVBiQwKpfq5KwCbLZcQ3dsY2aphm/tk1eM6+m7QFfCl8tERzI1bCtev+6K6LUrkqhHqgwRsWOKi0peUPAIsioOPqomWlLFiPLqv+Ekp5MBsjAiIyFeNy0vSn/xMoDAhXp29jcXFeyY2l5DYlkChOHj2ojS1khJsKZvM7lLFlC3wHK/Xxy/kOsLi07oGIAlFpim0+cOqPFprW3qzLpc6L3VR1kAqysrimJxCSJFbIzic0EPqmB5rXAYcCFkx4EVWkEyj8VDagoMvnNivlkBajQyhMiUJFHuCWO4dH9ogjS2HXJARXxUATzszPIbm1j/8gIZm7dQGtfB9Irq7jw0Xlpnk9MUPqpDYcOH5J/BStPmWg2yREzWCKQQKkHSrgQqODPWOkbDEyZvCgWQgIqmNgJhQlMmP72/Pyi+ovGres0Js3nxBZggkpa6bmcEqIb6TReefllGcCeOXsWI4cmMDQ8Ivkj9huTW17yglUUDACM7mpm4746lckj6UvSZHRjG9PT0/JpkI5mjpWwZDswmRSR38XOxhq+/zffQX9/L574whcwduCAGBU+IOYYZiKdycFysYRuJ8/E8bW6nsbM3Jx8LujfwU8sysQh0NoWx42rl/CD7/0QiXgKv/O7v4/xg0eQ2ckh2hJBsi2hys7FhQWBCTR37e/p0T2RscDxwOrZlXRaoNT87Cz+6s//An/81a8hFg6b14RLHuqVohwamRg93ejt69Y4Y3UGGQTPPfcTye888cSTVk0dKgskmJufF9OGFfP0YGBQffL0KfUlgYpDBw9JXqevrxfDo/sQDpcRJRU6FBZ7ZnV9Azu5LKavXQfyRTEqyKTRO+3MXiWfFYng/PnzuDE9jccf/xz6uruUIKQsSz1QQTNtD1S0xGMohMvIlgr42auv4/DoAUxOTiJXLsrQnrPe95/9ASYPH8PxA4cCQEVYQMW+/l4M7zMWEIGKG7fmMXd7HmdPVYEKSj95oIJJvus3pvUOjAwNayy//uprMtOWv4MLSCv7inuolAvO81Wwubrm1K4DteuCbST4DFnVnVMikXOJN+atFgLsBp2rm0LHtgtBwA8N1Jkg5lwnCShWAOWLMrJV9VA5R4s46fvP3LyBD99/BzduXFMV99FjUxge2Y/rV86jJVbE4YNjkj+LxNrQ3TWI9u4BxAgCckNAIG95CbM3r+P61cuYW5zGTnYJ3d0p9PUMCKRgYl2gXqoD8/OzmL09i8GhfThy5AQG+8dx/docEqk4bt26jrfeehNnT59Eb2+XzLz3j42iHGaifxsPPvAglpeX8Dd/8y1MTk7g85//jJL1XV1DSKYGkct3IIw2/OCZv8K5j3+Af/HHv4didAzZbAjzC8u4QJDsxedQLGxg8ugBPPHECewbPoT5xTzSaYLf3BBtIhTKSh5n+/9j783f5LzO68BTe3VX7zuWXrA1FpIgwF0LJUqWRdnOasVJnMw888PMM06k2JKT/yHJT7MkM5l5nnkmsew4j+OMEzu2LJMiKe4SN5Aise9Ao9Hofauurr3mOee996uvqqtAQNF4pBmUBKJRXfUt997v3ve+5z3n5Ddw6doFXL9xB+VCAn3d/UgnI+gfiOPY8ROoJnehXOmSgTifpY5uB1Qs3MS5D7+Lxx/Zj30HTmBxPYWVtbyeL85PPWRUEAiv1gSuah4ulcltEVBKlp9VpJU1fy6vLKOKqNgAnEOsPc1XgpvhdBfl5aIoFEpiVBhQQUo9s8Jkh/XKC2nhzm0s3rmNWqWM6emDAqU57xH0oIyOque4YVRlm8VTTMrzGv3GL5VIyysglYyKXUWZIbL9uHXfyhYQjcSxmdvSuTl+uSHjeOZay/GdlrxWRc9cfx8lyjiPGFBBkIZABaWfbOxb4sPYk1xTmbSPYGVpQ+BsAFRUyfgwINv7+fgqOgIV6VhyB1DhZZgIVPDxZjvntvJiVbCSkGtLsZxHLRICKpxMHxMGBBK99BObivdHsKK3p9far1STR4XYoK5owSd0IlHb7PN6BVQ4g2+OidkZmlKXkOpIBEUAnD4JVKysrYilJ6CiWsX169fMp0Mb1pyAbYKUTMozucENsuadaFSMu63tLd0n29YDFbwHJgakXa4qUYtTuNYz7OO4E1BRdDre9KaIllFBBbQFUAVipSJgmOO1qztjm30HVEQicdSq3Fxz082NO5NDBmpT+onJOq75BGU5RxmjgkFUSH7ByUTQNJxjjUAFX7wP3j83+wTUt7ObBijpHlityPtICHRlXPWXClTcw5pxb5vB/68wKu4jOa7Nx/0lx1UY17ZB2yExjV/4fwSoaNqa7fRYvLdraF8sEYoxGjdljRts/cszgO6jL/4ygArOPQH75F5wEV5UGzZTMwvDP4ctnkfLDTcxDupB311Gk2vzhmHVnlFx70DFp8g+3SUpoUr5EIPH35dn0gqA9kx9sT/qtxeOKgNPBncs32xmML1T+skfxfs1eHa1BzBaxdDKWXivBPcBVbtzLXLGzHw77K9g4LY945rHQwVmNrRbgCDBsYOrCG7ax+MeWPFt55PfvB6uLR4Q8UCPPu/9nFzuhTEd2bFKCntPjaYCUrVHMN4s+W0MDpZbGbikeEem2lahX5cMsuP6e2SuwBLOtr7z1skO4F7MVB/qBuLh6xbA4uSsvBwTE+TsC0t0Ow8D5+Xg95ZsNMkoielRNRNr+VQQMKEqQ9nJkJp3h7E9bA2279mxmSPxpt7GwI8HDBoPRPhRHEgpce13IIgYEs6bwxfr8vhhoOIf/AaLViqKlWUq7YAiMUx5X9WKch2JlLEuCNJY/GMAm2S7JP1KTxFL9NPLw9rZvEB8+zLO4zV5qUoryKiaz4u8SAws8UAWCx+NhWKeEkYnMgNy+oqxUIfnYxEt8138mcBU0G9ikzBGM7lqxjfee83LSvF+DbTyhuC2j7AH3vpfjJgHQMW9hV8PPvXz0wL//O8cD4LAcI1K488mbaHngcmlkDGRFgUvx7gz1+JDqOBv/5G6pbO9Y+er60i6U4WS9F4cwz4dLGwB/a9dmzdGkyEiRCN7w32sfn3N7I46o6MOrjgwwd1B/Zos2PJov11Z+PqtLZmo02/0s/+8ARUeXdY6rYXfUSkDyiN/0waoCG6yNVARvKu+q4NB6t+gOsDer1dc1CMDfUWGrXV9RzEqKmUl7j1QIXCiBVBx6OnPa4JlxTgTzZy4mUAOzBZJ7SfFkrt4Lh6k0lWrWFtjQpjAQRzZzTz6h4cwvncSq+vrkhWi3AUXFNPF5sa+U5v8c2dPY225DlREVU1fxdFjDyOZTiHT3xP4rXAR4ALERZdSPawmZZWAKgScPKYlJ0g/ZPLbzLT5PQIlTNwYVdJYFQRpyKjgwu6BCtFjnQElgYpYMold4xMy4SRQQUZFiokOUHroBtKxOPp7ezB7awY9o/2tgYpDB9AzNKwkBjf5vH62MUEEPrOU0WD1P4EKPrM0lPWGg2QoeNPU7a2ikk4EKihtxETXwvySFnHqoa+vraliggbmZFQkE9ZWXPDpUfHWG28gQ6Di0UcFVFCuiP3KNvIVseaFYR4OvrLWEihMRETF/vBURwIVN2/eVJ8qwVfM61EgUMFELQ3FC1ub+NM//o8YHRkWUDExRaCiLwgUPJDGSnMCXwM9fWoDjtm1jXXcvjOH1eUljI3tVr/SOyIW4/UmcPXSBbz4vReQ6ejG3/ibv4Z9+6cla5ZIJ9Q+DCIXFhbUZgZUDGr8ENAhUMFEC4EKylgtLy7i9/7Nd/DNf/APMdjfh2wuK5ktbUTcs0RQhwlC6t0zeUM5MY7lF1/8PgYGBvGlL31Z/VhT9WpVFdmUf2K/DPT2oVgqS/KISaGXX34ZTz/1tIAKtn1nJoXOTBI9mR50JFKab/PFEuYXF3H+7FklcL/2/POqeDaKKfXYaazK5FMc5y9cwMzNG/jc5z4rRoWMzKqsGIkHjIq33nwLX/3FXxSbgd/tJKOCoEqtglM/eldAxeHpw2AqXfNINIrvvfgXOHLgEKbH9zUAFe+8/SPsGRvB+B4bs7WoMSpu3LiJR2SmbYElgYqHHnpI454B5LUb1zVW94ztEvj5Hj0qnnhCVe/3A1T4iqtmoIL/Dqql3LTYDFZoXvfze9O66DcUYRC61fcbz2EgNj1hCFQQsPDyUbUKrweI1mJKPs/NXcZGdkHJ1Yvnz2Nh4Q6m9k3g0ePHsWvPfkSTPVhZnMOp997GntEBjO8a01y8urqBWDqD4bE9SHb2IBKzSnNOfGRlETR9+4cvYW1tVn2fTmcw0N+Nvr40+rr70NWRwcLSHWxsbmBigoyDY7h9ewm9/bsxNrYXL730Ii5dvoRHjx9FV4bVTRXMzS8L6HryyScwN3sLb7/1BtaW7+Dxk4/gqaefRnfPCDq7RxCLE2TqxR//xz/AudMv4h/+xt9DsmsSuXwFFy9fxccff4xrVy9hsL8L1UoWX3r2CKb2HcNGLoqtHNQWl6+cxcrKHZRLESwuLyDVncbuXQcx1D+OTDqDO7evo1pZwUMnTqAUG0G52i02HxlS6e5ebBeB5YXruPDh9/D4owcwse84FjfSWFvPY5BABVljAkG5Ca6iWCgrmc95phKtOUZFt0YMny0mwJeWlyT5xzWN8nFM6srsOJnSxi3VlVSckN8uYWN9U2srwUZK7hE478r0CCQWUDF3W8v34emDSKcJ9NqGjKCHARU13Yvt8DxQYUwLn1znfEYEhEw+0uK5BpOFsF0oI53uQjyVUeU752omyDm/8T7ItKBMEZ+/dowK9gHBQoI1Xk/ZNpkEhwmyRbG6vCnAhtfDNatSteo3fk5J+I6OgO7P+TYVI7XfVax5Y2vne2GVduYTspXdNvlCAhWJBApNQAWPT1YI+4WASFheQYwQsWG61S8EKmj6zPeagQrioGGggr/XZyJM3pNRUUJHhiwO9nkC5VINJTI0BFRE0dPbo3jv+o1rWgtpfl4obgugpywX4xUvU6DNeCyGXKGAbHZTcz7nbppps9+VHAr0og2o4DFZsMC5l2y6dkCF1ZhSxqAkoILH8YwKk1BgpWWdUSEOXNRkGzieZaZdraE7kxHAwtiS40ISE01Aha4pTaAi1haoyHF8KQFhSRKyeshSJYuWgFgjUEH2a1JtI4NWB063Apzb79TuIv30/wOgogVsbonE5sysVS3d34b3JwIq7gfcsP2S9mMh+Zm79nVbU+nW3wqDC8F56ulK29P52KD5ELbhc9tC5w1T3wj6jVbwrR19EW6K4Ge3fwxv3EPnbcmguRtQ0aa5A9+Mpntq16WWZLfx0fozzVkH89Jp9WoAdNqAFOGv+rhaM5lnvd712a3zduofs4Zoy6hoczy7Vy9X5tLY9zJv7Gh3AxB2AhVO7lN7z08HKpTKdAydxm5ngphy3q2ACtuX+DjV8umNvhhBn/g0Cz/kgAqlLAKvCwMnxARUctxkpTxo4H8OzKSDavEWjJkG3MI/S1bMI6DcMQOs2NOeQ+6DJTMswKCi9ZHXocS8k7QywIaxGc2z7Xtca7wHgZePskS5JdmZmNaa5u6T7WimxyaZawUMPkdmv+P3CH6ofdhcjgldZxqYaoOpMpgHg6+W94ltMczlb2frdPilhHaNBtZMmlfsGik3WixZYaBYGcZ44GcotcmCQ3tE6Btlkpx27W5/74AQY1RaAYPGpO6FYEZKiXUxDVzfiSHD+MwDY24M8vy6P4KYkp4yj1LdhXtO5T9RKeN/+Vf1HNe3v21sBUk2VenPUJcA430xxhXTwslemTl7ndlBWXDtqVyRNdU8OEAZywam1vIHsfHBfmeRkS8MMa8NKgwYM8SzIXjPKsAskmlBIIUeHwYASSK8Skkm+l6y6ISS15ZLEhtDQIn7mUAewQ/nM+klyKn2wVgnv83ch0mH8f8CdzQIlZCzeI/99ACouL945MGnf/Zb4J//7ePtgwJn/hPMqG6hDTMerCDfaHH18FAzjgvEQpTHICapUxh3VJRqTq+vRPYVl9APCjIag1B9OjRXh1katgDXTVH9ChSOGfwGxioVQtFlQ6TZFHa6+64HT83ZKLdghsLO+l2EP1v/mRV+vtGCSVsruL3bAO6E5EgaO9CtzC569gt1uOld6YJ1qw8wmkeBC6T9r0nO0DX5uIBos6uMqDMqHFBRLIpNsbWdDySgAkZFfhsEKhiQKJleKKpqkMGN1zCOJeKIpxyjolxRsohOm6trC1hZWdSCmEh2Ynh0VJWbm1uUeepCd6bL0QHpwUDzy25sb2/h3NlPBFQMDw3Lo4GLV6lSwfTho5K9yQyw+t6CCv7hYsNkiZIWGSZVnCQXjB7IBIMCmGrZURitgzxQYcGcaQkyOcNkBBca0hy1iFskEUg/xZIJ7J2cUjI7u7kpU1hqcfNsc7duoYvJh1QKs7duoXukF+ura7h45rwYFQcPHEKmpwf7Dx5A9+CgFkEPVLCNGaAlU0kxLTgWRkfGdK30qPCBFNd2Bi6saM1tFZSwicSqMqClzqIHKhoYFf0DAlXS6YRkKarlipKZb73+uoCKkydPYnRiUuwGJt85RpToSXnTbjIqDATylF8GLwIsUgkknCbj5sYWZmdnxQDhiyZTHIepji4LqqizTqDiT/5I0j5fFFAxJT1xBSyuaoEBQbnCILUsoIJ9RFBtZX1NOvE05B4eGTVT7ygrSsgASeLKxXN48XsvIpPuxq/+rb8joGJzK4dEKo7Obia0LLnCe1xaWMDY8KjGBvtIshRpMipW1S9Li4v4zv/5b/Dt3/wt7JukbE1BlbkEOTwoQO1zVb46wIyJT0p5eUbFF7/4HJJpGo0xIInpvBwXlJ2i/j0Tzsl00pgEP/oRvviFL2D3nj1KKBZLeVSqRTEqjh05glSyA5E4pXPWcOr9D8DQ/atf/aqCLraPycXUDFCNxXD+/HnM3LiBz3/+cxiSObclMulLwOF8/sxZ/PDtHwrsGB0Z0T1lKF2TjCNbzOOj9z7A/t3jOEyJKsIfnMMiwF98/0UcOXAQJoRX/wAAIABJREFUh/ZOaX4pxYEyonjvR+9ianwP9k2OG2QajeHa9VlcvHQJDx09ovPz5RkVHPfs56vXr0nChmAJgYpT772n8TgyMrIDqGi3QjdsikMfClcxNX83DED4n8OfuVuiLFiDQguTVfr4jaHVI/GZMZ8KD1TEEQWrb1hJFxWT5913XsLNmfPSfk0m0zhwYB8OHzmC4eFR1CIplGqWBL8zexPvvv06Hjl6CPvGdyFf2MY8q5cLFQyNjaOzq79erUzJm0IUr73xIjo6oIQtfU1mZi6hWssKSN01ugt9fdSJp3ReFQMDQ0jEO9A3NCl2Qy67jX//7/8Aa2vLGB7mnFuU38reveNKOF66eBFdnWkM9vXijddexVPPPIOTjz2Jjkw/Ort3IRXvxX/+T3+E0z9+Gf/oG/81uvv24c7SKi5epgl2Vj4avb1dePP1l/DM45OY2n8Y+XIKFy/fkkTalasXsblJ74Ux7DswjT2T49i96wBK+bgkwq5c+hiRyBIeffwEctV+ROP9KObyquAiUJHLV7E0dxWXT7+AJ0/y+w9jfi2B9a0y+nt7kZC5b68z1jOggklyVlNVYxCDiXOCAFcPVCwtSf6L8n9kS5BRwQ0NNzuMY9JdndrQlYo1rK5tqGKMsjeJVAzlUkGJYC/9tLK0INPPw4dp/E1JgaqS2pxz5YmjscUNXhmF/KZJGuWy2jwJUCmZbCOvg5s++jgQ+ZiY2I/t7SL6BkYwtvcwUikzg2bimX/z2B6oYL+zL/p6jTnBCkEv/cTzkVFBRqQqypyRsl2nARXra1sCZDxQQbaIrbmUTkwF3hhcJ9ZWV5HgKumeEc9esAQ+wWZ7fgj0Uk5K0k8dxuorVpz0U8qkn/gdzsMCV0Nm2nxf3hViNHQhnUyjWqoKnPY61/5ZV5FD3GIIz6jgmma+GTHMzS5ILlKSWmTtaYPOxAj7dlVygmS0sN+vXb+qpIZ5eWyjUiqaRweZBwIbTLOYQC/XMa4DZKzw8wQ0fMWgTygQzGFSg+tVImnSl1XKztE820k/VWqUfSqjGq0GjAqOU0o/sR0ZY+le/LwkBhfjJUo9KBVmoHYkrueNRSYE3lhAwrfpqWQSdsaoUBWkkwPhfbE4ZXHB/LQ8WMT74b1trq1qDeM9mEcYixziep48UIFcB8gKYqxTBypMCkxbhFC2thUw3G4t2PF+u5z5fSfg7yf57vcA9/+dVvfVKFV0D3feLskaJGRbHKPlpXoA6KdzHzv069XR/lpanKPNfYRlcRp2Z20vM7xL3bF5cuXh7n23iaofqr6TU1wTOkdzjr7lkGqbyGdM1YaQ0PIcxjhobBL7YLvxcd9AhWaEnY3Y0EXB5tT3Xf0b9+INoaKvVv2kvZaXfnIDw8dTbYa8zwF4uRt9zK2bLb/ik/JNvzRpnsaLCt+mHTeo0NSYbQmqBTkXuw6rNrd7qTMqLJnONLvt41jJ33R25kBipu1vt2SMRqtit8r9cNmjWNRtfEQ8AcCf30vXaq1xjAgPkiuF6vMv7ry+7xWNCCgwph9fkhpSYr8+LpWM92uOW8esmt6Ss6p8d9X5VkVvSgJBgl9ATP3lY3veuxL6Shgzoc92dFX+qhc1AEhsBsotyUzZphf927Vhi+EdtLGeJAfweNaL2CQ+D+ANtl31fqBqEb5gJaVpHl1X2JBxtLyn7IIY//PF9d3kuE2+yoMv/p5ZBGFtxqICMmzJ1ihbJb8DGXzlPo9n0lEmh2TAhclUcQ1mO0tVRabWLECw9vJjzxtmG7PF5JQsDrEciDej9n3rBzfPo0LPWg3/6/9Wl+r95jcN7PLMEv9o1hP+bGgn90XGh/qN7FOTYuV5+B5zGsrzOK8HL9/tnytjRFcCHwyeR+NCZFGqGfjiYYsp/PzpvTksrquzJawoxAAjnsMzmAMA0oOBaj8rAGYfsZ1ZvCHmcTwpxobUJ8isccOZ5yqUipKD9UDTA6DiHuKZBx/5+WqBuwIV4eA+qNIPVxr5JSe89Pjlrv7ezkCldaK+DhiYLI5/BZRa93Q2bzKCOb0FWLEDqPALuPfZcAu1X7zb9l4QCYWuKzCZckFQ6MvcfO98hdsrdLEuQqkHgd5nolU71Y/RMlSW78COcNfFRU2BU8sym8arbmWRrqO4hUYV1zV6VFRUaU9zVW6cPw2oYEJEuoyuYpUTNJOKWizjMdBc0TMqykxSVwgeLGN52Ywde3oH0D84jHSqU6wNboYJFJAlQFogkyMDA33Y2trEuTOfYG2lEahgdf2hQ4eR6uxE92BfAFR4kIILO6sTY6I0ctFhNYT5WBBwMPSaiR3qK+4EKjyjgu1AoIJVstKVbwYqimVEEnHsnZzUAkiWwvL8rMy0WTJ759Ysejo7HVAxg8xQrySWLp69YEDFwWl09/Ri6sA+ARUy8ExZ8p/JFSalCMZwgSVzgowKvpi8YRLJTEedT0I1KqBCnhKRsoAKJloWFlhRSSmozkD6idX9vNZ0KqGkFs+zub4moKKrowMnH3scIxMTmGgCKnz1AgEkS7iwmsEqbQJGBRMNBK8AbKxnlRTKZo2BQaCC10uPCi70ZOSUt7NKYFJ+5blf+ArGpybRx4p/JgQVzJmJF2M5GrNT+onXSzkSMiqW11aR29jAwOCQAjdWLBOooBb/tSsX8eJ3X0BnOoOv/9qvS/ppI7uFWDKGTDflKRJYXlpWMmVhfh67RghUxOTXYeajcQEVkrVYWBBQ8du/9S1MHziAWDKqZNetW7dkzipPky3q6DOQrYlBYXukCC5cuKgk6Gc/+zkltJgSIqDH8UWgYv7OvIy8vT4mARoCFc899xx27dolKZit7U0liVcWlzG1l14RxzA+OYXtYgGnPvgAGytr+MWvfCVgBfmqZ4GU0bikn25cv4Znv/BsIP1E+SmaaXOeOHP6tPwgfun5rwmoYCDNqmiwDTbX8eE77+HI1AGZiRdFowUqkRpe+P73jVGxd1J9XoxFUIlE8O4P38X+yfEAqGAF8PWbszh34QKOi1Fhz917770nM20mRkuVkhgXZFTsHhtTexKEOXnihPkIBFrFP9k6HYCZ3GyE1g6tAG3+XWcuhfyD3OnV103fa74y2xD6Cqya5GGYNCQgpop0bs7KFYFwV69cwXvvvIKlpVsYHRvF4OCwnt+hoRFMTu3D6K7d6MiQbRRTwd/VS+fx5msv42/9jeeRSsVQ5Thd2cDi8ib6B0cx0D+I7s6MihHKpQR+8IMXsHfPGA4eOIyNtQ2cO/shTp9/D7Oz15Db3MLw6AAm9u7G0GAfurs69czGOwikPoxdIxP46NRH+L3f/Q7Gdg1iefk2BoaHMDk5gbX1Nc0BTzz+pMDnf/v7f4BcdlMSUMeOP4pYohvdnaP43p/9Gc79+C38xm/8feRyCRkCJ51sTLGYR24zi++/+D08fmI3po88hJX1Mv7Tn7yI1dWsnoGjR45gYHA/Mt39SHak0NO7C7mNsgCMy5dOIRFbxMnHTmKj1IVYYhCFXB5pMhy6epAv1LBw6xKunHsJTz12GLsmjuHOegIbuSr6errFgqNHhZmcw4AKJv7pBRGpar7x0j58tpjgZ2V+DTFV0ysZ3kFGBYEKVuFznusQq48eFQTPOdey+i2ZoiQBGRhJVIoF+VOsLi8iFY9i/74pySmVuMaWyKyrYH1jXWwbGUPnc9jMLknCj8l786pgVaBJ5CViScnBManOefjYsYfR0dmN4ZE9yPTsRiJpzAaT/jOPCgIVbE8+k0zs93QTTOvSuumT6Lz//v7+QAKQ5+T4kOdQgj4JBlRsbmT1CIQZFTyPPBvc2iZgYW1drENLqPAY5gehY2pNsxwT50TvUdGRzuie6A/EbLz3qPBARTOjgtdBQIZ9w+S5Z1RwrufGkX3ln32TnDLWgpcyrIMnUUk/0UQz00VPBZ9U4oa5hpX1VZPU6uzQ8W7evKEMRAcB5iK9vPJK+jOh70EQxXnRiGIurtkEgng+trt5WJicgAeoeE6tsymTdWM9ngEVTHrUZFxeByos6vZABa/J5pyYqvg483LvT6CC9ySiDqWjdNX0qJiVrxivmQCPST9ldT1eusASSTb/0ZcqlkhiYcHLTHYKyGG/cw4nUMG+J/ikeS9OECdhrMUOY1TUttJIJUw2kgCdMSo4HngnjXHxzwRQES6Musfl6G7p8Xs8hI3XdmXr7Q7y0wIqgn3UTwGosI1Imyu+P5YHU5D3BBI0nK31udu9Wy/wCx3EqxG0uIv7xr1U/NEEVAQX02onF24+98FP6ZZWQEX4OneAHlIK2JmwD263+XzqBP9mvXDQd3VLjKatObZrDJ9d9oe+G7MhKLh01d3Bv9s0jFc7aBoXnwpUtLjvYAw2/c4KLa3a3bLABBkMaODLNPSlHdv6WXD3K8jI+Tjwg6rO9zken1txR1AS/i4Tik8d+GvQ50PtWgcqDFCxBLz1ZxhE8XJMvIE6WEEpwVCeRbJENioY4wrccEnduhyTgS+BjJJPqrtiCH8rOwuQrC19tlkJbMcekB8SQQx3DL7v208xuwNebDbdOTI96OV9KSQV5NgIvq3CabV2xVEm68NrMQNvz6pQVb4D+y2Bb6C8vKbIsGa7BcVO9abxhTI+4c81XvtyxwCoAxUs3ow5mSom7u2Y3FsSqGCPsOCTe2bGE8aWMbaFCuZSFg/6bhGTwxUNKBnv5LTYvsZssfsRsOD27v/yX9XNtL/xDYtlyDBgAabFETFdi+SlnP8HwTrGtmob+V8wHiPgZMwPH3PYtVWVCyDgUgdArN34h/GxB2h4b5LMDLFl1O0OC5W0l67PF7QaK4OFHGRVmFeZgRgNc2ITKKW8BuNwJ/GpPJhMtg3g8XJTBiw52TaBZ87k+wGj4n5CoQef/XlogX/2a4+0vMzwghYO6hueqWBuDrnPs0oreN+Wl7sDFRY2679u1g6WyCawohULYkeo2rxeONqk93ywzxstIHyPn9ZXVnHvPxUGHJrfCx8pvNTXvxO0pxrT3jcanbKSdoCQJ0eAsgua99QGTlAtQokdQEW9QdptcvxitrMN6iaxQaznqyxcICOgQlr1BlTkC+bbIE3qNoyKg099zml314EKos3U5/ceFR6o4Ga3Qn+CahX57XUsrSyqgn/v+D5tbJn8z21zE98h82IC31wcKG1E80kCFRfOndkBVHAhPHDoMBKpFHqG+x311aoveQ00xmaSiQlaAhWGqBsdsh1QQbCEm2mrtDA9x+08pZ9YoW9SD6xQUPfyeDTTJlCRjGPP+LjMT7e3clhZvI0kF9vtPJbm72CgpxfJWAy3Z2fQNdwXAipKOHSoDlT0UNrGJXS4cDOBxMVXUhtVA1RaARVWMM+sDvugKOmWarUoCSJu+hfmmTyoyaNC0k+lEgYGB7HNCk7qL8ow3Dwq3iRQ0dmJJx4nUDGF8YkJmZRycWaSTtqYHCf5nNrSAxceqOBYJ6PCBzlkVDCZt+UMViX9RKAi2anFnO1Yyefwx3/0hxgZGcYXCVRMTqCXHgpOToljlwAUw3ICFX3dlEspyzdlfXMdi8vLqBaL6OmlJBTZDKxMgRgVN69fxgt/9hfoSHXh67/2dwVUZHPbiCai6OzqUCJlZXlNiaI7t+ewa3RE/cwkWl8fzcNjkvWIxGIBUPGPv/VtTB88IPNdtoXXO/dVugzGybaYmtqn8cjEHbUtmXyfnj6sBBtzTNTiJFAxMzOD61evaczwBjgGyaJ544038NnPfAaDQ0Nm+hqvYXNjFTM3ZlDcLmBkZAxfff5rShafOvUBVuaX8Atf/rL6isk9X2HT1dMj5sW5c2dx/epVfMGZaXNmIVBRrllgeeaT02JU/PLXvmZ+GQQq0klUosBKdgPvv/0OHj4wjSNHDqMUqalihumyF18yoOIwpZ94TJlpR0Hpp30T45ia2KN+KVVq8qg4d+E8Th5/JJA2ISBDjwoBFeUybszcULJu1+io5HQ+PHUKj508KdkZq/f5yV5hQMFvKlqBE42/49pom7TwJsdfASul/HrQKnnmk4x1sKKmhHtf36BJwFCmLALkC1s4f/YTnPrgfWQ3VnDwwDhOPPY4bt6cxdmzF7G6uimW0ujoEPbvH8f45EH09Y9qE/LBu2/iwpkP8df/+vOIdXYimc5geWUTly5exdDAEMaGhwQCs06P8k3j4+M4dvhRRJHC+toSzl86JW+G9z94DwuL87h65Rw60nFMTezC5OQe9A31IRpLIpMeQLkYwVtvvI3c1iqm9u9FfjtrOrIAjj/2GKYPP4yBgT348+++gg9P/Qil0iKe/+Xncejoo8hvRfDyCy9h5son+M1v/ndIJPqxtrmF67M3cfrsWayvb2B4cEQJ++mDvQI4cvk4Xn39Q0xOHMLw8JiS2YUi9WxhIHXXEHJblFWax+XL7yKd2MCJk09go5BBNDGAwlZe0kmprm4DKmYu4ur5l/DMk0cxuucI5tYT2MzX0M+5LUozbfokWeKAkj4CAwpFSZ9tbecCjwo+W5yf+cyzAj0MVJgJcwIxPstpo64TQOZcqDRw3OanSmUL8WgJ+e0trW9bmxso5rck/1Sg7OL2thgY3q+I86UVFlRQqll1ViFPoIKARVlSUolkGvEYZeI60N2TQd/AgOaJgcFR7Nkzie0SzaBTStpzjhDlPp/H5gaBiqTWUQIq3V29SlATpCNQQb8ntgWN4FU97zasXBcFPCcIvABrq1lkN3mf7YEKz8Qgay0dT1plYUugwp51xgL8Q2o+TSS5RjYDFVwnvY8Mr9u8POyZFSsmn1fhAscPpZ/Yb2zLMFDhGRUtgQrKOM7MScKhu5cm42a8SBYj231tc13Pclc3wZ2qgApWJ1IWk0y47S22aTdoOu0ZIPLDErhUVgFBNueknzozgXRVXT5OaR6tV6l0wpiGzqOCQAWlKBoYFUIcCKIYo4KvTJN3h1QUhGJTSoJtTXcLM9O+NXtbQEWms1PjgGOZgIOXsPBghU8a8L7IqGgHVGTX1xqACm7KPVDBAgrFVD9vQMXdEqZtlqifFlDRbgW83+S4bVfaJUhbnOUBUFFvlBA20Coqud++4H5wR1X+pwEVtvkMXdPdkYr7Ayo4h+xkVETCF+mRFV2BR1nqiWNdXuiSfhKgIrzP1893ucVwsljx2F8SUGFZEmds7W7Y36vtJ409YLGFJautbXzlvPMn8ybVvkdDjackq6vIJpDP/alSIY4x4qW9dVwm5XUBreNli3tdpbnL3bBan3K0fHnJJIerWO6kCaRg2/o1lNfgmQu+w+3SLfPgcy/hcwbShg58YaJdzBAVP1ii2arq60bJ1iw2AFT97ySAlWx33gV8TxX1zlOClx4wKkIskxCU0hYvlaG3Y1B4U2axn53EtqrgKTcUSGy1nplrVWMs8NKZKFfyPGLeDN4DwgoT7Hf1l8vB+THlACOfUK+zYqgyUTI/K2fSLmDGMTA82MCCJcVfYjaaz4KAgqL97WXK2ZZkNjKu8HJLPKdn3/Bnxrh8EeQIcn9+z05GBYB/9b/bZ/j65jcMWDNgwvJO/ON9LtnvHAMyJK+RpUsTbcpSW0Gm+jdG2a6SniMr5qBygPl/eKDC2DoW+/kiSpP6NqaKE5CxixJQYWABj8fh79UReK8sZunsTAuo8HJajIFMzSLc18HTLul3f19saxbTkI0uZoUKY7xpuOUwKU3FPRTzb5oPHgAVrR+iB+/+/LbAvQIVwQLetHg1UCS1BjjQIvQQ3itQEaytDaCAr2yoGw75J7wObNgZAlQ79MzXqZzeT8JQfbc2m/zRPTEL6iUHDlZpWsRbICTBsGhcOBrR9xBQEQT8/j07QNivok7QpCRLi4jLARw7FytfcXC/Y9XRLt3XSMW1+KHZTJsyMCGgYjuPLRpqy6OCoIUlTvjvg0+GgApqR8ZiSgwQqBAdMB5DMp22CZ8b6hKBCoIIG1haWhDK/eiJx7G6vqGKOQIV1PRnRb0Q7IoZN6ZScVXxXb1ySf4Jkn4aofRTQhP6/oOHZLLaOzJoOuIOdCFIwQ09kysCKuilwcyWq8oz6ScuDlaR6l+qeEzTo8ICSx5P2uAVk64QwEG03S3GXOwJVCAexdjuPZaQ2s5hdekOUjRXXV1XVfFQ/wCqpSLuzN1GzwiBig1cOHMOpUIJ04cOB4yK3uFh0yRPp1VJu7WV088EKmgqztfIyKiTwygG0k9W3clgLob8NmUkCCwUZKbNhZFm2rw2Jsopt8HFk8nvvCo4E+o3Lv4bq6t4843XVYH9JD0B9k5g7/heVaSar0Wf2lVsj3xO1+P/rSpR51FB42/vUcHkHJNCZNuwkqAs/cwI4gmyRghUVFEr5vFHf/gHGBsbEVCxd2K8AahQwsVV4VBzkswDAhaUDFvbWBOAwPNTLkjm1qrarKEjHcPN61fwwp+/gE4HVOzbf0geFQQqOjIGVKyuGFBx+9askuMaOx6oSMawsroi6SRKP/3uv/4d/JNvfRuHDh4U4MBEIhN5TD7TRHZxcQGrq6sYGOyTDwiTr6srqzJL7usfkHRKd2+XaNzUhCcgOHPzJhbuzGNkaFgyMwxa2O+vvvoqnnrqKezetVsVq5EIK6tXMHP9JtZW15SkPHL0ITzzuc9iduYWlucX8JWvfEX9wj7zc0hXD5PUUQEVrNh/7otfwMjgoAJ+SWpR+qkKfHL6E/zwrbfxS7/4PHbtHtMzwOeyGo+KtfHuD3+Eg+OTOHb4qIAKBm9MbH3/5Zdw9NA0Do1PaRNZpP9GJIJ33n4HU+N7MTm+R4FmsVTBrbl5nD9/AU8/9YQSV0x+/uAHP8Cxo+ZRwXE4MzurBNmoAyo+eP99MSoo/XQ/QEWrdcFvgMJghE2H9bm4GaiwzaWjVjezJyImXxUO1P18EqbAe/DTNFUTYkqkkmnEopSYy+PVV1/ChfNnkUrE8NiJR8UwSXdmFJivrmVx6co1fPTRJ1hZmkMU2xgY3oX9Bx/C1L592DM6iO9+9z8gFqvisaeeRBer4Tt6kcuV8eH7HyDTkcT4xAjS3Wm8+trLmJrYj2PTjyMZ78F2PovTp99HTx+By7zk1/78e38sP6GrV85KompwOIMDBw6gq2MAyVg3qqUSVpY5zhcEsJB1dHB6GkePn8SuPQdQi2Rw+fIcfvj2D7C+egn5ch6/8Itfw8TeQ2LZnP3wPfz3/+1/g4X5LfzgjTewml3HZnZD3gm5TXoRFPHYYxP4zOe/iJ7+PVhepr/CALKbZA4QIKDkVAmpzjR6eghUFLC2dhuXL76DzlQRJ088jc1iF2LJQWxv5sT6Snd1o1CsYf7mBVy98DKeeeoYRnYdxp31JLKFmrGnInF0ZbqDjWe5SMCxpPWjVK06oKLLDM+rFYHYAipYucdNDRkV9EeIxZFkAp/m6WlKSOWQz9M3YlmyfGSjFYpbAqTyOYKY22KaEeAkkEsZPgNpLSryiQ35SJE+XougEo2B7ILe3n6Npb6+ITFZRkZ2IZMZ0qaNQCw3SdVqBLlcUWvr5va6pOfoeeNNrY1RsSmggmsef+ax+DxyXuDvuZZyDeD8ZesTgXPoGZaZdjKKSglYW9kUe47PA2XzvEdFmFHhv8u1KJMwA2/ONTpWiFFBkJgvggzeTNuAiriA4DCjgusyfR44nwqo0KbTzBTlqbRN43Cr1K8UqwKXw0CF3+i2k37iBn9ujkUW2+ilj4qTrSOLhJvbza1NgVXdPd1aH2dmbupcBJy5Vua2yFLpEYDPGIPTjQdmyYLZ2FgXk4XvUSrQKh4tMWXzi0llyP8knVRfhM20xajgBjpaRi1qUirsAw9UaP3PGENKVXyKoc2Em+w/Gr97oIJxxOzt25J+ItCi9oxGkSVbkJrMPIbz1zCgAhoT9A7zQAXHl2elMJbzQAUln+TNE4MSHWRUdNCsm/eaTf18MSp+noCKtsndUHFV89ai1XfCxVj3uxVpefx2F3Z/jIpWANDdgYLW522fA2/RTm2Aik8DKMKxRkOTtNwPKjqxOSD8YX+hLoFsv7qra7n7xM52bc+o4El9oWL9RAIqAnSk+WcvmWQXGOSq3bW3vIe2tf8eaHBSW06Cp337Orkhl5UNAwVtUwQ/JUZFePyF+9dL95hMjSXh1U0qb7eY0pLzTuYnLEXl5pdgTDqgws/h0txXYtqNTTfnq93vClT4HAoNo72Jr603VnRi1fJeLihAmloAYrwGyhX5/bIli012ySfNbf3yjAxbp9gI3nuBv9f5ZJxsFef8Pb8jA28HVARj3I0lAhFcS/g3982+ACJIWEseyVX+C6ywa/NJbKvg5yhxcttN85MvdPDJfkk0uWR3MI5Dcj8eFGs5LRKc8jJmrvRXbeKux5tve9Ntf11WhGqV/uofMTKMfVFnczsPDG+QLVNmk4r240v7D7UF2cKs5I+h4IoGzZicIIIl7AlOyJuBHhX0xHBjzL5r4JT36NTxCZ65uE2xnAN22I//07+st8ZvftPkl9TcVEdgkWKF+3UrKqEfhvlH2PnZFgJGBB4Y+5UAR7gwlwUWLAb08ZsAIPmOWFEP70kAjH/mnPF8nRHjYyGTGpP0GL0tyvQDoSeKnc9Ew0xCyz8fis9cv5hhvTEiBCCihlQqrWJZxoEGtjjpKC+hJYN6enw4zwreO/vhAVDxXxpZPPj+z1oL/LO/1ZpR0ciKqAc7wfU76pv9uxnBDf1bPzaHb86YWg+pm+jDthUtPt/YbnWoYMca0RBR1HUOGxJM7rwBSuyZHCFaZHNMx0qSBoDBodtmbtPcBj7A8vcXPppPlTUCGwQdGmJGNZuvJnBtFG5n367NURc3j0Fg6s8RBkP8tbjfNeMrOwZoHTTRnUqzPgRUOCpiS0ZFnuCEgRR1oCKP/Sc+owCCCxmTM2wRGVBVKihHbCNrSQ4zwqRElGQpCjksLc5rAXj44UewuLishmZFKJMnQ8P9WlysIrwgvW1K6jAJWy2WMDxJq8lyAAAgAElEQVQ8jJHRMUYcust9BwhUJNA12CPkncfp7emVbAUPvC5T6YQWPHaF3/Qbhc+q4Qs0cIrbAsLkKJMlttDYQkrdd+qLk0lAcMPTAqU56XS6GUgRQOCCns9vKYnH468sLWmR6+vpFdXx9uwsBkcGkd3YxNkffyIAZ3p6Gt29PZjcP4WewRHdj692pd9Fd0+PEgWSgapU1AZ8+X9rcY2ZVIYMVgslrK2t61qYPOAfmjUzwOCxlr1edU+PtMypR88kDhMQZFS89cbrknugOe7w7nHsnphAjom1UgE9XRl0ULqjWFKSTlrTMruyoJvHYvCV6uhEuiOjhCMrRSkrwntRhQMDCFBNKCGwgeSC/NYW/uxP/1TSPl/6ypexe+8e9A8MuEXfqrUVHLkgySp9ocTU8vKKjk+dawt+GagwCcJqmyquXLqEV158GZmODH797/19TO0/IPNSSjl1dffIT4KyKis0tSajYmyXjpHdzMojhewQytqQ9Cug4nd/V9JPR48e1X0zqcdEnjdhZ6Lq2tWrkvswaYwalhaXZepFaSrquxfLNO8dEEOFQJmZjZdkYM57nV9YUMj4h3/4H8Rsefyxx3DowAHM3p7B9etXMHPzOtY31rCVzSEeT+PA/mmN5Sgq+KVf+qUd0k8yJKP00/nzuH7tqjwqaKatZ7JUBAX4y9EIPjn7CX70+pv4K199Hnv27EYxQnkqS+4xWfjOD3+E/VNTmD40bWEb1YeqFbzw4gs4cugw9k0ZUMH5hf3z7nvvYWJ8L3bv3q0xy/a4OTMjQ+9nnn5KiS1+9uVXXsG+qQOqruazf3P2tu6BkldM3p06dQonTpwQoyLlzNWagYa7rcvhCi3/uUYwwmvHtj7K3YDweiKxUZqEc3gVpAhHEaklEKkZbZzVq9FIBYOD9DKIYnb2Jt568zWsr69heGgATz31NCYmDqFUigpw7O3rddqoUY2Va9cu49z5M5ibuy1QK5PpwOTkXoxP7sFbb7yKRx/aj+lDB9HbsxvJxC4UylGcufQu1vLXsWdwAh999K78TY4efhQxZDQHfPzJ+xgeG8LmRgmTE/vx6qsv48ixA5pj3n/3I5y9cEobyL6eYYwNMykeQXeX6fnnslnEk3Ecmj6K4ZG92NquYWWVvj5RdPV0olRew1tvval+/PKXv4SxkRG8/84P8djjT+Hjj2/j7NnTyBXWsbmxomRtFHH09vVjaDCBr/7yVzAwuAu5HBO7/djaLglMz2aZpOVmq4rBwVHkt0pYX76DSxfeR3dPGcePP4bNXAaJ9BA2sllVoBOAKBTLuHXrPC6cexmf/9wJDA0cwup6B7L5KjJivaVU9c7ND2WTuGnaypKdVkWlWBOgywQsf8dnn/0xPz+HaiTHGilJM9FjgvMppX62c1ls51ewTT+JLA2dC0p0q2pNG0dpspmJIRmNRcoiuCpLavMmUshkuuVZQNm4/oFBDA0OoaevX2bptonk3MjYgxVmtnZwreIawCSwNv1k7Dgjv7V1MnMS6Mx06nr5swcqUgQqqhUB5Dov59mqVdJvZjeRL+U1R5P5yHXfR04y006yKq+K9dUtbGxklVAno49G0jwGq+M8m0DFAREIDM44I0Q+eV460CSYTH6JcQXnHl4D50jGFbaJpZGiASWeFcE1iffZ1d1tVZnucZZ0VJ7G4WkzcaxC4DM3ielUWqCxWBT84wpfVJjgmDE+Xrhx85a+z0IIMS5pBulizs3cpuYyMirYl7Ozt1QZyHvO5bYk10WPig4HFnDTT9CiUqygtF2SDCPbmPfHtUzMTkoz1LwZuUlssX8p/cTNPIskaiWC/TVUy9xcs4qR8w6fjToTmusa52WyqkxqwM/R9bieFamqYCUAE4lg5pZ5VDAm4pgXUMGChiorXNlWLNigh5RVM/K6E/GU/J7YTyyukAxELKZiExaaUAaL8lgm/WQ+IFwPU5TLYmdt/IwCFT8BINFuPbpfRsWnJb13nKc5M/ypG9b2qfm2ZcY79nefepLWH7jbtbaTA2qz3wn2THe7nYZNYWuA5q5f953R5kM7+qrtwXb+Qu+0PX5dcmdnQ9aPpf3wp3TFfTMqOAvdk6G5P7El6XyBod4NPT8tr69tX9dNjOvy0U4Cq2XbhoEKVzziFRnaNUxLoIKXbAUoLdu73bl3jC+HMPN9Jnsd48LyBJY4Fpgs/wB66joZRCcVpaYLHVPfccC1AR5hfxLHNAnlQtrOQU4CSSwABxgoqe2KGFU5H8j61SWfmvtSQ9aB4bxOL/1kMkbuXkLm2DYU6gbfllT2uRGrfucA9mbWXu8/GNXheTjMjNDabf4dZlJtIIfF7SbRKGnMcFu66/CgfaspTa3jvSJ4Pyp8sEp6xmz+/n3hrZe0aj1sLMbTPTt/DJ5TQJEDcjyY431I6jkvb7xuRzZmgwFJ9jMZClSPMOAraFdXXMXr4zG5R2Rb8PfKf1QIApl8o5egsjnErtEDP5bwN5kmD0KEJb/UDo4F44EK1zj4lyGPit/6hjERPIRp3UmvLzORVkFvLCoWA9uEhTnce/Iz3KeKgVqp37uxFky2yvt/2P1bsbXt8bx8lusv53fBGMnOzr2fbVgFrlHRhOd2hTga13GLoa3YzBmsE/RSMavJ+vriDY4PxjUsbuLv5BepceT9MNzPvFX2Bc9F4I75Q8/SeQBUtJu6Hrz/89oC7YGK+srsGJA7AId6AqYZqLBH2D3JLYGK8ETgH3jfhjuZAs1RQiMnIViM/SnDi637pX+IdV5nrOMXF/87W6BaRyThiclPoqIyBp9vAh6aL0ondpCG/mo+T+CSZZNkqLpF59B3veyTaymVvTVFPU7Syrdlg7F4wykbz9/qtm0fYOcMIBdfdNPAqCCbwlUeFsPST2RQNAEV23lMPvKkBRxVVosWHCXUqveqMZtwPVDBJIEFCTVsZzexurykTfiRI0cFVPA4lMVhQnhweCBIADF5QqCBC+Py4iKyaxsBUBGh5EK1ioPTR7SgRjvjyG7lVIk40DcgA1m+uPGvoW6MFAYqzLSqLMYEF32+jFFhFZ4e8WfVQbnEBdF7VPhKRws6POo/PDyia6KMx+qqARQry8s6XmdHh5JCc7dvY2RsWAmacx+fFlBxaHoarHif3DeJ3uFRJUeYjGBFPM2ue/uoFW7Vr2xHVpnzxWSPDwg1/t2YLORLqto1oIJJDwMqeG09vb26Jv5M0IKJN2p2M1lJoGJjlUDFa0rWPfnUExgcm8Ceib3I5XPSPKc8V2dHGpViSe8xuLHK1SoiMTMOZYBKs9YOARWmvc0KYhqsSr5JJlsVJa6qlCuRNFgR//lP/rMBFb/wpTpQAWfg5c2w3N9sD/UvDbCXlpRoo+mwksBRYSZIJplIqeDc6dN4/ZXXBGD9+t/7rzAxNYkCzcficWQo8xKjCasBFfSJGBsd1YaBwEpPb5cSeQRC+N7i/Dy+853v4Le/9e0GoIJjnBXDDAiZxJK5dqkgYIO01LU1mm1XlGxknyTTpJQWTEYlncb8/LzuZf/+/ZJVYVsnYnH8u3/373Di0Udx7NgxTB84qHF18+Y1LC3PK+gkE2RtLYtYNKm+PDy9H7/yK7+ia/EbAgWbDIydR8X1a9fwrIAKe9Z4HFSjKEej+PjMJ3jnzTfxV3/xeezeswsFVBFPsmKaRsEEKn6I/fv2BUBFNWoVy99/8UUcOTSNKQIVbuLifPPuu+9KZmjPnj1B4Eg/j9uzt/DMM09rzNC876WXX8HU1H50srq6XMb1mVtK8I2NjalvCVQQxGE1d9JV9dwrUKENndtQhdeGnyZQ4TcUzWtPVbIJUUSJ6CgvwiCamWgCGDnMzl7HRz/+SBIrBw/sw1NPPoVRArGRNAqlGj744JQSfgcPHgwqxHndBH7v3LmD8xfP4dbMTc2THR0EUsuolO7gC59/GlMTx9CVmUIk2odasobrt8/i1pUruHLlLD7zmSexf+ow0okebGU38fHp9zC6exQb6wUcmDqC77/0Ag4dnsLY2C7MzS6jWMmKwXPu9BVcuXwW6XQBwwMZ7No1JrAtmY4j3dmFeKIDA4Nj6OkdlLQbAcBLl88rQXnhwgWBtb/w5ecw0Ee/iCrefPsczp45g7X1JbHb9uwdx0NHH8Z2bhtXr36Ar3z1OUxMHkShQJP1HmxtV1AUUMHNaAWReBWDAwQqilhdmJNHRW9fBY8cP4nNrTTiqUGsZwliGlBRztdwa+YyLlx8Fc9+7lH0ZiaQy3dhbauErv4MUrGoqs65JvP55fqQy29pTBJk55zASjWuCUw+M3lO4Hc7uyJQgnNvgeyLUkmgAzdaZJMoOeQqupjw1XhkFWU8KfkqAgseaOjt6ZcvEOf9zq4udHf3al0zersZIUdYMYYocrltAdOqLKSXSDypZDir+Anws2989RnnKA7Bjc2sARqZTj3TzUAFN1qci3p6+rQOcW5gJT0ZA/nitp5BAhWi6RcNsKGRdixBSYEqNtZymuu5LlB+ygMV/LeS2ZRtcprRqysryKRSZqTp2HledqkZqCDQ5YEKO0YLoGJ7W+sswQIPTvJ54VrK9ZLrBjfB5UpN4DPbjYwTvnxFXjwEVEjCK+l8M2JR3Lx5W5t7Fh5wnjM5SYs517fWFWqxzfk+GRUdAhzSYgvlCg6ocEbfPJ/m6XINha0itre2ZKZthuMdBr5w4xyh1Jf3ojLmAoEKrjXbhSKqxYpACv7hJt4DFZRs8Wmuhbk7+rGnu8ukRyQx4wpYnGmpZ/1ybW4PVGyh7Ao0fPsGZtrptICKpSUD5dkHnh3DgoLc5qZkBM2Xx4AK3n9fX6/8zBQePwAqfNgf/N0WqLhrErzNL1u9rWFwr9n9YIe34zp/ojf+XwQqtP63A6Bavc92cjnbVvfasp/aNWubxLzfIu7sjrsDFQ2X6/7Rbh/8lwFU+PXOBX31sdxmkHhD5uZfhxmpXvlBe/y7jH2TrrGXfd/LK7U5+f0CFXc7t/NJCX9EHkP0InDAuQ15S9YzOjT5I5urCa2bcbVt5xpACrcGMKbw65VvX1vjGVPU8x9hv4kddx6SKbKktiWrmfDV5skl+r0fkQfAdE1Nz4ZV7Fs1ui8kM0kexxbxvhveE8LlbpTkrTJBbr6Rxg6xhK+xK8x0mC/uMVqNcf7Oktm+It+8DQLWiits4zqjPb1YGq6gKJRX4nlbtZdnGPj247rGF/tM7AiX6PYAg9qmPXVHHgt+3VdxCuWElCg39iyPa6wBk/X0II4lyO188phQ/GSFHNy/2f0RBDDAQcwPFqBqjrNclGdDKG6jH56AHosbucfiPkP973JijJN8rMbzku1grE3zauAf5iR834v5ohg0rj5U0Wq5jP855FHxW98gC9fl0Bz7gJeo8UeQin9zLOmZqKjwURKXLMSJ0DOuKM9R743m778uqcSYjNdhBt62B7bj217X4kwevwGoUIPxvFR8KCse98wZzWXO1yKcX+T4ZPvwPuV/Kj8Rv0AwtkkG0t38HtuPY9P60FQ5PMgkP444cwJFxX8PGBVt5uoHb//8tsA//frD9YtvVzXQ5vaCSbsh6b4zAe+FmfxhLHlulDRFbwGmYT8Ek0CT1l6QHPIoZwO1PQyMGNK54xW81UTVCwMc7YCKUIVE/djhc3ifDn9Wn9oPgRMCERqvygeE1kYBHOA+VN8Mqq0V6drLJkD/nXrL2k/166rLYdWZFq27M/SdUDv5y3XYsk2QNotrsZIGI/XxWNFJiYRiSZt6D1AEQEXOZJ/IsBg99Igt+NQnpIakozBysUI8ouRvM1DBhSe7voqNtVUlDA4ePITl5VUtqFzA44ko+gf7tEAoAbS8rIpOJkuuXb6C1aXlAKhgNTyDu+kjx7TB3a6yMjSlJAoXhGSCMjkReStUa6ZdacGALfYEKfiHyS4CFb4P6VHhr9tXZ5C6J51DVrjSTNt5VBglkIu+BQ0CKmiwmtvC+saqzklpCwYAqYQFH5QWIlBBn4gLp88q0TN96BAy3d2Y2DeB/tFdolDyGtgGrLIks4DJCQ9MEKjg9fp/qx9aABUMfCzpkVbCnO1PoILJIf7MqlMCFJRo8h4V66urePvNN9DrgIq+UQIV40qy5Ap5dHV2oItAhfwhslrwrR0tUOWxOBYIFHV2dKlfmWBikowSTUy2mUm9GXjRu4RgDaVk/uSP/wQjoyP44nPPYff4HvRTLks0yjqjgvfJdpW5J5ND6+sCKtgWiQSrro1eTdyJiVv2xUen3sd7b7+L/r5+/N1f//uY3LdPMi5M3ndmTIKJQAQTe/NzdyQvFKeMiNgsGVWAsi8obzZ3ew6/64AKggd8inl/DNh4PQzS2N5MjCUT5mlBAI2a7RxDbBcGNHsn9uD8hXN6DpjYYvsQQCJ4lO7s0Psci7//+7+PRx5+GJMTE9i7Z68S3AQrKNfDZA8TlXO3F7C6Ykbgj508jl/5lV+2YMdtFGQmxsAsEsfZs2dw4/p1fMGZaXMOMKDCGBUEKt5940381ee/hrHdYyjUqFtqciwEJMmoIGvCMyqYiBdQ8f3v4+j0YUxOTjbM2u++9z7Gx/cKqPDVRLOzs6o2/uwzT8t8vhaJilGxf98BZJIdGlvXZm4JsOFYZ9sQqDh+/Lg93y6wvxegoh1I4YNYzbSfYoT9aZGBD15bghVuXrQNHjclZURqZSws3saFyz+WTBjlyh4++ohk7dIp+vT0oxqNoyPTg7m5OXz88ccYH5/A9PQh24BVY6hVWC1mdG9K6d24cR03KB+2MIPc9jXs2T2Izz3zOQwP7kMyOYRYqhvRBA3i5/EXL/wxjh49gNGRPRjoHUa1WsLpM+9jdPcurC3ncGDfMfzFC3+Gg9OT2LtnHLdnl9GRSWF87zi2Ngv4nX/zf2B+/iKK2+vo6OhE/+AARsZGVRnNPuvMdGNoaBjDI6OS6PvxR6c1Hsf37sF3v/td1Cpl/LW/+leQTHXildc+xDvvvqdqKfb1k089I/Pv69eu4+L5t/D5Z5/E0YePo1qlv0Qnsjlbpza3qM9fRiRWw9DgCPLZIpbuzOLqpY8wMBTB9JEjyOe7kOjox+o6weIEerr6UMlHMHvjMi5deh3Pfv4EejN7sZ5NYCW7hY6uOGoVMpRMbmB7O6cqeFaDc37M5TbNg4lrZZESiQVjGqxv6Pe2DiYkxxOjRKD7E+/o1Gac6wfXAc4PBMQJKPT09aFvcEBzfi5XwNLCkqrs9+3bb5VuNW7WUmpXevxws2mmjFYNR1DEyxryPVbwkwnBRDbl57j2+GeAcxLXe85HvB6aPu8AKjpNP5fzKiWlBFTUoprjNrey2C7kBK6KqcH5RXIWEcmVRROMBYDN9W2srq5pE0eggv4MLNLnplJsgGQymC8JfmVSyWDT5hPbrRgVvAbOZVwbbTPfCFTwOtgfAiTkUWEMJkY7fJ/zCK+dG3BKLa2srgZyU7Z5NI3jVkAF74X9MTMzZxKIPb1mUMkbM19QrGysSsqT8znnhFszMxr39F8g+43AvhgVIaCC90t6YX6THhwcY5QpS+m5ElDBDXLEEhqSBokag4TsFY4ZMioE9pfI7jADTg9UELLg+sR2Wbwzrzirt4f+K5FAh9wnVWxcuYTJ3YAKsloqxqjwgJLAmkACLCmGo/ez8gkrrq/bZDalWMhg+ufeTJugFyUQFQlvJCWH19JMu8m7rV0i9tPm67v/vrXcUFtCxX3THe5y9jYJ0LZburYJU+cMeq8N4bOirT7f9sbbASH3C3jsTHz63VG7+27HSLnfdrK9685Xuzyj3dnO+wvO636leCDYzoX3qaHvtmvX4ONut+az1a0+70Ce5ivy567vtRvv0e/NG3acYcmgHbfYvEe9C66lyzaN/Oa2apXkVlK0cbvb1CH1iwk3Qfu+rkshBfsil/Jv7u/g0fVVnA3dY0ncHa+GwsbG8eAT18HteMWGUMFiXULJRrHJydRf3tI5DAaEf1YiNQxUNPgiRARUBAxfl+T3IFCQp3Df8fN9+PzG8mi86/r4bj32zQeBEkyugI/V7fJLpHdB2fWv7Y0sqes8GJxXA4El3hdfTFabTI8l1vkd7b1UBGZDivtoFlfwZ4EkTiJKSX0xFMybQjWhbk3z8j8+D6A+cuCOEtsu6e/lqrwxNLuQn2PyWtevhLMl+nc+Jv6duveojz/sHk1yidfGdiFLlrEK98TcN/PamIdhkQJzD1R6YJEDpZLlyeUq/AWShEzBNQrFqrAGYnyizExIad1A2XB+yFiVzG2w3dS+kv2yvhEwolyJy+cJJDEgyq6J8qN2v+xTxTGU6CwUFLf493jN/yLEqPjWN41RwUIZxvzGiEhY0YdjQlQZV3JfWmLxqjPOdr4ajH0Y83pARBJi7joMlPBsCp+zc/cSsHpsnAn8kPyVz8cZyCBJrIjFQj5XpKakCbqT+tQ9O3aKvs99P+N7B9zw9wa+WSELjyVAo+o8XARYuryRk9DUfSiPY16oD4CKnVPvg3d+zlugGahou4i7+wwW/JC3QziB3swUCBLwoYgiTMO0z9eZAjY5hxb5MGMhdPKGhdP3QXCYu9yFD970ndDn3I/tNjBBoBJK4jfeayuggpOxq4B059L07IwKw0GJDz0ar8lFngrgfBhiN6vPfwpQ4abbhhHacivQ0Dfu4+4+Q2GztVcAVDDJaAsEF5YSEzClEgpF/mkDVMijIo/BfUcbgIog4OQtJakJGA/kZ7gYy9OAWv5rKzIMZaJm+vCRAKigZAGTTkwMK/njZIIo/cIF6OK58wIqmEQeHrUEGBcBMiqoIR7tMLkQJnUkPZTs0PdYoVitsdLTKiG8XiOT68aiqEnayScZeV1MhPhFj98To6Jc0WJDPw0uZFaoQMomzagMJR8eHlXAxkrbDSYmHCOCFfZcjLnwMhHeP9QnRsWFM2eVqD8koKILE1MTGBjbo6CNCR22AYEEb6Ts25EJPS6QTLw0MiqsUoTyV2aYXQ2kn1j164EK/o7HYsUuGRsMjJhoq5bLWF9bxRuvvSqz6ieefAL9oxMYn5rA5vaWS7R0oIuMEybyivScMNomX0E1hRJXTMbRALyGTUqeFIpYXl2VlBeBCuryy/wsX1QCY2VpGa+9+poS3V947jmxOJSwdVJRbGsGDmwbjlECFTwfwQUCWgpeE9Rip7FxHahYWlzAhx+8h3Mfn0Vfbx/+9t/5dRycPiT2UC1KoCKj4IDMGx5rbva2Eqa8Nkq1UFYnkYorUUepKkp3/R6ln771bTz00EM6F/tJYIAzFreKFQa/NVW9M0jd3i7Il4FMFco/TUyN4878HY2HYQIj8ZhAB+mSR2sYHhlGd8aAimNHjwqoYCI7kaAk1bp038kYYfy4srSO+flleU8cPXJQjAqOn6BKihsbVeYm8PEnHwuo+NJzX8SQl35idrESAUfxJ2dP490338Jfe/5rGB0bQZHeJ0y4xmKqDnnn7R+quv/g/gNGXaduF4AXX3wRxw4fwcTERD1wBPD++wQqjFFhz1RNkkUEK5556kkBFcxcvfKDV7Fvaj+60xk9JzdmbzcAFR988AFOnjypJGAspDEbnuub533/71ZARLCBuUeQoh0oEj6H1oLm49VUI0c4F9FIFdu5Ndy4cRUXL51HdnsFe8fH8cTjn8HEnilcPH8JS4tL2LVrVMlGyvtQ5u3OnXl8+NFHAjT3M4EdTaFaptyagfkcvxz/NBueuXkVN2fO4s7tqxjfO4gjR6dBDf1CKSFZJlbmv/TKn2P37iGm09HXM4jBwR5cvXYWg8NDWFnKYnL8MF548c+x/+A4pianMD+3BtrYkw20vprFa69+H4n4NmIoo7OjByvra1hZX1USkolgXj8lfwhc9PYNYnOjKN+AI4en8cO33sTbb72lMf3Vr34N+WoCH5z6sQzDOzM9OHnySaTSGVy7eg0XT7+Gk08cxcknHkc00od8sRNb21WUylVkcyUUKwXEEsDgwDCKWyUszt3CFQIVgzGBJJ2du5FId2N9Y1nPSme6G4WtCu7MXsHc3IfYPzUMVLqxsRnD2vYWythGcTtrjK8yqwtZyWUShFy7mJSXYXVA9/batgAZfklVwXeIWZLq6EJnVx86OrswOGCm6ZxTeAzp/lISh5WDyQQyPV16b3l5TYwubvQI4ktPGVWxI5i4JctE649PwNMjI5cTo0LrQITVeAZyJlOxAOgX463GOWhbm7PNzZyOR8DEm2nTV0nyeZm04pSN9Y2AUUHZJjIqBDgXt9HX36f1WwmRqhkqEpSNMOdeBrayBawsrxowkSETpohK2YBszkv+vHxeKAvY4Ta5qjpzkowCDZy8kF/rPCDMY3DDSqCCc5CXfuLnPOvC+yP455NrMX9H6ThWBJYrVSyvWELdy0aFgQq/lnHN5x8BKDEaTM/pWevp6g6q6Xzss7S+rPCKTAKed3ZmRj5djCcIVGRzdTPt8H3GEUNuY1uAGK/T2qhD/a7NLv8nI0dNlboWAhW8HjJDKP0kkKIBqGDL2FrI19LComQWCVQQ0KLUQLi6lBtt/5JOuKSfZtS/mY4O9TfHLD2hGO94tksgF4GaJLTisUagguOe+sv0acpJnjGlhEoYqCDolXZm2tWNxM8kUNGOcGAx/E9pA9kOqLjf3H+LJPFdr/Cu13+fJ28LbLS/gnAitv6pxl1L+Ns/LaDCURzvufMsXd/6usL+4o2fCTdu2D+idbtaLtGqgD2DwHsK7uimnzJQcZceairA80lPfz/hDTl/ZvK4McnfDJ74c9XBgruMszCAYOWRDgNpMXB9BbnprFgBmru8HdcUPmXT6RWr3gtQ0dAHJqMUSgfbqf0z0fR3HagIf8Mu17MqNBpCz5TS8s6fwBQBLPHtwQjGFD756gHkABwJMeg8mNbc6h6oaDklBP4KO0eK31f7c3s2gIEmVtDqGReSUvILkzc690WPFZol21pkxslWWe+LgVf/WgsAACAASURBVPwarUR6kKy3fXxYgtXvfVRAZ2iDeXaI1GwziAH/Jg/pjbCNgVAvy5XptSuMoi8W29oXy0n6sBmOc1JawXrhxl6QFPcyZIai6FqYW/AxiE9s22WYTwPjNg9OeClFfs7LNdXHiEkQGWhR97fyUkX1NcwnyohdWPGm9YeSVEHnahlxb8vkXJKkENNd8k5ifBgTxxrCJi09O+53ZFb8jyGPCko/8TRe+oqf9SAQ4xIWwrIIldfDvgjYJfJqsxyD9w8NA22S4tJYMx8IG3MhdlEYqIiY+Tdf9XZyY0LFfU6xxVJ2xg6pllUgxbhFQEuiHi9xfJAJob1YCBizZ8FM3a2NnBSZa1PtFd3YU1uSlRyPKc5/AFTc87L84IM/Ly3wT7/+kC610X/hboGh+53WcD8xhSWJWi1TzUta+DP8ufk7rswsOJV9JjATcnTD5oU4uOpwWYtfqN17QVgUANh27iAYanvr7gvBpTZqiocRZztg+J6b7lG/CrUdp0h93gdoTZ93wIYPPm2BMzrbzpdnToR7tOUHW99p00GD0KkeLVo4JXMnx6ggq8ExKgoEKwoOqCCDgtJPuUaPirHp4zo3AY4CpZ0opVOziT+ajEmz3PQEmdwx5FwazOs0DzWd7+PHH8XCAhPoXBk42W8rSUuggoloHoubfE7458+cDYAKelRQtofJpD3jk5KPGdozovNFhIZHVc3PcxOoIEbh5Ql8gOMrN9lf1K4WbS8alRGqZ1Swh1htTsYFE1SqZKReInUfQwGBqhIiEQwOeUZFDmtrq0pg87wD/f2i9DLZxYR8V29GVbg006aEUhioGNq1V/fDZAWrWpm0JVDhKZhsS4I1/LcHKnzlkBmQQfIj/C6vmffC6yZQoSrH3l5sbmyojZkgJ2jBZH0ht41apSKg4rVXXkFfTw8ee+IxDI2NY8/EBKi/vV3YRqazAx3UNN/KyYejoupKq/BgoEKWhrEBemQcTVYHgYpcoYSV1XUXIJCaaVUvy/PzWF5c1vnPnTmDickpPPvFL8pMm9XzfKIIRFlysKIAgdXM0syOW9UwgQqjTNKImdUWEemMk1Fx88Y1nDn9Ma5euCLpp1/9+q9h+shhlBi4UFe704AKMm8IVNy8fkN+CpRdIuDU0ZGScSmlnGiOTiDj937v9/Dt3/qWzI45RtjPXv7L+1SoaghVARscj5SleuWVHwiwmp4+jJ6+boEWH3/8YwV+TPB6LctSpYiBwQF0dWbw+//230pq6fDhwxhiwjMRxfr6Cmq1soxyE/EktrJ5LC+t48zp0xgZ7sfzzz+vPufLvFlqAh8p/XTm7BnJVz37hWfR18UEack8KipR5GtVXLxyCR+//wG+9qUvY5DG9nEgm2OVTALFfAEfnfoQh6enZe7NNq+66tjXX38djxx7CCPDrNC3AJZg5ZkzZwQ+EagQK6NYFHgzNzeLxx87qdmSSbE333obBw8cQk9Hl5gbt+7Mq/LYMyoIVNCjgkBFM6NCM3EIIAj/7IPVxqC2cd5vB2w3T65hYD18znYAiceh6UcRiZSwsjKHc+c+kSQMA959B6dw/PhJjO89gHg0jexGFjeuX8XS0h3EkzH51rACm8/AubNnsbKyiocffhjRWArFglVEMTnIdcho41axRubG3OwNLMxdwoEDAxgYyuDsuSsoluIY230Am1sr2L17GLlsAYXtCnbtHkIyyQ1OWUBFV2YAp069j/EJsiToGUR/EwLaNSzOL+Hc+Y/Q35PA4QP7sHvXFBaW17G6uY7FxUWcP38G1UoJu8ZGMThI4/ghpDp6lMzuynQKJLt54zquXL6Ixx9/El96/nlUa3Fcvz6H7FYZ4xMHSVLHtWtXcfX8jzC5bwRPf/ZJJJMDKJW7sLlVRblKb5ocipU8Uh1x9PUOoJQr487sDVy7/GOMjXUpYV+L0JOigmyORvYFRDjGtyvIZhdRLNxELFJCpUR5ugwhCpRrBVRLJtHo12muQQSjKbWUSveIUcc2SSbIMkrpfYKQ8a60fHmYOO7qJrOkG6l0h9a2ro4kqiWT6aOfB+cvShXwj/q5r1fP6fydBczduSNWDdcE75vEZ4+STkxim/xg3PSuq2Un/VSQNCHp7vxuZyfBVQIVSwGDgePVgIoa1tezSHemA2YDqwkFVGQ3xLLgzXNOo+SUQPvAoyKLQrmAoaFB+RZoLeUmm4n8WERARblcQz5XFlDBOYBzZ7VGwMc2mWYU3am1i9+n5F6Hk3HkNTYAFS7pwj7g5z1QYUAMKxCLSiaxOEFFBDGaaZs8FD+jJISbFyQjub4uaUGGPqVyDYtLiw1ABT+r+KVWDSQNPUih64rHMDt7R9V4nJvld8ENqDPsXllfoch4cO7ZWyZfx7mY/jNcQ72ZtgEg3JBHkYgkkNvIqS14nWyfRkaFmUtavsUAn0TSpC4qHKsOpGAigfMAwV8Ci3yeBXZVKgJACVTQo4JrG+XTlLZxeuBhoIKxDX9HLyHGdB6oYD9vZDdRLBetnSTRYcweviw+SolRwSrR7u4u9Q0ZiVxb5VHRkRZjiUk2AhhsA14TYxC+KhsEvcgYMV8kxhYC5xif+Y2+31OE49x24fH9Js6by4nb7iX8RTi/t0/73L38/qcCVDg5o/tietxFAulervu/5DMucbfzEHcBKu7CRtixZrtEst6/2xa24Yvtk+bNIElDMzecy+81XfFbcM3u/Tan4B5S5wgBFZ/m77ADuGk69s6deQsQoe0tK7Vre+GgItslNHVPIdBCbWi785ZAhcMXWktktWa3NGyQw/3uTt1u6PlEfP37rl2bvhDaEjdkMAyoaNEo4Vyu/7VVjLgB1vgdNZt+5fvd/g5/yjerP4xPXlrbNl6wT5IbU858FYPqeVc4YN1gifkwIOD3h0rYh9oyOIVL0HPub+np3mpuFCvCkr6eGcG1kntzL2sk3wSX4Fcc7lQNmjM29aIfq9z3ptJWUMhj2DG5r+C+WMlsFa/ZWmSFqGZIrjXM+zdwraHygZLFjnHjRiqvTXI9zn8gzKTwEmJcQ7lv8cCEMSucFJWv5g91kwEi1qo+g6PrYYJbe2UryCCTg33oZYyYYOd9B4l/Jd2t8t6knUwKyoye+V2r1OcYCFg2SrRbFb8NO0vWh8lj4ZlVxtVu/ebnjBVDCW+ThuI9e3CAx1ORjZMV5nUyhmWbsT94IZLWdPke5jv4+7D007f/kQFKVhxrIJDkfxm3KO6Kq6iuUjMZcsYc3HewTxn7Mgb2klccFyxwteJEZzheZWEdQYSw56Cbk0JzqoCXJqBC0xzPXfZSZr6YlcBKxApiZUBeULtrTDkwzfrQckhiBVGalW1YNbaJ9YcV3zBXZgodMfOuEHBj92wkrNoDoOK/JKZ48N2fzRb4p796rEEXr6VkUngi9fFE6L27MSrs0XETb0MS3E+GPH0zG6GZUWFsAh8AWCVoSAYpZIzU4vLqV9oAYIRvIBSOtQlkzew69LlmlCBEjQtiLlbNhxkh7pTeGEcrnF8UNOnYZGOvOlhhYLNLgITko3Y0m/teECQFSZPwMe9hHAbXVP+eD0g8DGKVBR6oCHlUCKgoYDtfMAPtggcqcpJ9InCx79GnteBwgeLiUcqzHpsLShSxVAyxRNwtrsbS4ESuisytTRTzlBtK4sSJk86jAtqULq8soqhEyJASt9zcClCIRHD+3HmsOUaFgAq34BOoYHK8b7TfLVAW1HQQqCiXVSnfDFT4igOh47WKJBd8pQYTMEwUmCEXF9SSGApcfFnlyOtkXxK8INuCSSGfpB4ZGRMIQL8BYzRYwmRocFBBHNkRy4tL6B3owfrqGi6dOy9GAT0qPKNicNdeJUS46adsFJ+RPhqnJo36GQYqPMPCVw2FgQom1llpy2QKj0XpJ/YXWRSsYt3Y3MBA/4DkYvbt2xcCKlbw2is/MKDi8ccwMDyE3XvHlYikgWxhO4crFy9i5vp1bKwSZDJdSq8xzgQSz9nb24fd4xNgmwwMj6C7bwArqxuSXGICJZ/fxJ25O6DU1EBvHwb6+vCDl16RZMyzZFSMj0vyii9SWQWoiVJsCz3blcFCa6ACiNPYO5XA5Uvn5Ydw+dxFdKQ78Te//ms4cPAAWKDhGRUkTBGU4Hi7evmKJG4YYLHCmMnVpICKdSRjcczfuSMz7X/87d+WbwQfM45rX93igQpVxtRoqDqrQIsMn9dee02JTlaTJ1JJJWfYx/QPSaRSGBwY0HNDyY7u3i709/aJUTG+dy+OHjmicdSRTmJlZVHjsrMzpWTi1iaNZov4+OOPJFvy3Je+qD7nM+fHJp/ZdGc3rly7ivm5OTzy8EOS8eIzwqAtEUliu1bFlWtXcOGT0/iFzz+L/oF+RNIJ3Lx1Gx2u+vrS+Qs4eeIERoZHNEdI5i0axTvv/AgPHTlqRuHO9J3j4szZswIbCDr56igm7QicTU8fFFDBP2fPncdjJx9HOmZm2gvLK2ofMqp4nnfeeUftzbkhrWfQ2BnB7OZB7CbAIlxVE/7s3YCLVrOrrxTj78KVW61Ajvp7NcRq1Ccu4ObMZZw58xEWF+9goK8fDz98HLvHJ9HTN4SB3lEk4xklntfXF7G6No9yaVvjisE8k3YEgwkuciMxPLILK+ubMiyenNyHdJpJY7KILGlIObNqoYZL536Mm9dP4cixXdjMZvHqq++hlsyguzeNPbtHsHtsCnt27UOpzGMvY3Agg9mZeUSQxMbmOoaGuzW+UEvzgcLSyjLOfHIWq6tzmD6wG9MH9mNjvQRE00h10ey5W0bt//H/+g8YHhxAdmNdknZDI6MYGxtBXy/lgoByIY+FxQXM3LqBfQf34XPPfgnRWA8W5rNIpntRrkZw5cplbCxcQy2WxWe/8DS6e0ZQLGWwma1hO1/CxtoaCsVNFKsFmW+vLa1jdXEelfIqDh7Yg+WlTVy/fgfJjg6Uq1sq9Y9UuCmMowx6T8yjVsoD1X55X6AjhmRnEt0Zrj39Yl+xXSlDE3Esurwz3RsaHpUxOvd3ZK3NL8yjljL5ArJaurt7xCijvi7nx87OBCrlgjYuW9ktJY4FUuhPRD44BC/m5xdx+/Yd+RoYUMG1jybVTGonkdvKm/ygPIFMi5eJbT4fpSI3R5Sdo/Fxp5gmHqjwoCU/y/V+bW0TlNoxGr1J1pmZ9gY6MuYVQEmmvr4BzbMEGTgWmaQmiEqWD6vgtf4Xac7IREA18KggUEHvHB7XAxUEO8JAhdc29oyKcAGBLyIwth6T1MYe9Mw1z6jgesSYw3tINAMVAplc1RoZPZzfOQ/xeSqWKuo3bba12TfwUuCG03kWmER/CoIKjulx6/Ydfacz3SHQhQ+eNqT00dpYkYygB0noR8Xv8/rW1lfFSCRQQQCLCXq/gY1H4ihkCwIz+Iw3AhUR1KImr2dZKwOB2wEVkqtkUofeOLWymWuWzeOL10mPCsqDUb6JWtD+vn0ShvMbN8wcJwIqyKjo7BSjoiVQIY1sAyrknZFIy6OCsQmLTQReJOICiQhUiFFBoILSUbGI4hqOJY55vsqbP0WgIpw4voeQWR/5WQQq2l1TyyqnnwCo8Anne22jn+bnmvZ99UP/ZQEV7RCDVjfZInkd+nqw7WvYf4ZhgtCH7wZUuP6wOCKk39JcDhhgB00H+4mBijYgSsjrpqFV/POlfXN9dxnOFwQxV+jQPxFQ0ZRY1yXd5eVjw4bikhYn1pW76nVfEc3D3hWo8OdtuCZfdBg2t/b4xU6QIsB9vOBC0JYO6mmTw2ChlkkE1RuAe25JLjeND65/vrrdfmnMA7VN83MXSriH4+pwE9v33DsBSEU2qSV05XvgkuRe319FYy4uVSEAk/Guur3ejHUDdEsyG0hh67fbWyqDy1yFSwJXjYXApH2dcWFHFIuCCXYnzeiNqU1myGIC+5z+q88TxFCbio1PEN0q571nBv+WfI9jWHBP6j2d7Cj1F9vAkxN0LidxRZ8FH3N57wkVKqhPzROTnzd5KmNU+CPz3H6dNR8KA+/5OQIZ/L5Yis5Q3OIe25uRZcNcRR2Qcu3kngczkGabG2uTLyt6csJkTnXD2qxuGq3CQcfWpZwm249xEmM73qfyLPE4/od/UW+d3/yG5ccovZmMJyUVxeumXLcYzF7Ki9cE+kxSJrQY5BfYhmSayqi6Wg3Ow3YKMyo0boJnpBGoMI8u8z1p3L8ZCGTsJDKTrDEs98B4yQpYDJww8EEAFtU5xACOKTfBNmKugddYH8e+OM7a2heGsEiW4y2d6VDBLGN6xpUPGBV3n98f/PbnsAUEVPhXwDpoX4HfnI+3r4Y/3+q7zZFVvSrVJvzGKlWTxQm9XNDlNfuaP28T1M4r8TPnjmP56owd5whVLzT1ZdjgO+z7sIMSZ8tYA6MizITQb6VZYs1mP3Hya6wkqX/H09Dqpq7B3qAZ39HBd/ZFI/jRepAa7bQRiGmo3PC/c6UbDBg4CVv1gfeoKCPvgAomNz0wQcBiixrKDqh4+DNf0uLOBJoqHbeZ9DET7UjCKGxctCwAMFYFEw3RahnFgkkpPfTQw1hbW0dBIAdNPtcxNDKkRAgXr8XFpcAYitJPYaAiSmZDJIIjxx5S93UN9GgBqwkEiqiyVD4blPSoGPLtk5NaKJR4oGEXJVPIqLDqS2mHZzpVEai6xFpZgA3Nvm0jTnmhGnLb26pEZ4W3Bwx4Tzdv3BSbojOdRrojjYGBQQwNDjnvim0sLyygd7AP6yuruHz+AkqFIg4dqgMV9KhQcoRsgRVL1lJnnAs2z8MggIwKT4n0upUahyFGhWSj8gRXrHKWQAXHB+WxmOSjyS0T4WfPn8Ojx08IgOAY2FhbwatiVPTi8cdPYmhkRPrzq+ur+PDDU2InrC0vCdioFrcR8VUQLjJTdQAXbXo1ZLqQ7sggke7A1NQB7D98GP2Dw/JYmLk9g3QqhV0jo5I44mPw3T/9M7XX5579QgBUsE9aARVep9wDFWwHJunE8HBm2hFUcOnSBVRKRZz+6BOxWn71638bk/v3ocqgnRW+mYwCC8p/Edy5fPES9u7dK5kngk2UIuO4kpl2NIalhQV853d+B//kt/8Jjh494qqCN5xBaJ1FpGAmWsPMzIz6jAyfN958U1qkhw5OoyPTqWeVx6aJ9//N3nuAx3Wd16JrBsAMMOi9d5AACBJg703sRRTVuy1Z7rJlp9hW7Nzc+25yY6fdxIqbeu+iCimxF7GAnQSJXkgQJHrvdYAZvG/9++yZAUjI5eZ9302eJpEJDE7dZ5+9//2vf61Ffwn+jRXNZh8T/GxWYVDs27cPqUnJSE5JRnhomEi69HR3gkaprExldXd/H43QTSguKoSXaRybN28Wo1wGkjQvFgo8E9zRsai8cgWlxcWYOSMboUwcG/Vv/r4BcHibUVJejounz2D9ipWIiomCt82K7t4+SZQy0Vd06TKWLV0q4IkEqlZqm44LCEPfCn4vixRDh/ViQYGAF3wHeK8M9Hi/BCqyszKFTUFN0pOnTiE7cwZMDidCQ0NRVFom7REXFysydMVFxZg7b55iTRmVUpMXVDrpJsOykXicvGD1/NtkqvitQAf3tGqA7JPAEU/Aw3NbVQ1HWZYBFBadQ0VFCeyjA0hPTUXezNkIDYmA08sX3pYARIaTwWMVYMvpHARMwxgZHsDo8LCYZLe1tsnCiZ4lYtruZ4XTm+NjB2ZkzURgUAiF7GFiwnN0GL7+PhgfsaDpRiMqy86gpaUSc+bOQeGlKvRjCFeulcJq8UFocCwSYtPkmfUPdCAoiIsaC4IDwyURajLT0yYUba29gJcTNddrcOnSZUSGB2De3BkYGRzG9WutSJuWA7vTKdcWFxODz3buEtBldu4sNDY14XpdtcjncRyLiYxGZGQYAvz90NdHTf8RREQlICUlB3a7BUMjwLDdgWs1NRgdbEdTWzVW3rYENv9QXLnSjtq6TgwROB4ehGNsCMOOATBfbR8cAxwjiIr0w4zpqbhe04zi0msCCJq8RkD4z2L2g49vOEDGn1c3MtPT4e+XCKcpDF7+vrD6W2HzI0DBRDIlBCnVBJF+4qJo0OSQcT88NBLOcRNGhshoGEZTcxMsNlay0dSaVetB8LNYYZUF6CisNi4yKc80JnJy7EIWkR70ho8XEBwYKPNNa2srGhsb4Wu1ifQTE+RcLDGxLEAFpZ8MLVyRxBtzCjDC+ZNABxkVrMTn/GX2Hr8JqCBrQrEYBgSo0HOKi1HR1wc/f+UVwHeUbBh/gl5kxfXRo6JPjJRDQ5VHhVT7aaACTnhZvGC3OzA8OCqMCn582VcpJWTMCxy3mchnX5E5v6cHNoN5qXWNBTgQNoUbqFBAimKuaaBCiglMXBwraabJQIUAARKamUUiq4tARWiozKk0oSazyxOo0MUKZt6LoY8tjApD+onHr61rkDYkU4DvI4/PYg0mArr6uiYAFWRUELjndVD6aWR0RFh0PL+WcBD5L3hjbMQhoDULKwgKT/ao4IkkASLmq18AVDApwsU1K7NZacgKwdFRYVRwTA4K9IevxdfFqNDJOc+xT8lMmVBbXy+gmhuo8EYvfUI8GBW8N51AoXY1WY2M2whWa6CCYMQEoMKLlZuskCTT0AJKYwqYxqTLnwpU3DIkvjkbvHbjIszKm46qiuvYs+vEzXv9/xGoMOaqW68q/oO+nRKQmOr4/4dAhaci1xRJ35spFr/vXv8AoMLzXOx+roXbRBDgltX6xnpSJU/d0k+ejArPjKgbHpgkP/YfAFQsWLEA02ZMQ9GFIhRfLJR4Uy5v4oJyygabssknH0MfYQq/ENV+7gS5K0fAH6YAe2QJbVyAXg3LkzON42t/+R054yv/+1kkp6di6fqVaG1qweGP97qkW/T+UzEqNONl4s17XtA4nvjJ9+XPL//Dr5A8LQ1LN92GtoZmHP5ot9rNAJncexnP/BYsCs/70ZX/nKsWrV2B6bNm4NLJs7h08pyaU3QS1kMuyRWXGj/cZBpttFVKZgZW3L4eLfWN2PfuJzc/WwOoUPl948qN+UZ3c3e7uyvaOZcrKVx3jkgVrSoGhI6hGY/rYibO7eJ1wByFET8o4EIxN0Qay2TCYz95EhGxMdjx7Ou4XlFlMBJUX1W+AArI0ElnJqI5f2rTYwExODYZmCCva8sj9yA+NQmf79yHysJSI9GvlAP4EW9FwzdRP0vdGVWFvGZEGfdmfCecQII2LmBBSUi7QR4l2aSki1QnUXO+kqlijKjviftwX3V/zG2YFbtB2BFklTBRT7aE0cYuU3l15DufeABJGanY98EuVFwuUYAHZbeMc6v93W+A9vwQxofBEtBSWopxofJ9uuBEACeCHw4HfvOs8r/g58nv0Kia8bAChpiw1wbXwjIRdo5qQzJX2QeUgbknuORmiuh28lyHKXaNlvnWnhUuZSqXsouwVA0wQhUem5VMmOtcyuBdZLvIGJb7VOCMzldqppCSM3N7UsjxYFISUQImKW8OzYjh9YmPJBUjqHrAgVUMuxVD90ug4ubh58tv/pO3wM/vcgMVE5ItU2IVbpknd0DxRUCFCtDcyX022MTtb5aQmlzy4DkAKFBCURa1Z4IbpnAd2aNK9uZH5GFS5pmb/8L4xSOymcCS0EHkpAaTwcN1pROYiirXT913lRTT8YUGaOR7D2koqexV2eTf09uMa1AHMD78eVL73wJtUs/o5mejC17ULp4eFW4zbS5ItUcFDRpJb1NABaWfFLPCDVQMYc7ydTJZMwk7MDgobAFdRUENYqmG9FETBiUa6E3ApARlBGhwzKRDXFyCTA5kZNB8Mzg0HAnJyUp+YnxcTJJ1/7haWYmejnZER0chJjpWquE5cczIyxNgJSSUBqK+KsAHqxQUEk+UGiblZ6Guz63hqCZ7h0hS6apKVvyxuk+h5hIqiL46ExFSXWsyy3FZOamrM7o6usT0lvdBCqPNz4qw0CAM2+0Ii4iQCmdOZPbBEXS1t4vUQU9PFyoryiXxwqQUDXUpexQSEymJEd4DzZwpI0JdeU9gIjY2Rp4jzbY4ybP7Ce3Q0Ee0j46ht7cPI6MqKGCioLO9DaOOcYSERaCvpwc9Xe2Ii41GceFlzMqdg6GBAfGo6Opqw7HPD0vl5eIlSxAUGg6bnx+OHD6EwosXYR8aEEiOskbSI106sOpZK3kGysQoDWwm/VT1gZfcS0pKKnwD/BEeFYXElBTZhgk2Gmrv/Wy3yMUsX7lCgIqw8HDRi2T1hdBLWcUiwZhDklV8nwhUEGAQoMIvQJJGBAi8aEA6NoLK8lIE2Hxx4XyBmMLeefc9SEtPg4PvIaXFbDQuc4ipLI9FqaaY6GhJDrK/sj94W72lIp3PoK2lFa+//DL+6kc/QUY6GQFKqkwBc0p+RNgUZmB4jEnMRvT19gmT5cTxExKcUPff6u8nVFaprKZxd28fWpqbpD3j4mIQGRaO7s4uOMaUoZiXjw+CQynF4iMeLwJQ0YuFJqQGQ+tKWSmCrFZs2LQJJm+1OCCQ6BgZFcmviLh4FFeUiURUXlY2wgODRBfT6QX4U8bEyxvllVU4e+IkNqxaiZjYKDh8gNGhUZgsPmjv7kTxxQKsWLAQaSmpcJjH5T1j4Hru3DlJeCcYXhQMttk2BZcLxGQ+Koq+Hz5SrdLV1YOGpibkzJwpSUQGtcePHUNCQqIk6Wx+/rh0uVBANla38z6uXKnCkiVLxOtEfAL0QnRSVan0TY/qaNcIKt8ptpXnd56D8YRknaFhqo9FyRX9mQyQ0ANHaZ1Ss9+QaBHZr3pcvvw5mptrYYIX5uTNx4wZubD5Bcrvo+NeYOk7WSL+vn5SPe8YGxZ5F8eYkgrivMJjE4Rqb2tBTHQYfIO8MO5ll+eeEJ+GAF8ajBOYova8E5ZAmwT3o8NDqLlahrobVejqbMXsvDy0dzeirKJQ3qe21gE4HAp8DQy2ID0lCtOnpUmwvRDm8QAAIABJREFUzndyoH8IySlZaG3pwkB/M85dzJdnTVPzuLhEFBVVobfLjtx5c2D198HB/QfQ1NyA4f4+aYfFixZgZk4ewsKiUd/YgKNH83Gloloky1KnRSMlJRRW0vqdrEIPRmRkophlFxSVobGpFUP2TlgtXtiwbr14YZw9W4SyiusYcwCjI32wj1L+yYFxhxWDA3bY/MyYPj0as2dloG/QiZKqdkRGJCHQ5ou4mCgEh0dhDFbUXCtHV2sJVi5bgHGvCHQM2uRZiI8FpYn86O+iqvkI9g4ODImnwbBjRBLs9DlgPyI40N8/gMamRnnfVBwwjkA/G/xoiOxrkefoZyMg7hCWi32YRs6jYjxN7xu+E8EBoXLc1rY21NbWCbBHuTfN4lFgs1XGGZ2Ql0XkOOQ7JvFlzAGllqySIOa1dHV1is8LAXNGY2SNcbHd190v4xXvU5kpmjE4MCgsO19D+omJZY4ZTMar8/Sju7dHQEOC8wT0hf7OnmwYApINJtcyRpCkUwAOXgvHbS72eO28F4KojBt4zRwbfS1KKkIl4SmJpYyreV1ksfFeyGCkb4ZmKcp8yOOa1IKP1f7cntuwOIJ9THknqRiH7wMLCAiWsU0IdrW0tsorrRknEh2x6lOug/1BgRTCphD6vhn1TU2yiPb18kGgH+Up6VE1hpFRu7AOOfmxfcxOoKm+wQA5vNA70I3RsREBfrR/kIzrEmQoXWQyYMiqCLQFCFAhPibUITeqBVW1Kis+zSIZxnvj1WqdcjL3lGyBMVIxKUMJAqcDbe0tMvYGBirgnQkN+lRoPXB3lamqTPSCl3hUCCPI3/Co8DZLHGgXmQM15vFfravNAgt6h1Gijs+XBQgsRiCziPFeD/uj4VHB50uggr42jIf4TPi5SfrJrAA9neTyZG67x+uJVcxTBdh8nvc/shHRMWHo6e7HZ58cR3NTu2vzpOQYbNq2DF3tPdjxzoFJh5liMUVAaMp11q2vZCpVpqnz6bcuH7+Zxc7z/QmMii/O+P7Rq+OklDhs3LYaXR3d2PH2HiOXdHPa151oN6rI3audL17F/QHAw4RHMkX1vbqiL8h23+LOPSWNJqyAp0rge27ksc0XAxVGIthgg8lTNZKfHitC+fFWAkWTu+Pk37PzsrD29jWoLKnE/p0H3eCDy7sQuG3rasxeOBuXz13G53sOS9GWWjvyf9Wa2Hiwxs8Tywxv9YiS0pOx+d7b0dnWgR0vvTupdSc0jsfhJz4flSSfBJjc6jl5ABXqCDcDFdNzsrDh3q3o7uzGm8+8KFvpKnlhIqgFjfs2XT9OZha4IkNZL3K3b/zVU/LlS7/4d0zPy8GmB7aju6MTb/zrc642lN7HNZsBTLkGbgOlcp3aszENiSKOfevu3oq5yxfh4omzOPThpxMT5B5gjeu4LiaBHiMmsnWmz56JrY/eKxLLvG5+JmeFFD7h0rMy2sik5hLDkFqbiotiA/MeUuVPk2JDYom+GvI3lUTWAIT2UtDJdplbxXtQyR7p7bV3A+edrz39FCJio/HBs6+juqRcFUoakjwK6FDJeu0toNgWKlbTSXXXczYULx754bcEADr44Wc4uZd9X0noCkPFACoYY2igxRNIM7qnMTfrNYdmR5gkj6DuR/luKFaEWke7WCgCNqn20YlxbsdrYDGAqzjRiFe4jZBBmOgWOSWjaFEelpJzUvGVMdqNj+PrP30K2XNzsPutj3H4k32qYNVgROjkvEh5SVu52Qm8LuYdGLsIEGGACYolwEIVVRjHD0EIxgvPvUh5WvX53ncUG4Q5FOZPjEtUviFsD64HDPk78e4QE3HFMGGbiQSxXcUfAmII+8TNjNDPV5ilYmTtVnsxXisXUMH1qTB8XH4nCtxgP1XG2p791wGzNyVIWYBBeSvF5uU2XAMzxuVHMS7Ioudx3B52uv9psEK/0vxXwBEv1ccEOGE/9I5Z+MfNTLcYBL/86ssW+L+pBX5xJ6WfPK/oFrOr3mASMCDBvkYRXW+Psb9OAv2Rgbh72tY/TQWCTIriPAEHDyBBXfKtLkK7/ajzTET1PRNSRqzhGV9N8QAVuKA2lKBDmCHqOxdUoJNe+niuEUWFcK6P4AtuMEYd04PzIG2vJiR1/VorcaIkKI+hcQsFRXiCFhqwUaGvYqxMxDj0AG1g627ap8ujYtww06YuIBkVyvhagArtUSFAxZDBqHADFcJaIFBhGDuriUIt+Gn4yGvlIN4/0CfMi9CgIDFwZlI4Pj5REj0EKZjEoPFqeGSUSDlxEqL3gExOPj6oKC9Fd0cboqOiEBsTi3FqO46PY9qMGbA7xhAeGSqJF+WnREkBNaEzweEcVx4KurqC16gqGs3i08EEjpab0EAF96UsB40j9WsxMEDzahpUU3fZR2iLTJK3NrfI/TJ5ywn0WvUVmMdHERAUJLJHTK6LadbQKLo6OmUBT6Ciqqpcjs8Ke3//IKmaD4pSlecspCD4Y/MPlGQ/Ezwi8TE6KowKXi9/d2lTCkFAgWBM7JOpYh+jVBJlpHzQ1dEOh9OEoJAw9PX2oKezHfGxUSgvLUFW9iwM9vdJBWZzYwNO5h9DZEQEFi9ahAG7HadP5ON6dTWkvJi0U9M4vJnQsbi1IFlhLMk9VhFIUoedkMEl2S1W8oMlkcZtwqJjMHPOXCSmpig6pbePSIft/WyPAFFLly9BfGKSABXcn4CLfnaiAWkAFbxfVv7yGbAf+tmCpD0pf+RtdmLcMYrysmKRODp//iJYrHDPffcjJS1V5DFg9hJmA4MKyn8xOUcZJsqOUdqDvzPJ4uPnI0AFE1oEKl576RX87McGUDHuFKNZJeOiqnoVUGHCoL0fN+pqJZhhcurkyZPSr1NSeN+K1SPJvnGTUVVtl8rf8NAQYYF406jdbhd/h46eLvj62+Dn64OhQaXDPs6/O8aEScKE1tWycgEqNm7aKJ4CDCLpJTI6NIyIiCiEx8WgiEBFaSnyMjMR5h8k+uFObxP8rRaMeXmhouKKmGlvWL0a4RGhsJtGYXKaYbJY0NrZivLCYty2eAlSkhJBKEpVmTgVUJGYKFJNOlgkTaawuBgxMTECLhKY4bvU3dMnWvzZM3IkQOZzPHXqlBhxa0+V8rIqSdiyPZnkqqmpweLFiwU0HBikNr0aaVX1jPpZQAUjaNWLEZ3MUu+GdMopp25PoOJmeaeptQbGx9knCZDx6Aoga2yow5kzp9DTWycV9osWLkF8XDKsFlZTM0FpwSgDZJikvwUFBAhgRb1VSbBKsM4xS71P3mYzKqtKcfb0cfj4OpGQHAmbLQChQZGIjoyHnyUYoyMOjIyOw9ufiWrGvmMoLbmM2NhIFJw7A7t9ADkzM9HaVifjYkBANJob+1Bz/Tqa2+thhh1hwYGIjY8SEC4yMgZhobG4ca0OZ88exvBIN9LSUzFv4SIM9Nlx/nwphofGEZ8Uj5KKQhReLkB8QpywybZt3YRdn3yC+QsWITExHcEhweju7Mfez47g4uUC2J2diIqyITsjE8lJKUKVpp+E2WxBZ08vKqqq0dJ+QxLlyYmpWLJ0JS5cLMHx/IuAyQJfqxk2fyvCI6IRHZmAyIgYdHfWY3CgHqmpMYiKS8eQkx45frD3D8i76xsQgFF4obqqCF3NhVi9YgEc5gi0Ddpgd3Dh4wV/P7Iq6G+gEuRDgyMyv1H7n3I5lO+hfBA/HHsJFDQ0NMp8IEjTuFNAJybfbQTOnaPwtXljzD4ML1gw2D8sIK7JaxzevnyuZLCEKaCitRU3btyQ/pCWRtN0NZ5z7Oc4IUAFJYPE00ElZzmniqSTUWHI+yQ4wE93T7ckgLmoZCTDcYrv00APAQv6ONnEZ8YTqLDa/OS+yZ5iwp3/8dis9O+m7xGLAkLIOvGVBRaTEyK9xMUdjQCHhmSh1t3V4wFUEGjmfPr7gArIOCbjqKGN7COyUmYBVDRQIWw6MdNmJRrNHQlUWGTMFV8oSgMG2GR+l7dIQG6C8BOBCrY371UbWWpQkvObABUGm0L7X3AurW1olPbw87LA3+or8xm1iwlU9A32y3hIMEQDFQQ4eB0DQ70ia0lGBZ8J25zPSiU/TOJt0tnRLnNZoJ+/+PPQS4L7K8cIlexQsg+KUSExqZMJDmWIKf+KZrMB1jq0xvUY2jta5PvAQJuKL8ZVm2hTSxlLjQQJkx1eMIv0E0EOf39fwxPKZAAVvIaJHhUq3rPA7E2GYJcA5PTxIPDM+Z/Ppbuz4/cDFT3eIpvmTcksAlYiw+ENL0noKQ1p/dFVsvx9qty1JyiQk5uB1esXCABLpuTZ/CKcO13sOl5SSiw2TgVUTJFwnnIy+VP+8Ack4D0P6wLMPYuiPLP/N13DVKmPL07YSyJIF5VNPqY7++N6CAJU3HGbAireMirIvwAQcFWoT859f9GDNa5jwmMxbu8mIGiqKX8KxEgnYyfvplppYrGTjNHM22pD2cntM6mQwvVnj2c98R50UeDEA6nNjRWelhB25Yw9YhOPRzzVbefMzsYaA6g48MnBiS+PJOfcbA4x5yXMPamtXMfWmUbj+eq1qmfVvm4CAhVb7t0mQMUHL70z4QZpGO5uG48wzaOqW8slqdrBPyAp4XFMdXQnHv+RYlS8+i/P/gEYlQcrQNbVE+VGJeZUgaeRtHR7E3z9J9+T87z0j782Crgmgqkys0sF9UTzZtXl3fGsbhP9HdcN7n6gHp0Ay9IPPdvQ+Flka1i5rsZrJojFG8jbYBuwcE88E1TCVpQHOG96fKeT9GQ8KjlK5WGgYw637+jUuJ+OrfW26rZVop7zDosOGDfIeshYU0hsb/gZMCZgkljkNA3pIwIaX3v6+4iMU4yKG1XXXAljDZ7rCnZRT2A7eKtEsgYqPAF6BbpTLndMYihd3Chzo5mSTAY44QIQ3SxrHkfWv6y7MRjfUqxlMCJU4luBWNqLQq/dtQSkyAgZcpUqea4T7QqkYIfRBZU8DuNSAv0K7FGeisKElniCyXK1xpSfGQuIFJgav1j4otmkQyMsjlIFJ1wzKo8PN5tDZ6x4LH5EthMqQa/GPwPyJZggcsMEDyhz5St96Ze/co9P3/supSuNAhLmZAzjbRZZ8C1ifKvfMy39pYEZxUZRzASRrxwblX3IQtA5HZ5br8X5syogVvKcvB62qRS4GNJhPAfXlIz1xkbZv5U0mYqveY9KuWPMqTxR2Nb8l2oaumiV0l28NiULPi4xMuMUu31YPWtjnJA2Zx8yXuqJ0707ayfv4JdAxZ8SQX25z//NLSBAhWvWnOpKbxF26XeDo+vkDLtrAv4j7nzK2GESUOGR2Hcd3UBR3cmiCajFJDkkHbTpyHTSifUI8IcEM5Nuz3MXNfzemhly62omBSHoj/pJ/a+OMyd4gRiMDVdgohdhUiGtFpuuxJquhjAOPuHWmJV0neXmh3BTc7sKIrSZtgFUkFUh1YEOScJPACpopk3QQhgWw8Ko4ITHSYQTJidZHeiQpSAJAKuh4zc6gu5uGizaER4aKlIE/JnVqlzAUmZDErxOCPuA0hBc3ApaLhROb1RWVKCns0MS2QQqWInMyr7EtDRhggQEUbJJ6S+zSpWTAgMLMfwdVzRGVV3B6gMlnyCLbZNREW8ECH42X9h8baqCQuZlpyD4TPIwKcAEDQMlSmBpySdWlVKuJjoySiZqGuLWVFciNiEe0XFxUo3LQMEx7BA5Jy7gNVBBGYXpAlQEIjk5BUHRETJZUnOcz16BFG6ggm3Cil6tdSnJGg9wiIEDtSZ7Kf1EORAvsyQm2HZjDgIVlArqRXdnG+KjI0UaKTUtA/ahEZFTqaosR9HlAsTFREviOT8/HwM9PdJOVm8T/Hx84GeljrQPSzuNgIb9h/9xQaPalQlwymPoBDEZFSrwNGGI1R0WKxJTU5GeOR0hoeES3OzbvRfRUZFYMgVQod8j9js+By0jxOQOE302/2AXUOHjxTfRgfKSIvjbfHH2zHlJ4jzw0CNISkl2AxU2myzCCAoRmKDMDg0/CSaxb1JL28fP4gIq2lvb8PpLL+OnP34aGWn0umACULEtNNgl764Z6B7oQX1DvVwr/0aggoEPPUHGjL4oz3FoWBJ9DI4ps0H5GCbc7QNDkuhhor9voF8AOT8b5ZMYEDrk/RketUvCmtXMtVVXEOzriw2bNoqZKqufydSwDw4hPiEBYTGxKK4sQwXlvqZnIcw/kIp1GDU5Eexvw6jZjPLyKpw/eRpb1q1FcGgAugd74c/KYasvGtuaUFlUguVz5yEpMRG0Y5X8BUw4c+YMklNShFEhVSmG/lZhcZGAF7Ex8S4fIzIqKA+SOWOGogybTOJBweSsJEDNXigvrxSGBQEemjSXl5dj3rx5alwaMuSsPOSdXMwHGTcVgKEWDwqgUOPl1ECFJ0ghb71xXe7vpwYqCDQRpBgbG8LgYA+qr1agpKQQo45hkRHLzs7BterrIqsUG5uImOg4+DEZ7qOqpVk9TZ8WHy9WgCkpm3GzpESEbSA6sGIaOI7Wlgbk5x9GbUM1QkNCkBCfiOjIGESEhiMwIBh0NLYGhmJcqqwIPNahs6NNAK7Pdu3EypXLERsXrhLVtnD4B0TLu3P0+CHxl2huqZcxj0a4KSnJSEpKQUN9A5rqq5GUGI1ZuXkICAhGW0cPCi+Xw+zlJ34q125cEaBz1qyZaGpsEHk/Jq17u3vlOXDcpXfB2KgPHKMEgHvR3dcML+8AMY4PDQ1DVES4MBFMlPPx8UZdS534MpBRFh+fgmmZuejstcNsCcDwIDVqR2Hz80WAfwgcI3bcqC5EU0MxMrNTERY3HUNjQYA5CH3tXZBxPSgYw6MOVJcXoKe1GKtXLoDTKxKtA36wjzHhboa/n6+cjws/WQwOKG8QYbA5FJBIdpSugNNAhY8hgaakcvyMcZKG9k7Y/C1iZMwq9eGBYVkogawvK5PyvggJCpM5lN5GBCo4l/Bd0ItWjhHsAxxn+C/nODWfjbuACv3OeQIVHL/IkCCIwvFGAxU0buZCSjMqeEw3o4LjIQSo4HhEUILH5rG6erpl0cv5h+OULPbpoWIYgxOQZ3twwUegnPUXPAbH9jEHK+huDVRwPnGxh0QSi5q/ar7QQIWWjlReUYZsFdtRfDAUUME+TeCG2/gH+ItesydQQVBb5IjotzMyKuMKz6ETBXq8sHgrNocGkjVQQRCCQAXbw+ZjhVUS6F4YdY5hzOlE/9CAXA/PoYEKGYfMJgzbBwSoCAoKluvnuZR/A3WvCSo70dnRIUUE/n70yfKHlUkbJhqMZIeq4FPSAyw+EJYOlQIMoELpdSuzUBkPPYCK1rZmiRM0UMFnzGepEza6/0i/ZoHDnwhUePkoM20mMwL8bBLH+flaVUFKR/vvByq6vYW5yiTIZDPt/1OgYsv2FUifloSCC+XImzMdjQ1t+OR9VTG7fstSzJo9zRW7sz+eP12CU8cvqe/MJoRHhGD7PbdJe+/84DC6OnvlTxu2LkPWjFScyS8U4GPewhzMW5QD/wA/afPmxnYcO3weTQ1tmDEzHWs2LhYmR2RUqPT1I/vP4GplLdZuXoz06UlSNcrYtb62GccOnkNHu5JRm/xhUmrd5qVIn55sVJqOorLsmuyjKj6B7JnpWLx8NoJDA+VZE6S5eLYYF8+WuA6XNy8L8xflIihEAZwD/YPGNgrEmQxU8PrWbl4+8byl1Th28DRWrV+CWXOyJrbjqUKcOnb+puuftygX8xbnCqjIduru7MGJI2dxtfK6Ubw/jlVrlyAnN1PGb27T2tyO44dOo+5GoxwvKTkOy9csRlRshErEDo+gtLASx/afwozc6VizZQWaG1qx441PXed/7MkH5OdXf6eq+vPmz8SCJbMRFBLouv8Lpy6h4Eyh/B4eGYZVG5chITlOQGKuKSpLr+Lo/nw5Xw4ZCltWoaG2CRHR4QgIpK+PE3XX61FWVIlFK+YjNDxEjkXw5tiBfNRUXcfS2xZj4fJ5KCuswMFdqh8mpiZg090b0NnWiR2vfaSub2EuFiybh6CQIHV9fQO4cKoABacvGcXtE4EKxvvrtq1BRla6S96vorgSx/Ydxx0PbUNyWpKrLThWHv70MMoul6nvjIXqhrs2YsbsGTh3/BxOHjqB+75+P2ITYnHo04MovVQikdSytSswb9l8XDx5QbYJDA7EmtvXI2VaqiHvMoa667U4svswFixbiNz5eRP6xbljp2W/GXNmYvFtSxESHqr6aG8/Lpw4i4snzk3pGRMeE4nV29YhITVJxkPeR3VpFQ59vE+04dkwienJWLl1DaLiyUAHWhuaQQYyY+dX/uV3yJmXi3V3bUZTXQPef/ZNuafw6Ejctn0DEtKSXce9WlKJQx/uFfDVBQ7qOzGZkJSRgtW3r0NUgjpPS32TzLtcC774D7/GzAV5WH/P7Wi6UY93f/uqbDN9VjZWbVuP0EiyM7lPowDYvLYXfv5LrNiyDkvWr8S18ityTdyOSfva6uvYv+NTtDe3YutDd2HWgjk4eeAoju85LMUgG+7bhrTsaa72r71Sg/3v7UR7U4tc09q7t2LG/DzFsnQ60VzXiEM7PkPd1RrMWjQXGx+6Ew3XavH6v/4OeUvmiwwSjxGdEIfAkCCZp6+XX0Hx2QKs2LoOYdGRcv0dza048P5OXCkulz5E8GDjg3cieXq6JJ8pcVxxqRi73/hAGKoc97LmzsLq7RsRFRer5siBQVw+dR573vrItYbQcRZjsfCYKGz76r1IzZ4m+3e0tMHOCvegQMWoKKvED//hvwlL/oNnX5Pfuf+dTzyM3MXz8Olr74lEVnhMNLY8fDfSZkwX/y/KFJZdKMLHL78tuYkn/uopJKSl4MMX30ThqQv45l//GaLiY9HW2IykaWlyP309vTj+2SFExkZj9tL5sPha5Vp4/Tuef0P6yY//9W+lnd/77auoLquSeePebz2KvKXz8cnL7+Dc56eQsyAPmx/YjpjEeGmDof5BXDh+Gp+88p6xjlEdTRem8Lg8xvyVS+ScLESrvXodKZlpOPbZIex++0P89Jn/JZLGb//6ZZRdKpZ++JUffBNzly/EB8+/iVMHT+CHf/80Uqan4a1fv4ozR04IiKHMnVUBDuNvzfAQcEP8KlQBh3iMsBBKfCxUzkhl4xXoJIAGk/n2USnieP4lN6PiO99S85IwX1jW5QLBDTaImIWz0E8pNMjaTQyulbyVlt/Snp8sWFGsFMXG4LvP65I8jYP+o8oDgtupNfOwzCWKAaHiJMZNjMN4TH0vSmJLAXdch3E7PneVXyEYY5djMsZVnhYa1OSaU+lNMOZlDoTJAF6LsFuFSaPBSI9cncvDljkV55dAhWum+PKH/zIt8Is7sz3u5QsqDW5VFSS5mymAChknjJ2mrPYxTu2ZOb/lJegkkUb6J4EXBlChTqn/5vkiTzqo/DpVhdAUj/YLizA8AAZ9ywLH6iBwImgwGY646WqMe9BotKqcuJlNofbTjArjHBNuS0np6I9LvsmzqOQWnhZqNuCOugrEqEiTrwwEfIKZtlP0BJn4FqBCpJ/4nwImBm4BVHByEKBiiHrhrIZVppdKM5G5aEO2YXgQHZ3t8lzDgoMlIFSV8P0iecTEJKV3xHTY6iuJdTENJXggCUeg5to19PV0iyxPTEws6FFBoCI6MVGSfVY/6nj7SAKQiX2r4SUhSSFqjXswKjT9TlVuUtZi0JBugSSpPaWfKNfQ1z+ojIMFEFIGSoqpQACBGtwqWRMRFiGTVk93ByrKChEcForI6BhpVwIVzhGVjBBGRW+XgAL20RFkZExHgL+SfgqNjZKAYGTIDl8/m3FPNklq8LycVFnRy4mYba0BIj5nqU6RqgiHaIqTiaAAIx/0dnXBPkbpp3ABKno62xATGY7r12uQmJSM0ZERkYe6drUS1ZWVYijK73q7O+DjbUZYUKAksymjYrP6SIU3kzMqcFftIkbqdHHlbwSCvL2kUpqV9P0Dg/AXCSsrhsecaO/tQ3tPL0IiI5E7Zw78/IOwd/deREZGYPHypUhIIqMiQt5wGp/qxDElazRQwXvV0k8aqKDMmBerbH0ICTpQXlosUlynT50ToOLBhx9BQnKSctAxGBVsOwIVTMYRiGBb8xkx6SX92AAqxOujvR1vvETpp6cxLSNDggrNttCMCgVUmNDW3SZyLqwAZiXP8eMnJIhjEpLBD58dzzXUT519RWelpEpwcKCAagFWP/T39CI5OVnk1VjN7cVKbB9VdTw0NCJ9X/T0zSbUX6tBqJ8v1m/cgDHx3RgRoGKgpxfpGRkIjY5BSVUFKirLkTctEyG2AL4acJjGEcAFnLc3ysorceHkGWzbuEGqTpu7WhEeEg5vPz/UN9fjSmk5ls2Zh2QyKkxOAeE4nhDQysjIEPaHAs6UUUhhUSFi4+IQGxNn9BO++93o6OxEVma2UWFklv0pycW24v6VV64K8BEVGSkyZoWFhcjKzpLAs39AARW64lzPGZKc82BUeLIq1JwyUXZv8qJzMljhug+1VHCNwZO385JE4Si6u9tw+dJZ1NyoQoC/BVnZ05GVPRd+vgECdhKsaKhvEkYFDcYjYyNgC6CnQAAiQsPgbfYRwE9AW5NTGeI6zZK4Y0UxAayxMcq9DePSpbM4ffo0enu7xbh6ZvZ0RMdEI5gGyEERhpRZh7zrnMMimAQAcPb0eczIyRBwICQ0Bv7+kTL+FZdeRGRUFBoaG9De0YbCwksSaIeEKAPs0AArUlOSMDAwBJstEC2tnWhrZ9W8SRKwo84RtWgZHUVfX7ckWrlwYCJbvBtYUW/2RaBvJIbo7TDQhZS0RCSlz4KPxRdXq6/i6pVKjA33IzTYhtiocFiD/ARsY5/IzMpFaEQ8hkbNGLQD/b30BSCLyhdWbz84R4bQcL0Yba3lyMnLRnjcNHQN+cNkDkJ/R5eMAf6hoRixj6Gq+Cz628uwauXvwqHYAAAgAElEQVR8OL0j0drvB/uoCd4WMwIo/WRjNb4GKoakfTRQwUQ8WQa6DyigosElxcNnFGizie8CE7SsTgsIYJLNifFRjqmjMm5zKvHiOOoBVNAzoba2dmqgol8BFbKokkpKN1ChKwg1UMG+z/GLjDE+B85BHEN43UP9KlGgwW4BKgYHZfwja4sfgrZM9oeGhMriirJQZFQwuU2pMno98Fj0qOC/ZFaQGs/jcCHX081+p4ylmXTlPOoCKmxKcooxA89po0SWUZGsF8y8fvGJ4HENjWsC0pyHufjnApB9g2OMABWs5jebBSiRJHkgWTEqcOJ8wbGW4ItibPnK3EigQlff6TGE7eJDD4VJQIWAGWYzbtQ3yLUGWPzA2kUtcceXq2egXxbwYqbtBBrr6g2wlO/IMEbGhl1AhYAwIstIdgOkX7KIgRJb/lY/YVT4WqziLSSVg3IvCqjgflZfVRFLoEIbihKkUGaQaqjiNWiQsKWVklWG9JPFR+ZnPkuJPw3pAw2MeQIVnIfol0TwhQA5WbUEVbQ0l65+5XF8LJQoNBgVIyPCLGIFLOXU6M3SQcDUTxUvUB6UptqsCKXfCcEjfhxdBGH+44GK0LAg3Hn/WjnHrh2fY/Mdy8U4fv+n+ai93oSY2AjEJkRi4ZJZ6O7qRWFBJdpa6KXUbTSm6ktbt69ESlo8jh46h9Kiq1Kw8eBjW+SZ7P74KKJiw7F89TwMD42g6FIleF6CBS1N7fj4vUPImJ4kQAXbr7W5A+2tXXKchUtzkZoRj/raFlSUVCMlPR5p05LQUNeCTz887AIePFc2m7atQOaMNNmGnhvZOemIiYvA5QvlOHborPxt7aal8nwLL5bLMXLnZolvTP7nF1BUUIHU9ARsuH2l9I2CcyXyPuTNy5ZCnsP7TklCXrMXdXHWpm2rkJmTjobaZlRV1CB7ZgZi4iJx+XwpKsuqERsfjYXLZqt2vFiGtuYOdLR3Tkjyzl04C8tvW4i+3n4UnCuWRP7MvEwBUj55fy+6Onqw7LYFmLcoT5L7RQVliIwOR/bMaXLczz46KEDklrvWIzgkEOUlV+Q8ufNmICw8BOdPXkJPV+/vBSpSM5Kw8Y41cm0FZ4skTiNwIfe/54QACnc9cjui4yJRVlSFlqYWzMzLRlRsJC6cvozjB/Ixa04O1mxZKePDlbKraKxrAlkL0XEsXHKgpakVFcVVSEpNQHpWGprqm/Heyx9OACoO7FRARVLaRKAidVoKNt61XpJoF09fkucze2GurD+O7P4cBCBcjBSjc2y+eyOyZmWiobYBVSVXQKmnmPgYXDpzGTVVNYhLjsWC5QvkZ15vw40GiTOFCm9o9m+4exJQ8cT9iE2MxaFdB1F2SYFcy9YZQEX+eZw6dAJbHrgDmbOyca2yGtXlVzBtZiZSMlJRU1WN00dOIi4pHotWL0F3Rzcuny1AW2MLImOjsOaODRJDXj5dIAnt3MVzJKmev/coCs9cvGmZz/Xhfd9+RJLEV0urcL2yGtlzZiI+NREVl0ux971PERoZhm2P3o2wyHBUFZWj4Xo98hbPQWRcNDpa2icCFbUNeP+5N2QsfuC7j8k2V0sqUMPjzp0lYEj5pRLsfWenodtvMB5gkuNvf/xehEVFoLKwDPU1tZi9ZJ6AI0ykv/gPv8LMBbNdQMU7v3kFkTFR2P61BxAaEYbKy6Wou3YDc5YtkGR4R3Mbnv/7f8PKrQQqVsk8f73yqgAWOfPzEJucIMnwve/tVEDFwjk4deAYju85hDsffwDZc2bhamklrhSVIWv2TEnq8/f3fv2ygBSL1q1A4/V6SdinZqYje16uADiv/+9nkTVnJjY/fBcaaurw1jPPy3UTqOB4XV5QjPrq68hdMh9xKYmyXmm8UY/isxcFGMmcPQv1167jlX/8lczHX/3R9xCdGIeKgmJUl1Zg1uJ54tVRfK4AO196B+HRUXjwqScQEByEc0fyMdQ3gPm3LUVQWAiOfLwH+XuOGHOTMjbmPPbYj76L1BnTcK20CqUXCgVYSc3KENDgw+ffRFVRGf7in/8GVj8/YVhUl1VMACp2vfYeyi4U4uEfflP2K7tYJMDK7KULBFC5fPIcPn7pLTz+k++Lf8NHL72FS/nnBKjImJkl/fXckRMIiQjDvJVLhEFIoIBtyfdn8bqV8A8MELDgxJ4jePqXfyf9+N3fvILq0kqJIe/51iNyvp2vvCcMkMd//F0BgPL3fY7BvgEBp3j8gzs+xaGP9hgsDGUOzjlm/b3bcNv2jehobcOp/celny+8bakkzQ9+tBt73/0YP/v3n8t5X3/meVwtrhRA4MEnH5M+tuOFt3HmSD6+/z9/JEDFe8+9IYCJrIWMwi8dizGeV0Q6zQYximcNUMIzT6cM0pXkFEENLbvEY/7qd+5115PfZXEFVRS8XOCHknU05FENSTCyKPU1ecozSTznUEAJmbNWX4vBNuG6SXnBSTzK/Qk0OMbg460KwPg7izsYc2gWhioIVtcsrAyDccMCFGE8sejO20vyNDpG1FJYfCa8NsaWzHEw78V3RZgfTsoT0/NDsZ8JtPCe3B93Uk8XJfMRUEFBYs0vGRWeoc6XP/9XaIGfb3cDFVOTCDyy3WrNo8SMXFX7k4CDSQ3zRZDAhPy/Sy7KTWVSh5qEEkwqUNVmRvq07uu6BfrourabKZJ64aUHlQm38YVAhevMHrtMddceoMXke/OkyHowImTQ1Qixx6k8dVJvCdAYyTUXXjSxsY2zT/HsDP1LTQl1O1i4gQoCKEz+MsFOGRkmGdxABaWf1H/9gwQs3IyKuSvWG9rPilGhPB28FC3QYFR4eSvtxYEBykZ0SWKEVYL0SGhrbUV0TJxR8TMmiyiRVbKp6nP2F0XXVAh0fV2daPPHRMcoRgXR6fFxRCUkYJzJCj8mKrwMI1SLS2dQEtycOHT1oMhAUBKJyD8nGhptDrneA5vNV00+pPaZldQCDUuZ+GdSQEAQX6vhveAj++nJJSQwWCa7wYFe1N24IqquEdEEHlh5SmNdVtc1iSlyf38PKirKhAGQkT7NkH5SQAWT3wQqqBHOdmDFtQYqeO2saGVQzevS2ojUtVeTJGUy6FHR6wIqWAkw0Nvj8qgY6O9DV0crIkKC0NLShKiYWDHTbmtuQm9nB8qKCtHS2ACTcwy+ZiAqPBgxkZEIDfKHlQkc0clmhQGr+83CYGFgwEDBKka0PkqqTOQzrJLA4LPlBE9JJV+bP/qGhlBRcx3VdXWwBAQhMzsHp06fFU+PeYsXISUt3eVRMWboTUpCxUiqiBGVySSAFxNy7H9W3wAXo8LPSvEKByrLSiQwOXnilPhk3P/gQ4hPTICTUlTsLzZfGZoIVLAfNzU0iT8HwSp6VLA9LTaLMFR4X53tHXjjlVfx9F/8CJlZmXI9TLZx8SQVoNpYzGxGS2cLOru6JDnG72k4zeeWnk4mhg5qzAImjAwMir8GEzb+gTap7A4JCEJXW4fo1RMMkaDLahbjbx6HTIrBkWFpdyay6qqrEWz1xboN60W7nfI+A3396GhpxaxZuQiKjETplUqUV5RhXnYOgqx+kgx3mAFfSsr4+aGkrBIFp89g05o1AlQ0dTZLxb6PzYbGlkZcLavA4tw88aMgo0KI6E4nDh48iJkzZyIuLk4xZ0RI2ISLlwoEaImPo/m2mm86Orqkwpb9XgdpBCqmTyezyF8Sc1eqq5GcmiIyZ9ymoqICkZGRIisyPOIOqvX+euzkmVUiTFVku76/hfSTDsgnzjmeQLnSHFXSfG7vi8kxg9lBVlYvCgsvori4ADExYcjNy0ZCQjwsllAql7pATpovNzY2obmlRYyvQ8KChTGTnpKK4KBApTHLcZsMDZoIOs3w9fUHhdOYmJeEvxfQ1taCC+fPoLGxDk3NdUhLjkdiUryqxPYLkvGPfZKJ5v6ePoSFhYo58o3rDThx/CAWLVmIgED650RgcLAfhcUXEBgULONcYFAgLlw8JyAITBzFHBgf1UAE2WFm0MeIslRMmBCs5UKJIKSAb75WuScmWwf7h0QGCyY70tNSkTtjHlqb2nHhfD4efvQBRMRmw9vqj87eXhw7ehRnT53Ajavl8LOYEB4XJsbQ0VHRCAoMQUR0PPwDw2GxBWNggIyhEak4Nzm8pMK94UYp2lsrMXN2FgIiktFrZ4VsAPo6uhAc5A/foGCRwyu/fBJDXZVYtXw+HN4RaOnzxZiDEjNAoD+BCia5lX4upZ8ILNC42u5UMoeU9pEKKS+VmL9x4zp8ON6YxsVrJ5jjh5USUgpgCgj0EwCNcm4cZ5kw7xsYRGBIGIKCw8VYnWM5jbQJVBAIoDwc+wH7sK68V+xDZRytkstK+onXMJlRwW0ILtC4mduSmygeSuPjwupQVflWma8FvCAA2N8vC1w9pvFd1IwKHqunt0/eTc4//F4kOcdUfyVQweQ3nz9BuY72dphNNPemB5BT9uN8S4CdLDFW2mmgQjMq1AJTMSpYqCDvsSElSABMM+e09JMAFSblg8S+LrFG/4D0CzKCtB0Y75n3yfvjuEn5CoLfBLkFmKAnlKFZLec35lJ+r8EEXTRBRgUXyME2f4DjmbE4Z5KvZ6BX2o7t5j1uQl1trbSLt8UbI/YhASpEDskw05YiAotF4gN6ZvR0d4t/VwCLLWw2MWSXCkdKQIj2NmNhBVQQrJbfncqLiPMrYwPNqOAYRaBC9VMzGpuUCTgZFawiZfwjcZ/WYjf0lWVsozY1zLh+44a0L8EF6jJzCO0nEGWMURpMYrzC4xBAMnlZRMqT8ylZN5SvIlDB3yltpYAKVXXI+JBVxDTTlnZgLPr/EVAxf/FMLF2Rhxs1Tdi54wjWbloMSkEVnC9D/ucFcttfKP1kgF6z52Vhxaq5qCy/jgO7T2J6dgrWbVoiYAGP+/Djt4tf2pEDZ1FRek2OS4AkPjEaRw+ek2QJgQqyJT55/5D8PSsnTb4jKPLxuwddoMSd96+TayKr48IZt0QV98nITMb6LcvQ1zuA99/cA/vIqEj2bb1rtez/7qufYsudq5GYHIv8oxdx6XypcS4yOpagp7sPb728E0tXzsWCpbkoK7qCg3uUufj8xbmYnp2G0qIqFF4oNRJGKmGVkZmC9VtWCMDw/uufClgYFx+NrXevVed9ZaeAFpOln1Qy3b2e2nrXOiSmxOH44TMCAPBz31e2ISY2Eof35eNqRQ0e+tpdwhQhKNHU0CLbbLh9NbJmTsPpY+elH89fMhtlhZU4vPu4eoap8dh45xqp2r50pkiAiiZhVOxyTduPP/mg/Pzqb9/F0tULsHD5XDnGgU8/l+8XLJ2D6TPSUXq5Av19A7ht0wq0t3Xik7d3S1FZzuwsrNm8Sq5px+ufCCixZtMKXK+uxafvKU+O6TnTsO7226Rg4OO3dgnYQjDmrkfukHHts/f3Ii0z1cWoIFDBsSQxNR6b7tkojIoPXv0Iy9YswcIV81FWWI79lGmCCQtXzMP0GdNQcqkMl88VTSjYmzYjAxu2r0Nvdx/ee+l92IftAjDc/sBWWae8/dy7yJiRjnXb1qKyuBL7P97vahcmGf8QoKK8QAEVSwlULJ+PiwZQ8fiffVOqvPd98CluXKuVYojVt6+VJN3ONz6CeFTcr6SfdryopJ/ueuw+JKYnCShRkK9YN9kEfu7ciB7xjnjZdX36ByZmF69fjuqyK/jszY/la47/D3z3KwgKDcbBD/cgODQESzeuFJbFp2+QmTKOsOgI3P3EgzLvvPzPvxVGxfq7t6CptgHvPfsGFq9dLoliVr/ven2HAL4+VgseeepxBIWG4MCO3QJYeH4WrVmG5ZtWCxiw87UP5Dxke9z7jUfkvl/4hQIqNtyrGBXv/PplYSIsXrtCkuQ7X31X3q+ImCjc+62vyD7P/71iVCzdsAo1FVfx/rOvqXeXQMKDd6G5vhFv/+pFbH34HgOoOIoTnx3CN//mz2UMJnPgekW13O+6e7fJMT987g089INvIC41Cfvf/QSXT7Ktx3H3Nx+V5PqhD3cjIiYSWx69Bw01tXj7mReQQ6Di4Xskyf7e716R/jlz4VzxsWCC/s1fPicG4dHxsZL85/y/49nXkJo9Hau2bRAQ5oPfKQYJr+vxp59CcHgodr/+gSSEt37lPjRcu4E3//U5aQOyHhasXSHMi5O7D6n5QKrrvZCzcA7ueOw+NNc3yfb0tgoJDcGjf/ltKQj86IW3pD3/7B//GmTNkGFxTRgVZmx/4kHkLZ6PT155R+K6bV+9T9r1lX/6lVqT+vvj2//jLyVuffOZF7Dx/jsEVOGzuXj8DL7xsx8KQPTRi2+h5BxZTON4/EdPCiPk5N4j+OzND+Uetz56D5ZtvA1nD5/AjhfedAEVfOa8Np6bbIjZy8ioeE/a/84nHhLGym/+xz9LLDJn+QKs3Lpe2mD/+7tcbcBtucb+i3/678I8eue3r6Dqkip0vOtrD2LZxtU4sms/9rzzsTAqBKj4t+flPskyePQHXxdGxfvPvYmzR07iB//rJ0ielipARf7+o3L9rhhIpJsVs0Gtrwwjah3rGGs+Sf4L2ZCxiEkxPBk7uIAHVVT4uxc8zbQdEq8w/tTFh4aaucQj4sVhyIpp9ga/JyhE9prEDV6KVUyJJa6XCDowtnTnGLUEpvImYSEfC1gYYyj/EsaNbl9PAUnEcN0ssZ02M5fCN8pojTNf5G4P5SHKwjFl/s7YXUlpKdaHqHaIAbdiR8hHpJ59ZF2mCkRUzk4Vy5kMFqxSAhCj+C+BipvG/S+/+E/eAj/frqm2E1kBLgUkGYU8b1JR4lUu6RYeFVMYPv9RYIUrYX+LJLpktyY1OgfDm4AEt2PETUCH7O7JdlASJPx/7fmg95HDTpJOmvzIJwI8+kK0VZknpUEnsiaDFTLsqMNOuGW13a2BCpVwk+udYL7tcRDtceFJbpkMVkxquFtVBku76ItzmaZxkKfxsaL2EQVWHhUODzPtYUmG3gqokAQIdfBFl3pMgg9OJlxM8yNShGLi2Y8R0eszw85tR0fFf4Jm2pw8KGEjVYFEu200XzZ2NGiInNDqa+sw2NfnAVQoSYS4lBSRULH6qcQ1WQ5SAeBUSUZ1IWRBGJRDYwLmtqQ3MpEwODikEtLUdxQDVeX9wIU0k3T9/dQod8DmFyBJKknEy0NWngx2O9kWQFhIqGKYDHTjRs0VkaQiUEGTby78yahoamyU7dgmZeUlMmm6PSpSEBYbLYloatgz4cGJ3xOo4POhNAiTNeo69X2pROqtgApKBBDksY86xUx7cKAf7S2NCA0KQFdXByJjYjDY34vWxka0NzWi5NIl9HV1wt/XgsTwACTFxyIkMEDYFH7Uy/cywUKtUjOTXRZpc07C7MSsXuB1+xi66IqyyrY2tDRNysDa2+qDfvsoKm7cwPmiEoyMjaO3fxBhkdHInjsPqekZiIiMUvTLWwAVWj6D/UhV8Y7Cx2KT9mSy2tciLY4rlaWw+HjjVP4ZASoeeOhhJCYnYYxVOmazJFP5/pHWzePQo0IMVy1WSYwxP6Glnxhc0WPkjZdfxdM/+jGys7IEPNCMCkmwGQEYE7hN7c1ShawTgkzGszKVTIyxcWXOxv9YjTNAsGJkRIAzns/XakFqQhKKLxUib9YsRcs1AaOOEanOZdVpXHwimltbBKhg1Ud9dbV4VKxbv16YFkzY0ZB7sLcPM2bkIDAiwsWomJ8zC8EEKuDEGJNRFm+Yff1QUlqOC6fOYPPaNZJwaWhvQmx0HLx9/dDc0YKqklIsmpkrQAUZFSKO53DiyJEjyMrKcgEVanQex4WLF5CSmip+NMo01ilABaVmCFRoj4r8EyeQMW2aJLcoUXOttkZYIGQecJwpKysToIKm9UPDqnJH93f9L89JNg0/UtVsaPxLwHkLQJ7XMmFWdG2nvpUKGwEq5C5doMfkuYMAZldnO27cuAb7yACSk+IRGxcpLKvxcavyVyLyYFCjuT+r9BuaG9Dc0ixjY3REGNJSkxAWFiKGt0JJJyMK3vCz0iSeAT4DczUusUL62jXKLY2ip6cdUZGhCA4mY8ni8udhptbfFoCmxmYBC4MCQqWy9fSpYwgND4KfH+UorOgf7EdTay36+/tgHyFrg0w5O8YcNEGmpJ8dTnmvCP5YYYJFNPVpihyXEI/MzEyEh0bCPyAQjU1NCA0Lx8yZeSI5ROmk0qIiVFQWICTEhtkz81BddQXHj+3Bd7/3HfgFJSE4PB79I05cq6lDU309Th49hJLC8wgIppGxCaEhgYiJjEZAQJDIxIVFxsDbNwBOmTu9EBWRBLPTCxWlF9HdeQ0zZ0+HLTQO/aNBcIzbMNDZq4CKwCAM2cdQWpAPe99V3LZyIUYQgtY+mk1bAbMDQQE28ajgYohzEiujmYyjFN/oOM2z+yVJL/r+NKEeHBRWmsXK/uiEyekUoEJ8KqwWAXQDCVSYHOjr7kBTQ70YZvf0DyAtIxNp6TkIDYmWOZTMDAIV7PP0a9FAm/ao4HjkZm2pxOFkoILPX89R3N4W4K/8CJxOkW1kXx7qGxIaO8FYgpkaqCAQwiS6sMTIdPAnoyJE9iFQy7GMgAPvn++pFBSIjKIXfDjZG0AF+yrlf8hp4zzFuZPjpAYqeD8sBNBABX1BtF6zHkMFdDeZ5bj8jgCI9iJyST9Rt5lFCgTJrIpR0d+n/HsoJ8Mku46FCDaxrZQvhLcAVgQqNLNBbyeSkIZ0nEha0aPIAIc45tQ1NsnxwwKCBKRxCRCbTejunwhU1N64IUUPTICM2AcxPMrkvb+0K8dzHk9iFJPZBVRwbg70D1TMDx+Lqhw0gAAVqo+rd9yqqvPYL7WeMiUfCajp6kazwbph4oAm95znAgIUS5Pm75JouAVQIXrWMLmAChZvEKggC4JABdtOj7m8P0+gwuxtdQEVBCjou0PPGs5tXRM8KhRYQZBTgAr6WDHe6yTT549kVHh4204Yzz1CcoIFNMs+daIQF86UCEhBv4qOtm68+/pe2e0P8agIDSUzY53IWrz35l6sWD1PjnU6v1AYEhu3LcfwkB1vvLjTdSkr185H3twsXDxbiu7OXgElKstrcHD3Sdlm2aq5mLd4JkouV4kMlP7MXzwLS1fORnlpNQ7szp8w7QjAsEQBDIf2nnKxHh587HYEBQXg8N5TWLl2gcTkuz/6HM2NbWp/E/DIE9vFIH3/p8clkUNGBZ/t1aobqCi5itrrSlZJzYHuPs5Yd+mq+Zi/JE/AhYMGOMC+8OBj20UCcP8ulez/fUDF5DmUv9/76O2IjYsSoILrCIISBAg+8AAZ9CPl8nLrPeuRNi0ZR/flo+RSxU2H1NJPXwRUCKNi+xpJKlVX1KC8uAq1NZQ/vNmwWRVfjAtjb83mldKmO97aheycDJF+qiy5ggOGhFNyagI23r1B5GBe+c1brmt7/HuPyHiw76MDSEhJ+L1ARer0FGy6a70kz65WVKO8sAJ1NXWuQsPJN01gYwGBjUtlOLDzkGtJ+tC3HhRpq3079sM/2IZ129YJULHvo/2u5aqMgUbSQKSf5szAuWNncfJQvpJ+SozF4Z1uRsUEoOLgCWx5UDEqWptahHVxpbQSfT19bu+StBRsfmAbOlvbBajgmP3I9x8X4JiAA2WI9OfRHz4BW6A/9r6zS6RtPD+bHtiGzNkzpKL8/NHTrj+tvWsjZi6cjfOfn0ZAcCBmzJuFM4fyceqgArHYGE/8+En5yROoaCRQ8bvXsfWhO5E5Owcn9x/FuSMnld8hZeHu3YLcRXNw/vNTOL5X9W/92fzAHciZn4vTB08g/wATvmqnbxpm2i/84t+RM382Nt63zQVUbHnoLgEBTh08Joluna/41l//mUwnLwhQsRZLN6xG8blL2P3Wh/IcKe+z7bEHRGaJCfXbH70XuYvm4tQBAhUHsf1rDwkDhNJTxWcuovJyiRiFi38FgFXbN0rVf1d7J4rPFEgynMfih7HOrMVzsfURBVS8+czzwligRFLpucv47M0PBPBIzkzHvd/8qqyXfvff/8nlx/fk3/2VgBEfv/gWcpcuEHDm6M59yN972PDoYCL/XsxZsQgn9xxB6bkCPPiDbyAwJFjYH5SSqiwodnkR6ribY47Z24wV2zZg5e3rUXDiLHa9+r4hT+SDrz39PZGEIoPiWnkVfvgPBCrIqNDSTwQqHkLe4nkCVMQlJwqrhIyNfe99YlTfqzyBmBmbTPjWf/tzJKan4KOX3kbhqfMCVJBl8+5vXgZlwLgNQaW5Kxbj8537sO+9nTKPbnpwO9Zs34yCE2fw7m9fw9O//J8CxJNFQ7aHJ1Dx0YvvoKbyKr7x06cQEh6GikslIjNVdPaiaz5XBZ9GsdU4kDErCw8/9XUM9vXjH//8/5Fr5trr9kfvxqrb1+HIzv3Y9/5O/PSZv5M4jn2kgpJuJhMe/t7jCqh4/k15JwhUkFFBhsWpQ8cV+3kcUpQj3mOGr6ZkwCgzSi9JnUQ3QA2JOwwjeO7D+2MuiQfiWlv8HgD88lcqH8TPd7/N9YVK6GuwQO7D8IRgjMi8AkEIMaCm58OIkvsUOW6JN5RKCEEFiWWMwgdRutDm35SXpueIyFhZjLMrrw8plPBSeTdd+EgGhfa/4jlY9MH4iDEu74m5KcbMbAcyTfgd9+Gx1XkVWKNzTqrQVb1XCnxgoZLyeFEflZDTzrLSZkahKWOLL4GKCcPsl7/8V2iBn9/h1gSVV0An5W9hyqTeEU0j10AF53BOZho9mJSE/4OYCJNacrJRmcEmUFn8Wxzwlnn/L2Z5uGWZPHWQFHrp+rgYHpO2+X0P3gja5Eg3ISiemueeB1KUNFcT632Naj2X8JMLFRlXh3aZaSvQaILKlshFudtBm2p7RJfq+lw7TWxbdXx1Tfo29FeshJaBmv85DEbF2C2ACko/DQ1igMlcw6OCjAqVpFQ6gBol50SnTcNNyQYAACAASURBVKBopsxbZcKUyXcyF2xkI1ituFZdbQAVrOq0K2mNUTusNl+36ROvSaoFHWi4UYuh3n5ExyhGhcnLW6pEUzKmSYLE18aEIBRqzlp6mSDU5MFKD14XP5w0NEuDwIQYdQ5T59/PZY5K4IL3QIo8KwC1USU1vX2Z3DXajHrwBDoYtHFSiwyPQF9/r0gotTTfgNnHGzbR+Q6T6xgbHBUmCaUOaIhcWlos1QCeQAUZFUyoBAeHGklvylEpRoVqW6fIR1CeRHtkqAf8RUAFE4Z9wrRgoo/JkNamegT52zA42IeI6Gh0treiqrQUV8pK0dPeJqyJ5LhYzEiMQFhwEPwsPiLRYWUlLitj6clALUiLryQWVFJY63pbYLZYJIkkgaaYiilNS1ZfWC1eUmXqpHwRTKiub8S+g0fQ2NqO6IQUZM2dj7Rp0xERxSS1FK66qhTYT7T0E4MCSjGxWkJpTwZJgpVMCqsPwapRXKksh9XHC6dOnoG3lwUPPvQI4pMoFybZKJXIczhcQEVrS4skiagT3ter9PW9LF7S/xlc9XR14U0yKv7yJ8jOzpI+y/OLt4LW+TQopE2trYqJYfGRpBiBClYjT58+jZbLIn3BZBipy71dPWKGxvfFi8Cb1YLcnJk4fvhz+Tc2JkaCmp5+mqRTt5+SQYGiG2+12jBuGkdLXR1C/Pywbv06SW4x2COw4rSPIiNjGmyhoSihR0VlJRbm5ilGxbhDPCpsBJJ8rSguLcP5/NPYsn6tSCjUtzYiMT5JnieBCnpULMqdjaSEeIwacn2U9zl69CimTZsmfhRKQoTSYGM4c+6sMEjIqNDSS+3tnZIIneZiVJhxIj8f6YZHRVtHu7A3srKzJWnL511UVIT4+AQcPHgI588XY9wwlGTfUkaA6t22+HhJcnXVqlUuNoYGKlTQ76YhKwBi4kdvqxN4ql+r9+tW23NvFsgMDg2IvjzVSVlZHxQUKOwhM9kuHpJTikZtaKOSfTU0hO6eDnS0NonHhdViRmJiHOLi4yQIJnuBQIUJXlJtTSmnrp5O9A32YmyUrKsA+Pp6wTTuwMBADzo7O0SGinJZIyP0r2ESlKwAmuR5YbhvGL0D9KsZgdPJZLw3hkcGMTjSDbt9SN4RE2jcPCiyT/HxsfD188FAfy+8TD6IjklCdXWdJJ55jTNyaIadhrCQKJFqa2ppxo0bdVi2YpWAGeNOLwz2DaKk5AyKi88hKT4a3R0tKCk5jSef/CZGHMFISMvB0JgF12tbpVKuq60F+3fvRFdXHbKzMlBceAEBVm8xmQ8Li0RYRBT8QgJhC+TYGoWY6GkYGTKhrPgSenrqRH/eFhKNgbEgjI35YrC3H8GB/rAGBGJoZBTFBSfgGLiONasXY8gRiMZuSuHYBKgIsClGBSnbnCcI3HDRMToyJkAF2zU8IlwWSVzY8N2vqbkGq5WzqhPeJpOcK8CfiWYf+Z0YbmtrA65fq0Jbq6oMjo5NQALbLTwRIcFRCrgygAqykugPpBfrHI+4IBPPHAGIdR9SRvPsQy5GhQFUcDuRbwoMkPnKMe5UjAoWDvTSdJHSVAqo4IeVvzTMVsDGuOzLMYagBPsr56Tu3l557iGhoWr8N4AKMZ02e0sIKX4UYw50tHdIv9dawTQQ19JPwg70ACrYVixe0POzvkfOHTRU5gKZcx2vifGAABM+PlIIwGdAGSiOsXx3+Xw4njMRy4WuXnwKo6KvX5JjGqggyK0KFBQbg/cp54aqlOPP/JsLqDCZUNvYJAvnyJAwjHPBLSarjK1M6OrrkQWpZlQQqGB8QUBveGRAgAr2Lfm78RyVhJ2XS/pJgApbgDLTZscx4mJJABjyjpwbKOfIBTeT4jo+ETBTpJ9U5p5lFLpfNDbVy/0FBLAveUtMpBf8elzTi2yO5zTFJaOCwyVjIDJUyOKghOOIkdC5FaOCHhWU9uN8TLCOCQxKoHHx3d1FM216SymQgskCAhWe0k+jHWQQ3Rqo8FzbyM8uT7cvDuZj4yOx9U7KGwG7Pz4m/hCs1KdkE9vj0L4zqCq//sVAhT7F+Di23LlK5J8O7j0lfhQExSj7FBBkw/rNS0WObvKHbVx8uQqNda03ARXrty7DjFnpOH+q2O2JAch3ZD/Qd+LgJKBi9YbFmD0/2wXGe56P8ezlC2WYkTtN+uprz6mKX/2595HNUt2/f9cxASWyZ2Vg/pJc8eAQ0HJwWCSbTh8vcEmP6Hlx9YYlmD0/Z8rzEmQY7B+82UzbJaGrroJszWW3LRKggfIdes3K6z28VzE71m5egabGVux40+0vIX8wCt2EgREfhSN7TrhYGZ73OdGjws2oeMyDUcHts3OnC4siPFLJ2Q0NDOHyhRKcPqoq/GfNnYE5i9g+oeq+jQXUjZo6fPjmLmTlZAh7gkCF9pqgzJMnUKGXw49//xHFOhCgIh4Llyu2xMFPDI8KSj8ZjIodryqPCko3LVg+X7wyRMee13euCKePnNYkfddycPXmVZizeLaMO5M/HAMPE0gxQwEVRZpRoUvYPIAKSj/NyTGACnpUPOAGKjSjYr2WfroguvccW9dsX4/07GlSOMY1Jf0fju3+HE219eLloICKDux4/h35fdOD22AfHsYr//L8hMu971sPIywqHHtuAVTc/+1HEJsYJ34UpRfdTKNlG1dh/oqFuHD8rAAVWXkzcPCjvSi9YLBOTLgJqFinGRW/fR0PPPlVxCbFCyOj9HyhMroGsHLzGsxfvRgXjp3BiT2fu/MrGMfmB+9A1uwcHNyxB8XnL7sW29/46fdl3xd//isBJTbed7tIJb3z61ew/bH7RErowAefouSsqtDnA1RAxTie/7tfivTT0o2rUHyWQMVHsk1KZjruePx+dDS14q1nXsTtX7kXsxbNwekDx3Bs1wHpV5se2I6M3GzFjOS6uaZWJIQaa+rkGGvv3oLcxXPhHxQov9N34cgn+1BVWCbeCZsfvFP2eePfnhOPis0P3YWS85ex7+2PJB5KyczAnV9/CMODw/j1X/9C+QMA+B6BCpuvsA7IGElITcaetz8SOSXdjmvv3IwlG1bj9P6jOLZzH1KyMrDmnq2ISUqQJDC9+krOFuDAu59ghLK2hjcT58fb7t6CpRtX49T+ozj04WfStpz3vvGzH7jMtCmP9YNf/EzunYwKynfxc9c3HsbsJfOx67X3pQ3nLF+E458dlPbXsbguWuL7/fWfPiXSTx+//I4AI9/86x+KLNd7v3lFmDMcI+751qOYu3wRju7ajwMfqOtZf+/tIstEFga9SP7qGXpUKKCCkmQ89v3f+aowKghUnPv8pHiVbHn4LsTTa8XHG8ODQyLt9cmr7wv7Vn3Uu5yZNwMPff8JAaKe+9tfuiSotzy0Hau3rRegYv/7n8p5Kfn55jMvCUDC3MwjT30d81YsxI4X3sHpQyfw/b/9EVIz0/DWb17F2SP5RsGELqgle0CBCdqEXMka0ejaMIw3igOY1JdiCgIDBrtCno2wwdX787sX3JJH3/32RLlJ/l3PLfIMGC+z4NWuvTfVvat1mGIeMMbURWjq+li85a3YENTyNgCcySCCloLi/KziXiWppU3FFbuYJRqqgEQ8UqVYjWtZAhX051AFbK61oNQae64pVXpV1GrEt9DwHGThIAsRvRRbxagTV4/Xw1NXF498CVTcNH19+cV/9hb4+22ZcguTK+kn/+55n64UjSIhTErGTwpyZLE0KQGuQRDPg3psMy7CN3JVxsuoN9SIhDqx+qvB8PDcRCpaPM85OfAyolUXEOGRzPeolPU8AiWC/pCPZ7tpoEK+MwJUd37LuHrXYTUDw7O5JiIwE8EKvb1mYkzVVrolPdppwvPwhDImPSePNvWEoaT1SJvj1DMJqBixOzA8aphpDxnST0ODYiCtPSvmrNogzcGBlYkSItesoCXFn9W3vDNlcuSUZA7BDC74ueDlKH3t6jVERUdJhTmBClL5qKEdEBSkmBeSyBiTCk62d03VFdHaj6b0U1wcTN7eIkGQO3sORsZG4R8cICg3k+cykUivUv/ngEMWyroCQLHQKQllFmYAqaVcUPf29WN4mIyPManwkwU05UzGRgXMIL3P16KACspOcX96NSjpjTGRR+J9Uuqks6NJ9OdJY4yMiFLJ+rFxUIc8ODhAvBCuVlTK9U6bnilJ56TUZARHRUjSioAMJ2SaT3PhTkmgkREFAlEaRMusaDNtXTHOBQq9O/r6KP2kkj/eVgsG+vokcR0WGoLhwX7U1d0QhgQbNyAwSJJt508dR1t9HSxwIjkmEllpKUgMZ/WnWWQoKGfCJAkTR1ZvH9iole2jgApqU7MOU6r7NUDENZ1hiso2ZVDDgMKb76G3CWOsUDD7gDFOSUUV3v/sU9i9fJAzeyGWLFuFiKhYOAjwgPJk/F/FYxGJMF/qlPuKKTOTdQwCfCw0o6PEiAk+VNtx2HG1slyS12dPnYOPjy/ue+BhJCQlw8nAxwsqoHcqoIJGuU2NTaKrTR36AcOjwtvqjf4+BVR0dXbhtRdexN/87KdSST40Zpd3gokPJutURa6qzmjv6hQvBgY9TIoRqCArIDMrC/BW622LF9ku/eju6JTzsQKbMjJMkOXl5uH40aPIm5krLAx+2jpaMDDYp8xjDX1MCRbpFzMyhKjwEMzKnSUJM7KIuro6paqV/ie+gcEoqyhHVWUlFsyejQDqgrNCBOOSoIavD4pLS3D62AncuWmzLIzrWhuRnJQqPgJ1DbWoKi3BnFmzkEz5rHFadqvA7UT+CaSlZiAuNk4AGwEqHKM4d/6cmIfHJyS6cOXu7l65runTMqTtGdHl559Eelq6vG+syu/o7kB21nTExcWLTEthcSliE5Lw+utv49133hO2AYFWLV8o/ihmszBp0lJT8LOf/VSkwzRrUCW13MbaKjE5YfKa4CE0TskjCUJVr/McO2XGcu2rdOOlap2BrVFRxP6gqqVZzeOChtWOBlChZjAVGI+If8D/y957QMd1ndfCeyqAQRn0RoAECPYGdrGoUhStQnVZki05kYsc27GVOO/FJXlx8vvZ/p3nJE7cJKtakiVLsmRbsmRJVKFYxN57AwEQhUTvZTCYmbf2PvcMBoVy7CRrvSQeL5rilHvPPffcc77z7W/vHUNrayNqa6vgT4qJmUFwhmAgx3lHa5sanJzih5fghMuNzMwg6uvrceTwYXmWkBVBEIzzAplqTABLji9KqnIMwwNMsA8jmJ2OlKQMeNzJKCzOwlCkD7m5k9DY0Ij6hmo0N9Vjwbz5WLZ0qUy+T5w8htT0TCxadDlef/MdZGZnoLunA9OnTkNPj5HbmT5jGgqLCnD48FFcecU1SEnJkKRS1OVXgvPQwYM4fGgPYuF21NbswZ8/8CnU13dj5pzF8CXnoraOhs39iCKMY8f2YN+ubQJJerpb4Yv0wRcjo8SD5PRc5E3KQXpmkjxt0lPzkZ5agHO159DV04J5ixYiJS0fg2Fu1pMk30FWQ2owFQMD/Ti4ezNcQw1Yc9VK9IbS0NDGeS0LYUrzZAXkc+R1J4nFMjhAttaQ2CyR2JCksWj8zXiIax+9m6qqqpCSwnkxCncsgmBGErLS+GwNoaOdoHWT/pDyXVg8CfkFxZJ8Sgqkw+NOQTA9R6y+xsYGnD17VlJpNJLnEs81NG6m3dsblzUz49cjNlffYL+ACFcUmqPpr0MWnTwn+IyzrQ5QwfHT2zMAmn8TqOA6K5ZF/0AcqGA7xahwgAr+hv/uIlARjui5YrJd4LiM6smkYyWcSybVZO4xWc1ECdklNFbnmOQmku0Ro2KIfUo2Zj+SZQ5uKlGtbJs105aEm8PUsIwKSUgm8f4M69ESUEHjaY9bYAYf1lQCFY5cEttHVgznV4I+XJNCw1E0tzSbtidIP8mzgvY6ZLYlMCqMlJxHiWbGCPR8QWzYCcy4sQc6e7sQiUXku0XGRM3ZavUJPWgGBnpVrMH/ZlGE2JuO/xbn3mjELc+Mnt4uAZwEN0zRhXpFAA1l+ng8gjTJfmfzHzWm2OxLMioiw5yPTLPIKbQSZReajPQT+4WJAM2Hzoabs6itiOQJhXNEoeeJcxsZFWKBJLnR2z+oMSBjS4EN3LybghfFBj6fjNQJfKUHUpVYkNRXKISuznZHBpFFCzTG5Nj2I4MMxpQUtdkwKng/x5tpK6JLCG9tzDOenj06yr/0qiUCFHjOsS/2Cb0k3nljhwEq1l8qf4QXnx2RxBn7G5pP04ei6vQ5TCmfpMp6mmsbRsZlmm8O7qUm+ehXe1sXsnOCEzIqFl8yVz4Sm98eMZ1ecdlCLF9dieNHzowDKsioWHLJPBw/UoXGegN+6uUwpOnXcNOH1+o+/+q5Deho74p/5WOfvk0AkQUqbP9xzZo9fzoWL5+HtIxUbHtvD/Y4htL2x2JUrFggTwjKXSW+mJhuqCOjLhPX3nwV2ts68eJPTRLPDMqRBff629Zi2sxynDlxFvt3HcGFxmZcs/4KzJxTgXff2Cq2sGVUvOAwKsw+dSSxI0bFjDJsfGMrju4/Pq6/5yyYOeJR8dR4oOKJH/7MSJQ6vyT4x98svqRSQMr7G3ehvaVDUlKM//ft2I8jB09gUmkRrr1lLdpa2vHSU7/CnMrZuPoGh1ExxmuCzJCf/OCn8bbd9/l7DaPiJQeocGSdNjhABQGOa+8w0k8vPjEaYGIievaCWVi8ahHSM9Lw/tvbsef9vXHrLV7HqjUrsXT1Ehw/eBz1NQ3j709tA0qnlmDtTYlAhflavH8RgzwqLFDx1hZ8+FN3yUz7HXlUHNX9FKPisqXYu8UAFXb88SbllxZiyeplmDF/FlouNOPZ7//EABOWUfGww6h44D7Ng7947Hl0tLTH2/vH/+N+Jb5/8+zLOHemNh7n8Zm/9s71mLFgtnwAJBclpqoLa2+7DnOXLcCud7cJqKBvxftvbsLOjYa5xEjuU18yjIpH/8+PMG9pZVz6iRXwN3z0FsysnCtT4r1bdsbn0WvvvBHzly/Eznfex+bX342D2lz7CFSQubH1jfew452tcZnQ+7/6gM7zyLe+J3mmdQQqaurwzPcel3cGDa03v/Y2dr69xSTL3a7RQMV6I/10ZNcBvPI0JaWAshkVuPm+uyTl+uy/PCqpIbIetr+5CRtfceYrJzlMH4nlV1+K2Uvmo6nhAh7/9vdNHzifU55q6RUrUblqmbwRXnr4aeQW5YtBQaDiyX98UCbR9Kg4tvsgfv3UC4opZ8ybjZsFVAzgR3/z92YPEg7jgW8RIDBAxYIVS8VseecXv8H7b2yMgxk3//FdWLh6Gba89jbefek1/ZZrCNcuyj6t+NCVkqba9fZm/OanL8X7mfdtzW03SA5r39ad+PWTP48D8Pd96XMCKugD0VBViz/9xpe1p3vhwScdoILsh3t0fAIVNAVfcc3l2Pr6u9jgSCuZ6ckkn7nOE/woqSiT4TVZDp/4yueRX1wowOHssVNq123334Mll62IAxWMX6654wZcfev12EtGxQ8JVPxvUIaKbaNPCo9/12cJVCzDS488K0DDnpvHJIBB2SeawLN9NNS2n/P4HM8EKljURkaF8dh0Y+0d12PNzR/CO796Q0DFV79nvDEo/XTy0HH178ce+BSWXbECL/z4GbGQPvd3fyGg4vmHfyr2kNgkjm8W5zpbDMPzM28S96lwUGILPgkwcIqQjYS46UcrgclcxsOPjUg/febTTvLf61FOhuCMYWzEdC281/Qq5TEYW/C55n6fLzJwLROBz4tM2iVBa9Q8uAdUQWiE78VU6EFfSualGMPz3nJdYQGqUa0wbF2111Ft4DG4VDEm5MtIkkfEYDU+s5S4TFHbLTPEAhVmDBkGYpT7Rso/ObklU2hiVhobn/G6LdBnpLFhilP/YKY9bi3/wxv/BXrgm+tnmqT/GDDhXwVUxK/fQgZ8Y3xAbyq7bCLdsVdzDHjiQY49liO/NL5edeTYRqbJJthNAt6khJxzKLeTmHQfDzLE00djwAoli5zX2F+JOPKBr5FfKBmgmcU1qnrLTDT8P3OwkW4Rx2AUqDOWRZEIKZj8FVkViT3lTGa2/XEaxAQgS/x+J9678d9z1pFRybZ/M1Bx5bp4IEEgwjIqmHiIirZnNP2srjQTG0bCwmgT1tTUqPI5N49mrkY/kEE9qzW5eDC5ZmWl2BVnTp5CT3uHEvjFkybB5fVp875o6TIlIdJzMnXcOGXUqZA0FD5S9biZN5qLNiki0yJ5aPQpccL3uUmWD4UMo02SkUk4VicnAhWM95jiZTKElc5ccPJzcgUmVFWdRm93K7Kys7RpzcjIVGKHEjBMRqXSpLiuHjVVNUjxJ2PGjJlISU3HlPIpCGQFlYQtLCrWosqxxoS8qUINqXqAyW4LVFgzbVZLs60MHNgv1BRntT/vs9fPCulehIcGZYJKoOJc7Vkk+X2qeiSwsXfXLpw8fACxwX5MygliwcxpmFyUjwy/eSYp48CEkJKvTEqQTSEPCmM+7k1iQswrwyhWXjDRpKfaGdoMHpR8YoJCtAEXIky2uLyqGh8Ih/Ha5o3YtGcfgtlFWHfdesyZvxAxjxdhBi8UM3LHHN3tqPqETJPW1jZ0dXULIEpKDig57vfSR4Na+kM4c+qEzFF3bNsJnzeAuz96L0rKyg2MKqAiSYENq3l4jPMNjRqn6WlpMolnxoYyVX29/ZLhaWtpxZOPPYq//eu/wszZBCrCksOgFjcTW0xQsQqYz3Z7VydaqNXudstLY8uWLarypyl0zGs0wvk7mml3trYpKSowxxODL9mPxQsXSVJp0YJKzJ07TwmftvYWmZJSb9hQVIcRi0R03uQkH3LoeVBU4BjuxqSHz/OXlE6GPzUdx48dx5nTp7Bs0SJJctB4RVM7K+mTfTh09DB2bN6C265fj6zsIBpam1E6pVxGz/RDOHXsKBZVzseUyWRIUDrESKvt2r0bhQXFMrpXUs/lwdDwEPbu24vy8jK9T1YA29LR0SXJsYpp5UpyMejcumUbysrKlSSuqzuHvsE+TCsvE/ARjsRw5PgpsW2eevpnePzRx5T4stUnhu4ryz0kJ7kxc3oFvvnNbyrRauZna7zNQNgkVi2zIXEpkERTnJ1ElGJkHTHAp/lY/TVCnhNgY4FsHTsBnI8SkbJAhY43krAx1c7Gv4LMrGRWloLJ2y6cOnME1TWn5GeTm208AQJJyToPvWH6KevV0YXp02fhwIEDeG/jFqNRHw0bYJZgcSyq552AEBPJBDty0rPR29eBhYsXICU5Awf3H8G0GaVISolhx44jOHToINyuEHJyg1i9cgVmTZ+L9tZubNuxCRXTZuGSFevwq1//BvnF2aitqcK0qdNRc7YG1edqkJERQH5BjuSmli9fjeLCMnj9KRiK0k+IFGngyOED2L39bdTW7safff7j2L/3CCqmz0JZeSUaz4fQ2hFCGEOorjuG4pxcvPSLlxCN9aO8KANTCrPhdiVhx74TaO1uQnZuCsomlyAvpxDJflP57/VFUTxlBjxJeQgP+TE8nISenpCqntOz0jDQ14P9u9+FJ3oBa65ciZ7BNDR1cH7NxmC4H2lZKUhJHgEqBgiyD/bJq4MslCNHDmPKlDJkZprqWgIVNdVnkcyK/tgwkv0upCTRk6gfzefr0NxEOQufGBTlU1lpmo6hCDckyfD6k+GKeZGeliGdWzIqCFTQn4KMCoH9LvoiGd8msho0bXGDRQ8NeNDd24vewX5VfNGTICUpGRkCKgzbguuGqOcqKDCm4D09/fAnU14uWYUA/IxAhTwqUgNaK2XEnZIimUG+BFR09WiMESinvJTYidQlFnsRkgQcoHRYhD40XYgMDyErIx1hgv9kkBHwdsys7XrLdYl9dzGgwsUNqANUkOHGtV5rtANU8Jk3cmd+zSOJQAUBB1utx/NxneecQO+kwXAUTc1NzvNE1pMpupBZuWOmbYEKK7fFooILdW1iT+XmBOHy2GeZyZaYgAr6fAWDQfVNbU2NxmR6RgYG+3oxMNgvoCIlJVlgI+cCJezdfrhiPjQ1NaOruwNpqZSHYgySZMDYiAvhCJ/rGNxel4oEksiKcGIZtpuVe9zIy6PC1r3AVAtyvCQCFYbxNjpxHJ8jCWqpIhKoI1ARNUBFSloA3iQP+vpDkpuyQAWPZedhA1R40SmPikEBEEQ9CPyz/zvaWh1JPohNaEA4A1SwEENJhg+QfkqMte28/tuieX5+573XoaAoB/t2HRMIYV/0glq2Yp6kPZ978jcyohZQ0d6NF59546KHpkH2zXeuNcUJXo9YEDSw5r/v/Nh1uneUdao+axLFZCrk5GWKtTFnHlkSo6WfRnlU/GzDiEfFXdc4HhX7xnlUzJpr2BbNTW145edvx39TNrVE46CuthG33LXOeFRs3DPiUaHzrzIeFY/9UrJP5dNKsX3LPhzae0ztJRixbBXlnU5jw6ubRvUDjbPXXHspmi+04uUX3hw5b0WpznuupkE+EdfdvEa+DC88bdgQo3c1wH2fvUsV+G+8/C7OVZt+uvGOdSirKBWjQh4Vn7hNTCnrUcEhe9W1lwrM2LV1n6Rmlq6iR8WJuEdFUUkB1t1Ej4p+7N1+EOtuuhKdbV147nHjZUDWxM0fuV5tpUfFupuvEqtj23u7cXDPEa3dq65ajuWrF8m3gvG79bB485V3xZik/wSBiebzLXjxqZcxt3IWrl5/JU4eOYW4KXZ5Ka69fZ32ND/5fgJQ8YURoIKFIJetW42qk9V47YXXFRpMn1uBtTetQcuFVgEV6269Rl4W29/dgYO7DXtg1ZoVWH7ZMhw7cBxv/vKtURpVZF9cvX4Nmhub8aufvixGDV9l08s0F9SfrcPsRbMFVJw6egpvvGjG+QhIYYKc0UDFVqz/yHpUzJ6GLW9swv7t+7QHuGr9WsxfXok9m3eJLXD1LevQ1d6Fnz/yIvfjMAAAIABJREFUrCkEc7lw3//4tJ7tN57/ta6PDAr6rr3w0DP6/NZP3InSqZMlqTTiUTEPa281HhVPffcxk5tkMp//c7uw/MqVWHnNZThz7BRefvJFtZ9z6t2f+6O4l0QwOxNkWPA79JvQvS/Ixe2f/IgK4ARULKnENbcbjwoCFSvWXobV664wfhM/+blh6Ccl4Z4HPo5gdhBvvPAqTuw/OiqBTo+Ky69fg9NHTuClx+iB4FLi/MP33yMg/eFv/otYD1b66ZnvP45Vay/HpdevUfL6l4/RqyMmaSFW2zOe//HXv4vL16+V7wCln16h94WL0k8VuOW+u0dLP61YjG1vvCd5rOs+egu62jrw9D/+OP7Mfubr/1P9/+YLL+Oy665WMvpXj/0MrReaNW/f+8VPY1JZqVgbjKEFVNTU4el/eijOqJAB9hPPKa9RMWuGkvQs7Hrob/9BCW7GKV/45ghQMalsMq68+UPyqKCXhqQh/X6ZUtNf4dWnfo7c4gIsX3Mp9ry3HW+/+Iru7cJLl8u3ov5sLX7y7e/Hk+WMbeZfsgQ3f/xuGVo/+Z0fqSCS1/XxL38e9L0g26HuTA0+9dd/hpyCPLz0yE9lAM7XvX9+P6bPn42Xf/K87p08Kk6ewZPfeVCfEwD8xJc/L6DluR88IQCodFoZfvHos2JU/MnffFGMCoIfJw8e1fV8+E8M4EDpp9ee/aWOex2ln265Ls6o+LNvfUWyVC89/IzMv3lv7/ufnxEY9tKjz8pInvJeW9/ciDeeo3xUFMuvXI3b778H585U4wdf+068cp/PLuOQv/zHv1MfvvDQ0zi4fa/6/9ZP3I0r168VUPHqM7/A//zO3wh0euGhn2L/+7sFJH3ub76IWQvn4NkfPokd77yPL/7/XxFQ8bMHn8TuTTtM/KNEvBk6g6Eh7fdNXDaSU2IcYk22DaOSey8jY6n4Ixpx5LxDAgoGh0J45DErvQR89jP0gnAK6+RV4dFzor2QAxoYD1Ejx2XjEsN8GTHqtrlCJvhN4YXj9+CAJNx/ihE9FI7vhdkeFnUwBzU0HJIENednkzcy+zTiDMwXmRjJgCT8nOAB13dJP/HflDyN+x6aPkssfGP7WNzE61AfiQVtDMAT+9PEfyaGYixu46k/MCpGhR1/+Md/hR741vpZJlk+Bqi46LVNkPNOfHguClTEQxozoY0CFuLRjgl0DJQxPgFv2yQ5DLVDDb/INxMbehFGxdiLTNDZ/L3u7aiSLXMlppLL8fIQauocmQBG/Brs1Y6e2EfAInstiVVhDuAz6uqdPonvNh0wZExv2nttkmIJ4E7CojL2+keKgAmOsHTOVMLJo4IV2Qlm2kzO00Rbck/8u3+09NPCK6+J6/ExqcHKTC4EBCpi4bAq4JkYYKKUG25K3piqRJNUpE4332f1KGVxuAhz0WVCjkkHUyFoNMGJbp88dgztzS1KeE4qKeFOV7rbZFQw0ZyWTb11k8RRMs/xCqAEARc5q5NtQHEjvcJz8PjWZJPJFyv5wIVDkg8enxY7sj5oysQEuUa4y9AbjXQUPS6Agrx8dHS04szp0wikEARhgqdX3hbZ2dkCtpiEJVDReK4ODTX1qp5MBCrcTCAFUpGZlS1GBRdKC1Qw+UiggkkyJlzYPxcDKijjwUp/XqfH78XAQJ/amZudpWRd/blz2nRlBjNwoeECdmzdjNbGOuSlp2DutHLMmzEVaclJ8IELa0ztlOGlUzHOKn2/yyWGCSWxfEkpoOwDQQqXm2CFTQibsSmzKlZhsqrR6PQATO55fIgNRQVInG5qxLOvvIya+mZUzJiD69bfgsKSyRhmX7PCnVUUTnKefcKkD2WEOMYIMqQE0lQ5QV17n5sbmwiqTtLEDNi+dTv8voBhVEwxQIXL50JyKrUvh6QlTHCs6fwFjUsCMwLdSPlk//UTNHILqHj6icfxN1/9CubOm4OBaETyTgQKmEBSUO6lDAnQ2dMtoIL3gIDdls1bZGosRoWPiXyCKj4M9Q/IS2Kwr08JSLiG40DFxo0bsahyIWbPni1gobunS/JiMq0VC8T4q/g8bmRlBpGZkS6Kan5evvqdAIkBKkrhTQng2PHjOHv6NJYsrESKn5W8lATiBtAHTyBZQMWebdtwx/qbVNXb1NmKKVOnIzocwfnz9Th26BBWXLIMpZOKjcmyMy/u378fuTn5yMvLd2RNqDM6iH3798kkm8wImuvymSPoRxP3qRVTTOWM243t23cJlKAPQX19HYYiQygpLkRhfgEiMRdOnK5G/qQpePqnz+PBH/5QQIU1w7bJSI60ZB8wd84sARWqsk7wsiAyNQJUmIr4xJeh8zo8B5EvxkPtFqCwYAV/T7mVeBvG+FxEwcocmzlMBCoSAFP1vwuuWBihoT40NNaiu7sNwcx0SV/RL4WScZxPS4tLUFQ8BU3NPTJ+nzFjloLmvXv361IKiwrFHDh2/DCOHzuKYEYAq1Zfgry8HFSdOY3c7Fzs3rVFsmXpqdnYv+8QorFBrFi9EFVnG/Dm66/D441h0cJ5mFpegcxgAS40tmL//i249IorMWfOSrz0q18jOc2H7q42VM5fiIz0IGpqq3Hy5HE0NV/QfS4sLMac2fNRXjYVRZNI7c9AeMijjcK+vVvxysvP4HN/eh86mprR3NqKmXOWoKePfhkuhAgwVh9D5ez5aGltwabNryMrEMbsqUXIyy+CKykLB4+fwK4929DacgFTJpVhZsUsZKQlweMNIZhTgEDGJCQn5yMcCaCzcxiB1CDSg0H0DXRh/+4N8KEZVxGoCKWiqSsZXl86wuFBZAQps8dqfD+iYcppdYuCH42F5Qly9OgRsVgIHPLe8J40NNQhLeCGm4DnYB9ami6grfWCQMCSkhLMnb8YWTkFAtwGBocRCkfh8SbB608SSEWDZbLyCFQQwCdQwd/Zsci5nusZwQILxtMTiMBpV08PegZ6JfVGoILAc0Y6WYlGrslI7ZhNG8/BiYkMGJqEWqDCMirGARWBgIAujt5eARXdqtrnWm59MLi54gZVcj4uSFqLQEVrW6eun95Gw0MhxRa8Bl6LihJCIY1X+WIkcQPoSAc4vg2WUXExoIJVybw/nLvILrMeFVwLuEaJOZCwBnGt5L2Sd43Hi/6hYfnDaO50quds334QUNFU3y7QPyc3Q1V20jmmHMFQBF2UVyQ4wz6LxdBQX2+kGoNB9Pf2aA1OBCo4Z/hE/SOwmySgoqOzTSA5N9HcGGutjLpUTED+2liggtdl1lcaSP52oIIeFaoRklTkSHFTIlAhqcVoDPV19bqH7Mtk9iclEPsHMfQBQAWLImimzXUpMz1D0SgBH65XlMQ0sldGUoLJBSv9xETWfwRQMXV6KdZdv0rsMrIeCEIkvghi5BdmY8vGvWhqbMUNt16h54U+Fi1NbairvTDhNoLyTzPnlKOzowe/ev6t+HFXXrZQ5tRkYB7ad1L3nx4WaekBmWmzzyXnlOBRwRPc/OGrUT6tBPW1F2TCTWmpqTMmi61BRoT1WEtszG0f+RAmlxc7v6kSIEK5J4IQv37xLRSXFuLqa1dpCFHKicdYsHi2gKet7+3Ggd1HsWjZPFx61TL09Q0IqGB7K5fMQWp6Kra8s1Nm2mNft330eoER9bXn5WnB5D9llnjeV55/A6lpqVj/Ye4P3Nizjd4draiX78XIenrLR65H2bRS1NU0oq66HuXTp4AgAxM5lHI6evgUVq9ZjiWXVArwYNsoRTl34Ux0d/XiNy/RWBq4/vZrtE4eP3xayX0aXecV5Aik2P3+Ptx53y3Izs3C8UOnxIDg57kFOWJKEKhYtGIBLltziVjMB/ccE8t8wdK5SOP1v71NTAoacrMy9+jB4wLWps+uUGxUXVWLXzz9ilgYFqiwEk6Tp5biQxMAFR//wr1G+umlDYrf13/4OskkHdh5SLHRvMVzEMwMyoz654+/hMUrFwnM6Ovtw6HdRsN/wbIFpn0btmL/jhG5IXuf7rjvdkyeOhn1NfU4fuA4cgpyMHfRXHR1dOGVZ15B0eRCrL35Gkl0EXSoO1snOabE1yig4u2tWH7FJVh19WodY/+2vSgsLcaMedOV4Nv13g7s3rQTt3/yThSWFOHM0VOoOn5aGvhkVNB74rmHntZvbrznVlU/79q4HS2NzRpnV996rebLA0y8hoZQuXKx+ncLDbbf3xNPoipW5Jzp98k4O7+4AKcPn8DZE2fkE1E6dQpOHDwqv4vsvBzc9Ee3Izs/FycPHpMBNVkReUUFaGtqwaN//0PDqLj9hjhQQVDiI3/6x/Hj0qx77tJKTJ42BccPHBV4YeI9Y7zLF5Pit33iLuTk5+D4/qMye668ZJGAh9YLLXiY0k9LFoh5QTDnmX953Pzmk3cJOKExOYGSypVLkD+pUADCQ1//Z3kOEGih9NPLT/1cycyyGeViVPA7P/3nR3Hjx26XjNP7b7yHbW9uwkf/7JOYVFYigIAgyNQ5M8T2aKiu0/Xe9ScfE8Oi9uRZASB5kwqxePUy+YiQATCpvBQ3fPRW1Fefw0/+4UdiDFAK6tDOfXjt6Rd1j8pnTcNtn7pHQPSDSqRHpS7wBTIZUlLw0qPPoL66Fp/40udRUFossIASTPTSoNTT0d0H8PyPnpBvx01/fJfm/N0bt6Kns1uJ/6KyUmx7/V0ZSZtqfZOf4IugBK/pzOHjuj76YEyZUSHpXHpUVB07iZvvuxvLrlqtRP/+rbswfcFszFo4T8/Wy088j2N7DuHeL96P8lkVOLb3sCSv5l2yENPmzhJ74vkHn8T9f/2ApJ/IwKDc16f+6gsCn57/0U9w9thpPYM0xV5yOT0q3sSGF17VdYjZcMu1+s3zP3pSTA6as9eeOiuGDqWb6CHCBDYZFdzD3HH/vYr9KWlFYG75VaslA7Xp1bfwylMEy4yJtpLjkSiu/+gtYg7xeX3/zc3Iys0CwTLOKW+99JqAirs+80cyeD97okrsiTmL5+v5ILv6+YeekfTTn3/ryxpPNNOmR4VlFbDKn7El12uyGs2+3RR0qg1ixpLNa+WhTP7J7qVYMMFYzDJUmMN49PERoOIz9xu5TgIEZDqIMSGJL5MvMICFyQ1yLeDaRRUGxjbKljlVt/IJtQwGjQ7DirD7SdOmmOKLoRDZIi4dQ2OK3hHRsJj8PIGeZ8lcmX62oIidD9ke9h0BER6TOSVrzB1f02KjVWFYLMrDU22CfSigyWP2guYc5uiWSUFAwxa8Mab+A1AxYdj1hzf/M/fA7wxU8GLHgRUfBAokgBL2a3EjGNNzo5gQmlJGJ4HGn5C1cPblcsgTicyAMY0c5xMxmokwiqnwb7mZifJVCVVnht7laPg54IW9JntuM/fEa29Nv4yRaLK9ZT6MIx5jWmzPk9Cv5mCjv5fAqPig61eLLDtETRxhxMSBCiG6wxgSCk2fCkrajEg9GTPtEY8KAhVMPPBIrF7iwsZ/M2E80NutzTyTEZyUuTllot4CBGxCQ0OjktnUr6fkga365PeYXFEFaH+/FgUmVI4ePoyW8+elgV9MGRlp4Ecxv3KhZC8ysjNHzCnJImDygZIWlKVyFgpLCWS7yHxgFaul/8ljwElqWn1CshaYdOZiS6CC7/M96RhKr9FUozPg4H2fVFykRFNN1RmUTMpX37CKmbIrZEGwWvz8+Ub4U/yor6mV1mRKUgqmT5+BQGo6SssnY9jjQl5+oZLlknwYIpPDyGUQqGCQEwwahgaDr4mBirAMiXv6eg2i7yXlsU8V+3m5OQIqzjfWoa+7G6kpKTh76jQO79kD73AIc8snY/6sChTmZilxSnYC+5HJICV0pAvB5EkMfkrtJKXIINRPsMKfIqCCiaC43rUDDNlnQXIRZH8w0UZ5HLcXGObYi2DA48I7O3dgw6bN6BsYxtyFy7D2uvVIz85ClFkwt6li4HXzPrBym6atllHhT0oR6OD1UFIJ8Lpjkn4iIPP+FgNUkFFRWl6hcU6gIjXNyJ9wg8SNI4EK3nNuSFk1xP6m9BO1wAlUtDa34pknn8Bff/nLmF85D6FYTMCB9Nj9RhaL1fG8932DA2huMSaWvE8EKlj5NXPmLLiSvKY62OcTSNLT2SUPFgaBUVBGzYPFixZj06ZNWLigEnNmz5ZMWN8AvUYGdS9Yudra0oKMtHQFUlnBdAQz0tQG6tzzeSNQweeydMoU+AOpOHr0qBLWSxculExMhJRYVXz44E1LwaEjh3Fg127cefMtkidp7enEpMnlamNrSxMOH9iHpUsWobiQ3hGUXnFpo7J7925MmTIVBfkFCvgEPDqMCj7jSrzGTKDHZ7K5uQnlU6foueEmbPv2nSgtKZWfy+kzp5CSmixQjYBLJOrCyapa5BeX4plnX8APvvd9A1QoeGcAS5sa9rsLSZ4YKufPFVAhkM4BLlnRwufJABWGIjwCVFg+nwMkyIR3gumWv5Zn0Gjpp+GIlZQyzI3Rc75dx0aDFJz7eX76SbCfGhsITnQgEPCioCBXzLLwMP0u3MgKZqD23Dns2r5DSfQF8xcjOSlDevwVFdMEfvH5EQOL7Ke0oJhbe/bsQG3tacRiYcyfPxOhUD8WzJmFTZvfUTLpQkM7WltZBd6PFasWoKW5DbW1tZg+rQIL5s/HQD9pz14xYOrOHcOatVcjO3sqXn71N+jsbcOk4nwxKpL8KRqTNNzlJmffvn04ceK05rD8vByUTZ6MsikzUVBYJsN7tuPV136J3Nw0pCe54E+m35AP/uRChKOpSnafPnsCi+YuQf9gH2rPHUX18e1YMr8MJaVTEHalor3Pi/6BkNgMB/cexFBvP6aUZmNqWQbcKW64/anIyqL+eT4GhpIQSMtBegbZJL3Yu+sdpHjaccUVK9E5GEBzjx9ubwpikRAy0tMktcXNWXR4WB4+XV1tOHX6GE6dPAG/z4s1a9YgNydbMnP0PWhqaoQn0ocLFxrQfOEChsNRebLwOSeYkZZZgJiLXiDD6BsY0vpKoMKY/NE3IFVJdEp4sf8to0JRlwyQ0/Q8kS1gK+S1DsErMLS7v1fPAs2TCVRQspBsJ8uKsEAFk8cMo7rpUeFIPxlpRSP9xL5JDoxmVAhgd7nQ292Nzq5ugYx8j4ADE0bSBXa8YdjW/sEhDA0DlLnhTEYfpBilEyXJ59W6xbVMoIlM5R1Gxb8CqEiUfpL3BQ3NMeJRwXYQqOCcwIQ8ZRlNAQ8wPDQsRgn7kv5WfaEhyTCaNd1srG3fxoEKny/uT6ECBo8XFqjIzslAIJUm4HxGogjx3obo3zCkYgs+2+cbjTlsWno6eru7MOgwKgiCJweMUTbHUzRKCclkARXt7S1qI+Wh2L/sU6/LZ4AKzkserrte+S4xfLR+W2wD78UHMSo496anBxwZFSOjmAiwahPPAg5HCqG+rgGuWFSJ7ThQMRCSb0tirGQ395TOYdzFeYnPRWY6JbDoS+UyQEVbC9JSOZbdYlTw3nA9pMwi7wFf/96MiquvXYH5C2fIH4LyTmNfRhZqDk6fqMVvXt6MNesuwbyFM/S1Xe8fwo6tTASPf1H+6bI1S1F9pl7+FImvJZfMlSwTYwu+err6xGigmfac+WQkjAcqCEpdfe1KVMycLICKVaUELTa9tRNtrR0TtkG/uW4VKmZO0W84FprPt2Hrxt1iVPBF/4kVly5GMCtd95rM0L07DmHvzhFt/yXL52PJygXGgJ4eNg5osX3T3ouf94bLUDGzLOG8rdj67q44O2LNdZdi/mJ6J7qwc8s+7NzMY40AFQQlrli3Sh4TbFdnexfaWzsxpaIUe7YdkOwSB+iV61ZhTuVMJZw4zprPt2LLOzviskalZZNw2TUrkV+Yq+PQv4FMiM1vGZNl+k+suGIpMrODesb5e0p/MGllpZ+WrVyEpasqR66/d0Dsim0bjQzXpVdfgspl8/Q7PmO1VedQUJyvPcFzj72IihlluFoeFacQl3CamsioeDrej/d94WNG+unFN3HubB2WrFqMZZctkUysPB3qL8g/pLW5TUAFX0tWL8ayS5coqa/709uPg7sOYdu7HM/jvbMYu669eS2mza7Qc8Vx0dTYhK0btgqU4Jxyy8duxdSZUxXzvv3yWzjuSGdZ5su626810k/v7cT772zVenHNzeswfe4MzYlMVLPAqbi0CHu27sH7G7YIALryxqu1j+FczzidIMWm37yLxlqyZmK4+pYPYcHyRbq3rOzevmGLkukr116KTO45OEa7ewV+0GuCL+1dHWkeCxBk52VjzS3rBE4wgUgQjqyGN194TXMNX5SauurGtSgoKdK/ud+iJA7XjUe+/UPMW1aJdRao+OGTmhdzC/Nw9a3XYXIFj+sVI+XU4eN4/flfKwa2LyUWnQR6+cwKeQQUlprz8JrNeSJ4hEDF0kpJXp2vrcez339CUjcVc2fg6tuuE1ih35xr1BzLtiUCFYd27lfCmsD9lBlTcfN9dwqoeOqfH8FNH7sDlSsWS3bqvZc3IK84Hx+680Z9T/0fHhY7gp4btWeqtabccM9tMgxnMlnPU8MFvPfKBoE5ZH6sv+c2AQ0/+c6DWLR6mcy16VFBGST2fcWcGY5HxQC+/1ffNknkaERABU2sX3rkGZw9cUqAEE3D6WlBiR72I827yWro7+tT+xauXIYrblqHnPw8x3ulH0d27cfrP/ulisRU2ObspTh15BYV4oZ7b8PU2TO0p6UROBPelPl64UHjSUGPEcpVTZ09Xd8hiNFUd14MiV89/pzAC46H9R+7HeWzphtfiIFBHN97SFJLlLSiJ4VlVPD7ZFQYM+2foPo44+kYbv3UR7D08pUCKt547hUl1wlU0Idj7+adYlHkFOXhlo/fpT5TWzq7caGuAZOnl8eln5Zcdgmu+fB65Bbkx/tg//u7xALq6+nTPbJro0203/nZP8LSyy8RODHQ1y9pNIIOG1/ZgNd+9isUlhTj9k99BNPnzYqfl2DYlOnlAioo0/YX3/6y/v3THzwuaTRTqGDkk7j2yMdriObV3McNax3nd0LhQRXucZ4w0kfcKBk2hfbMBAUkYcT1yLAEHkmQfvr0p4xcJgsu+RpdSGa8LgQMDJu9pZjDTnGwQBRKRTnLCN9nfoSBkPUptEAF4yDmAsjg7e8fFKuTx1TcSHAtSmlc+lqm6pmzjBVTrGYZ9wZQYF+wEMd4TJjn3sbUo/KaCXVtLg9lUEOaK/lHBSXO5/y9YaSygIhsEvpSki0SkT+l/O+8hcvHl8lNuBz/930zc8mH8PF1M5HVdhjPPrMRJ/r++/bFf4Yr/xaln8YkxaXK9EGeDB8EVIwDBRxmQaKshcObSOyfkWR5dIyckVo3pivHMiQSPp+IGTJBmxIrXv/dgQr53TjGQXZDJ6DC5GlHN9GyGvj3xECF+U1iH9jv8oMxzJMRBl4iBBQ/6agz2J346G+O6utEOERt+ECgYhj0qGASdRRQIRPtAcenYhCL13zIABWO0aZNmNMbgZvy1ECKFgJO7qwwZGJD8lA0l3W5cf78eQWU06ZNUzLVAClRZGVl6rsWqGBSkwv14QMH0dncgoKi0YyKufMXqNLeAhX2wlmhx8pK/p5tVDI6bFgeTJJwgVTlvNMuW1FoGBWUnmJFAaV8uFDTw8AYfstAVPIrBtHn/WZCm4nSgrxcnDx1Ep1trSgtLdJ3O9o7VWFIXfPc3HycPHkCgfQAmhsa0XKeptUeVdgH0tKRV1gAf2oKsnLzHMYEZatiAgOk6x2mHBZZJyOMCi6AWviYsnESsKxe5TXSAFoVGX4vBvt6EA4NSs5noLcX9XU18q1obb6AxpoatNTVoSwvB4tmTcek/GykJHvh87mU/GVfKeHA63fOoSAyFkVKcsAAFclkVFCixA8PQQjSGRO4kDaAUFIriVJRKWIV0CnbEzbPWb87hprmJrz8xgYcPVmFmCcFH7rxRlQuWwHmgn3JZLiYQIqVChaoYP9yrHl9ND4PS4LE73UhNjyEs6dPKCjZsXUnMoM5uO2Ou1FaViaeCDwxbRAJYDFRx4CFQAXHAGWWZF4eGdYmjZWkTF62UvrpkUfwv776FSxctACD0Yiqmjn/MPGvii+vGRu9/X1obWuLP/dkR7DKcM7ceXD7vcbbwsNAeUBAxVC/GUcRDCmRs7ByoaSfli1ZilkzZykQZOJ2QFrnAdRUVyMWjqiCWswlnxf5OdlKfBIYYPuZ3GRCtHTKZLh8Ppw6dUoJ1+WLF6u9UZqPSxrGBT8r8U+ewNF9B3DztdcJLGnv70bxpCno7e5BZ2c7jhzYhyWLaaZdAhc10z0ezQnbd2zH9GkzUVRU7JiwUWszgp27dkjGZtKkSfB6mNjj2BxUUnf6jIp4ELp50xYZftNEnn4pGZnpMiQuLiwmjoUjJ04jr7AEP33253js4Yc1dxhNVFMBY8aXC8EkLyoXzMPXv/71uEmaknG8RocWzM2V2WSaiZbv2w06pdzYbm6+pLvvMZ9YHx8yesiesYE6x6LLnaTva9OUlqZ2MLhVuyitpWfI+PUwMCUwQZ371rYWo1sf8CMp2Ss9f1ZYa25KDsCfHBCThVXYnLZZcXX61Cmx0bgJYMJ47ty5yMunZ41PgJ3XyyRojpF5aKjBqZNHMTDQg5aWRh27rCQfdQ012iz39oSRnzcJKSlenKk+goH+buTn5eKyyy5DdU0dImFWD7rR002T9z5cfuWVCIWSsHXbLrR1t2DmtDLJfWVlEgQIoqG+QX/TSPz9rZsdVl0vhoci8HtSUJhfgrLyacgvKEBKRipe/fUv0H6+GleuWY0hJl1jaYA7C30DEZysOiWggvJbjRdO4eDON1A5u0ReK6nZJWhqc6O3bxipaUGEQzHs2bYdp47sgN/XgbySdOQVFSI9IxdefxBJKVkIBvMRzMpDb+8Qdm7bjGBqCJddtgodA6k43+WB25sEV3QI6amUfgrQbQeRcBhtbU04duyPqW7/AAAgAElEQVQQjhzdj/S0VKxetVKAdDQSxmB/H7o7O1FdfQbd7U3yBQoGs1FRMROTSsuQGsiQB0kgPQtRFzcgEfT09mE4TE1qzq/0mTF+ChaoINBNYI+AvInpYloLOCeRfcCxwXFFoCIacaGnvxc9A30Ic5MT4xyUjCAr2V1RPftcN2winmshBxK9mPgMWDNtjk9u1vv6+5RgYYWZBTkME5DgBn1lCJSYcZfIVmJCnY8JV/C+QT6XlLrrlql8gAnGoRCGHZlEK60o/yX5ZvQJrOUzZ9cICzByk+pNZh+ZjSuZl9b4kLIPkdCQ5l2ZayeZ77HdXBPTUgOScOKLv+Uf9jFBBEo/dfX2C0S2QIUFLsWIc6SfJANFViUl/aQHTemnVgwNDSI1nYw+kzzltYTDUfQPDQioYOKdx7NABf0dero6EQ5TgixNbD0S56yxdCRC8N6PpguUfmoXQ5FAIuMQ6TZHxF3DMPvIFUMSTb4pjeAkyhgjWI1lFifGKwtd3OSbiKipuVF9l85kp8i0BBuMTJ1NFth5kkAFKyYp/cR7SjNtxizcRPeTeTg4nMCOHWFMalOe5ENvbx96unsEVFCiiwlYjj3GhUwciH3jcctLysosMp7i+SMd3t/Ro+LfeYeWqN/wbzn0Bx3nYsz3i/1mjBH1b23WGFmv3/r9BMmP3/rd3/IFExOPf9n1daLPLpqQGVuXlZCgmmhHOUp7I+FEFzu+3mfhjPzKvPpvUIaExQ+MCUYo6M7RjHmLIaOz0ptVsiaW0DOUeHF2kyZp39FX7dhUjesKsyO0rM6L9aIth0vcJI6+wgmIoGYtcQ5J+ZKxr3E70/imkexnFhKaGCu+h1VsM75ndW32Ap2D6rri2UXGUtyvaMeiZphK6XEJCX3G71pwQuuDw1hlzC4JWUeyL1GWWv/tnG+khRP0qx1PKkAZrf+gPfJFBo5Jzo6AJ1o7Io5fGq+JRdvaJ1FX30jFMBdjxHD5mQvpWUElxRn7cx2k58aN996B7s4uGXBb8Neu9/y95vWxY8neyImeYecCZDRMUN9jpHNoJGw87kwskXgutk3sRqfAzPj6uCQ1a75PiUcTo5Jtbtkl6l3Ha8P2h80/cT02EkEjHgI8Br9vJKMZZ3vEZjLHoZThCMNS65JA+RFpZ+1rdQzz3cTYwSab7ZizY/Zic5MZQ0YmyMYDJgnP2zySp+J18Lq5bkpSyOvX3pHvKXE9bOSZOC9wfNt9ieYJ5g0cUHHUc2THr5M3EjimvmaSnnOLKaLi2s1jco3lORlz8Cf89/UfNWbam197Fy8//aKRZnIMrTkYmaTX7x1fPtNXRjZ4aHhQ8QjvI6/PsEsJPJjCB+6zGVPx+iiJPTg0qHwV25eo6qE9lOLIUDzelNen348HHxnpQwIVKr5wQEDuy9SnYlYYYIMgBxU9+FuyMSlDxedJ7A5HbsmCDoY5wWszRRt2LrYsD7afhbRWpYPXR0lidZ76mCxvjkGfM++be24LZ0eOxziSRaMG4LMsjFHzaHw+4XJC9iklwY0vmyTSNF8aRRWBQgQ92GbKdbJwLUYVDyoR/BdnVJTd/XW89Z0PoSxUgyf+8ov49C9NVcXIy4+rvvhdPPWlpSg8vw1f+vgX8d2DzqepZfjIA5/BX3x4NRYWjVB1MNyDmn0b8aN/egjf3WTpgem49Rs/xFOfnInkvho88b++jE8/VzPRykpyHK776tfx1ANLkTnciJ/95Z/ij35djK8/+218dXn6RX5j3h488Qo+/Ylv4mfVH/i1//YffvMGC1QkhiMJQcW4qCTBQSz+mXWiH51oj6+DCcn6xMPJPEanNSuoAQwmAirsrxJX2tFghU0XjXwj4bsTRXu6jIkDnN97UNhNhAUqnOuzlWcmHrBeGmPDO9v/ti9G+kVARUI/jbRvYqBi5PPxpb02fho5u6HKXawvfieggtIs4d8OVCxde10cXWYSg4CEkuN9fUj2cYNvEitcFKlpbVFl6hly0WH1ID+fNWuWEipa1ClFlBVEqgNUiJ3hmHAfOXAQHWOAClZyz503HzG3GxnZQcec0lAIlcig3IU0xgdkVmp9L2xlJxO/mmfiOoU0cjSSGAwWrDQCF8/BAVM5yQSkMZ0ybBK+jM5hBHnZWTh0+BDS0wKqbufizkqSpiYmRLzIzy9EbW2NmAE0BidQQWbC7FlzJPeUTWPY3CxkZudocZPutCP9ZIEKJjopu8HkpWVUaDFlv8rE2i09a/YtE+F8UbKBvhQDfb1IYpV8SzOaLzRKO5w64qeOHcFgeycWlE/GgunlyEyjlwif4gh8LrIeqEXpUYUqk/CqVOVGgxWRyQElvCj9RCkTVgrTUJtVFnxkpUfJFwNLGa564KZEFD0tfB54ooCXmWj2oyuKlv4e7Np/EO9u2o627gFMn1eJ9XfcAW9yEjxJPvi8bgVpDJoIVFD6icbMZMckp6QaRgVBDU9Mpu5Vp2kmNoRd23YhJ7sAt9x2J0rKygwXxh1FShqDNEq2hARUNNP0dnhYutlK7DGo8nsljeByedHR1o7HH34YX/vqV7Bo6SIMRIZlMstnkRI9iUBFV0+3zLQ53hiwEHRg4D97zlx4kgl+9Esuiv4YXZ2dCPXSo4IMhTBIOlmyeAnefuttLF2yRPJJ0voeDkkWiUDKiRMndE6a59IolnJe6SkpWLx4saqyOSN0dnYIsAhmZiI1K4jqs2dlpr1i6RIElEQyGz7uC3zpARw7eRzHDhzELddeL7CkfziEvMJidHd2o7enCwf37cHiRQQqJikZKr33UEj+G3PnzJfZPcegEvWIYvuObWJ30BSaMjd8UeueQMWs2TOM+RqALVveR3lZuUzla2qqEczKEFBRVFiEaMyFoyeqUDy5HM+/8Ev8+KGH4h4VdpPF4zJ4Tve7sWL5Mnzus5/VfWR7xKjSpspW+3gExFp5OG7COK7ZDxzrAioiw8gIZiA9PU2bTLK3tHmhHjJBOZdbm8yOzk5kZOXi/PkLYktVVi4UiGSZHEwx0qSd1fcDoX50dXWio73NJIIDAclW0NshiQbqBPlcNDlOgy85gKHhiDYLrEInYMjqKV4vte5PnjyGqqozYlMUTyrSHz6xqWlkW+U74EsMZ6tO6c/wcAg7dm7H0EAXFi6ci6lTp6KosBwFBZOx6b23sW//NmRl+rByxSXIysrFkWMn0draKa16juFZMydjzuwF6OyMYfuuvegPdWP2rGlITU5DVlYO5s2vVAKT/dDX16Pq8aJJeUjLCKK2tgk1VdVovdAkP5WcvBwUFher4njThlexaMlMFE0uQQSpCA2loW/QhTNV1VhcuRiRGCV6zmDftt9gwSzKXk3CsDsNaRklaO/uhy8pCJ83C4M9Azi4m3rnO9ET6kDMa+bbvPw8VXGTsWb8j9Jk6p2eHMZll1+B1t4AGju98CWnIhoZQEYg4DAqXGhpvoADB/bg+PHDKJmUh8WLF8Hv8wiw6OvuRP25GrQ0NaGfrICUVBQUFiM7twApgQwkBzJkls0xn56eIe1bblYIVHBO53zNZAHXGFYyk81AqR0LVPCZiUs/pQaUEOM6a5lq3FjFom5091mgYngcUEHw0nhCJGl95frMtZHsSK5h1CDmGsGkgQUqUlIJ3JKNYYy4KfPE33CNbm/v0JrE98RA9Lj1/BpJR8NX6g8NIRrzoqW1Q6Ay5QOHhwYRdZvkNuMA/pYbUSZNWL1NSTvDDDAycHbjrzUniaC32aTyeuxmmjITY4EKVePSLyscHiX9lAhU0D+Cc1Z37wCaW1uMJ4UjEWc3pWOBCgtWcO26cI5AxYDYFPzDNkuicTiGvosAFXzOe7vZ9qFRQIU24j6aUXNe9MWBCgL/lHZRgQATHBHOPxGEo4R7Io5HxQijgnMfKwjZn8QuLFDBVKAtqrnQ1KjPM4IG9KQ0p+KbfyVQwWpuD6WfCFQMmISO7pO8UkyyS4UdDmBKRkWQcUoKDe2jBjTvMGbaBCqYnPL6TLEIpa4ou8IXGRVisk5gpp0oVWVC6X/n2N+JU37vvcPojdHFD/P/GlDxAdc9UTL69+mf0eK+o3Y/H9BPCbughKRxfM85itl48cNcHAgZaZWLUmRM5NHTzknwmoR/4q9Nstv6anFc2yKEcV/TAHXY6zZhn3AoPqP2NXoUJ5hfjbqkiyXOR78/0Y7UxN+JfX4RD8dRl5qQ4ndbc1i7hxWCYBRcx/SQye6PuQarvsD5XTw78x234/GoOeoiN8my3Nh6FZc422GbtDTxmrkec+rR0ET8qic6iU0sOga4Y+/2BLITOtyIPIzZa8oUV+PHmO/yPa4ZhjFrksZKkvOeu4DyGRW46Y/vQGgghEM79uozGldTpur9N9+T7I8FCuway2MyOaomj532pKTrvBm/fIO82Epxu27yOFamWZJKKt4x/WfNiBmr6jQOkM3/Nol4U3luZRm1ZjvJd+svYBOx3FPxZRQJTJ/EGcwJaR+NIbXdfG6fJ2Og7ORZ4gle9jVBH647Brixv2G8zn2nfAEcUGQcUOEMkgkBC8cv1SSojb+AwBCuvw7bkmuxvQ7jXWCY14zjeE+417fxGXMGFgiyAI+UhsbIzbJJZCxwP8c4ZWyi3UpfsQ9VLOjIeDIBz2OxDQIqbroG7/7qTQEVXIcZ2xHAYc6D5+c5DLuKvpoGNNHYdBvgVTESpTTlqWDAV67BTKKbAcfojk8uwQSTG+Eej2OS8yDf4HkI1nDs828VnHg9+MGDI88kpZ8SpdNsYa8BzJwYUOCv42VB1z6HucH2WNkl7vfZH7xW7uviWUvmHRzg2D7WZN8zvtDYctHvi+CSk8dzfCgYc9i+MmPSxE7GEJs5ByP9ZHzjyKoYAX5G5tcR+Sd5WcQMsGbiMsq9muK1uPl23KScoPew8gzsN6p9/JdmVPzeQEXpKnz1G3+Jv1pXDCmwh3rQ2TWEQa8fhdkOmNB+GA/+7TfwwIsEJBKACgCde5/Bpz/7PfyybnywkLz8HrzwgwdwXSmj0AmACnuuCeKMzuNv4Gt/OfFxLx6W/Pf7ZASo+N0C91HftsFzfKEf+VTrv7MQjt8cjE2bKzozptKjXvZ4ZlEa95k9b/yjkbS7iRcNjWGcGfVEQEUiqDEqcrtoyHqRQcNp2VR/6NzOpY001QS66hMVhYxUcjjIgVnwx7YxYaOiNF1iIGvQjATWxkVDT9NmrX62SxMAEufM5vjmui0QZOt2TJDCBctMqlzMuLgNho0nQ3+IUk+D+jsu/cSk/+Agll1zvSZcLiJMINhKRib6fW6XNuV8nxXGZFRwolalgIvViX60trbqD7X3+VsT/EWUuONvLKOCCxMXPjIqqGduGRU00xZQMX+BEuKsUJFRs5L1Li1MTBDSVNpoa5tqAWvorUSiEyj3DwzofFyI2H4mCkQ9dAJqJjWpccyFzwAVhllhtDPJqCBI04fszCCOHjmsqmQaVVPWgIsapRAoUTRpUinq68+pIp7kSeqZRsIRzJo1W/4KmTk5ooumBTNVyWArJf30xkhKkrwKF05W2LKPGFgw6DTBjTEw5qJK7wNW9/I+cWwxOT7Q26X+jlKGY5BtTVNiu6+3C4f27UUALiybNQ3TiguRQiaFL4ZIbAjJngA8LlPZyQCV8kY0gObL72X1Y7KAHRrD6o+XMio+jTU+D7YyQRWprAJlYE8gg8bArFaNxuAjq4LySJ4YusMh1NQ14L0tO3D0TA386dm49xOfRGp2Jtw+L/x+Q/MOpKTKTJv9yj8EFZiM5LjzuKKSfYoMh2SmzUTZ7h27VT1+0623yxw6yoDUHUUgNVmBk8yZIxG0NDXrWNRm5/jhDEC6aW8vQR832tva8eSjj+Brf/VVLF6yCP0OUMFnaSKggh4VNtH1zjvvaIzxfnsDSao8pUdFeDCEro4OmWor1JEfRwzLli7Dhg0bxKiYVmFo/ExU8X8cD4cPHUJ2ZpaheQ+FUV97DpHQIJYtW4ai4mLk5eYqMGpqakJPby+y8plQP4/a6mqsumS5gIphMiok3+SGLy0FR08cw4mDh3HrdTdoaol4XcjKyUNHe4c01jlWrPQTt5wMXVkBsmnzZixetFRsHwtUcN4ho6K4uEgeFZR+MuBJF1pamjBr9nTDiKA8xI5dkjEKBNJwtroKefk5Gms0H+foOH76LHLyivHcz3+BH//oQc0ldiNoNwwcowQqrrh0Ne655x49w+Xl5XEvl3BkUIE5xyGfWUowcHwygZvsS4KHptasOmNSkFJa2ZlieLm9HgyIkRVWX3EToCrvcFgeJFk5uThXV4dz585h9apVSEun/JZH329rPS8ZFD6nPT2dmi+YLOV3hJV5XKriF707SpYSgcFkePzJCKtqMSp/GLaZwAiBCyb6WlubcKbqtOS5+vt7DTMjNQWlk6eguKRM8wHngHO1Ndi86T2cb2jQxsTvjWBB5WxUVExFQUE5Bcvw9luvo629HqtWzBegW1ZWIfmX1vYONJ5vxJmqM7ji0pXIzipCc9Mgtu/eD7cvgnlzZ8FNj4XUDCxddgl8vhRVRp46dRLtHc0IZgZQVFqGlPQChJiIr67C2dMnJSF2obVFTDRfdBBTphagfGYZ8gopRZGOnj4CFTWopPzUYD8am87g5MHNmFlWgJLSMhw4VoXSshKUTC5D/xCZc/TdGcLxQzuQ5O1ERmY+Tlc1oq6uGrFYCDnZaSgoyEJaWgpS0yj/1IesNBcWLFiCC10EKnxISc1EOMzkKo20PQIk9+7ZherqUygtLcCKlUslk9bS3IRwaEA+FJxT0wg2ZQSRWzQVkagHUbcHSYE0pGZkwZ+cqnRMZlqqtP65kTU+EzEBXfQ84iadQBTXQEo/TQhUOB4Vhh3FijdKnfFZ8qKrt0dgBZPYiYwKAmRcf7lWMDnMe28ZFTQPZmKO45ggvhlbhlERSEvVukZQhGsliww41slmIFDBJS83NweBQKo2XnwG+FJzqN87xE2jF83NbRqnqUlJ6OvpRPdAm+ZXJd993PyTScJkvAdpKRmjNumGau8xYB/XdGdzboEKtltABZNCoA6wYVTwxeo5JklSU5O1xkqb2KkWZB+LUeF2o6t3QM8u2SBjgQoC3RYksNR98x0Pzp/juOVa40dKIEkbV8oPkIHQHzKMCppnc55obGhQBGGAii4B5pZR4fGaZL18KOBFLOKJAxU00yYwQABJVaMRzs8EKuhS4QAVfq+kvqRnzCQPk1Iy1DZ+Y0owx0zFLMNNARXRGDKDNEEn8GHkUX4bUMEblRpIVnsEVAyEJINogQpb7WyYLl55nzDeoqdJRipZcQHNYYwn6VHBsWikn8hcZbVh0ijpp3CbG0k+P7yKM3waY+x3Y1w5Gpz4DwEqRmWcE7YF/15Miw/anlpUaex3PoBRYYtlxh/2d9zrXJTN8Tsex9lpjGvPBMlV853xCfj4TjEuV2va4OT9R7uWjjrRB7R1outzZGXGJi4vtotm7G2fJ35H85kTC9PYfqLEtinAsu23Rx5dvp94PitCOdEw0bkTh2T8v0f6ZzQgMfoo8bOTmTW2tYmM/zHdaErIHADCtsCCOWPbYyvynH2s2Rg7X3IMsQ2Dggk/Mz+NBRjGXrthozpAhVP7Z/vVFhAmVrCPqli36gEaaXYv7ySMnU4w/Wr29/G9vZPwjA+8+CU4AI2YB+Y69HuuU0yCOklVk7R15Gu473GYC0pYuj3yFVh+1UrQ9FuV6P0DMkem6Tj3s/JCkxQf53KzHnFdM1iMAfRtlbydF01mxdH5Z77GuT791mkXfytPKentO8AATYotwMTjO8l0rj+qcg+HTSJdRsCmJnWEUeQRmzMO2CUwCfh8aK2HYRhz/YuDCw6TiefiZ9y3qcjdAQxHphEzeNhn1qxZa458lFg4ZOODYZNYj7LIyPSxmDtObkbMHG5oHGN2m/vQvl/+AA4rW98xiR5VunPM6BiGBSjQhWdl0lpAlAMAOKwOm7BnXxG0J0vEeCwMqz02X2SAFa85hnIPBhAxeQf2gzm+rt1j5ICs+gPXUs47usUx4LqP3IQ1N63De6++LaBCe2ALODjJcuZ1eA4m4zWeKHnpI3Nh0GSGHNUE7oX5XSbXWQwoRQufKSLgb/3JfgyTjemwY9g14SEzLhlrMTfAwjWOM8bRvOKHHzX5Ar7up/STo/ai63OOY58jAZBeI4kkQ215YTjm1iDIZiREJY/kYiGHR0oThsVkxhnvm2E/sJBkBFgU8MRxFKPEkhlzdg4yOTfHe9eZBAjYsB0qaHOYdCzi4ffI9LDrRhzYNrt3XacYJk6NJvM0hlHDYiUjl2WfXwJ5fKn42QERNZ/8V5Z++r2AijNl+Pg3vo7v3T0TyejBiV8/gwf+9xPYKNDBj4V3/xn+z5duwlVkWdRtw5e++DV8932MMCr4teE2vP5PX8Od390DDvuRVxk+/t2/x/fuLjMAyARAxYV3H8KHP/0EdvxBXmpUz/0u//jmDdQCnUiO6CJHsSwB+/FvqUwyQEUCDD4mkhsNHlhkfwKgItF8eoJgSBNYAlAx0noTHOgz5wv6t4PEj7pKVe1OFDTahP0EwexFr3/Ey8Fsikzj4owKC4jEf+9sEBP6Z8S7Y4Lw13bVuO9bjwrHxDvxAhPaYd6eCMiIh/qSzhAVN7FXJpJ+YmUgDazle0D5J5pph0bMtAcGpLlv5KAGsWjNWi3YA4ODkm5i0skabA6HQkrIMJlIbwZLfeO/OfmzGpQV5PUN9ViwoBLdjvY2FxAyKpiE54vVkUygcDN/aN8Bw6goLMSk0lIluWn4SKCCQWJqMENJRhOUkcY5pGpnaQDGaMDm16bYaB5ajUCWCgEEKlhxTb1on98rKR1bUSEgIhTCwGBIC4kJKLjQe5Wm5cBk0pNSLj6PB1VVVcjJyjImn5SjYDJSDJIm+UPU1lRLI5FV8LVVtYgNRzFj5mxJP2Xl5iKnqACB9DQlX1jwwEeVC64BKphMH1b/8PfyzggbCRzj/WAkbriwMynDin0usEOhAXR3dcgQOiczW7JIPr8Lu3ZuVhJ/347dKMnJxKJpU1GUmQ6/gBhWQ7iR4vMKqGCihn3HJJEBeVxI9tLENFmVDfLRSGHyyqdAQxCO81wwOJW0g8P4YDLPReoxpS3YpzBB17ArhhDNqXv7sPfQUWzavgttfQO4+c67MXX2bMklMTDhdROkoCRWW1sH2traxIrJCGYq8HJFh6UqxWs7ffKYAuQ9O/cgP68Y62+6DWUVTMQyGoxK0oL9xY0Cg1ZKO5GdwASdMdOOKaih2SLve0dbG37y6KP4/772N5i3YB7CsajMtBnYyWCLVUS8VrjQ3dsblxfhuNq4kYwKr7TrfSnJArAovzQ0MCCggoarqgahqgeiWHHJCry54U0sX7ocFVOnilERc3OTaSiuB/YfRMkkmlRTfqkfDbV18LmApUuXagZktX1hQaGCTRr1BrOCAmSaLpzHtPIynZtAhZg/EcCfkYqjx4/hxKHDYlTopvi9yMrMVvUxA8KDe/dg+aJKeVTEXHoCEBoKY/PmzViyZNkooILjfteunSgqzsUkSkKBlUdetHe2oaX1AmbPMlrgnMO2bduBadNnSPrpzJlTKKCckc8jc25GfJQCy8orxvMv/hI//tEIoyKR7sswMS3Ji6suvxQfu/dePZcEeBjYcz5gco59ZzxbSC0mi8Kt54pABadJSW9pHhwSUEHjZFZ1D5Ju7VTL2fvMJC3ZBpSpot49QYFFixfqGSWrgJsasiA4H5H9Q613zkN8XgiSiHUkD4JUU20W5ehhUi4Jbo9fxsXcuFjvB5qni1budqG5tRkN9XWYNq1C4GrThQuaW9juYHaaroFJ7+amZmkT0yuBIFtnRwcmlWQjOzsD7a3dkndqa23GjJmTsbByHg4cPIKeviHMX1ApY+yG+mo0NzXgmmuuQWTYj/q6Duw/eBhZuWlYuHAREGUVWwjLli9Fkj8Ij4eG751o72xG1Vl6jaRiSvl05GRmwefySHe3pbkV1TXnsHfPXvR1tSCQ7kZuYRAlU8oQzCpBLBZAY2MLppQUIxQZRiQ6iL3b30ZBZjLmzVuA3QeP42zdaVx55eUomTIDHe0hySkdO7QPqQEXZsxcjKHhAM43tqD67GnU1Z/EUKgd+flZKCosRDAzCTmZHmTnFCEUKUD3YBC+QDqGIyEEkgJoa23F4UMHcL7xHGbOmIJp00oxFB4Q2EPWA+8npfwml05BMCMLHZ3d8AeCAvvonZRCBkdaUPJdfGWmp2peIPDZ29One6okLBPyBNfS07Re8hmtrq7G9OnTdb9MzBEzjBrKFTlAhTY6kj1wa+7p7uuJSwOQncD1y+M2/jT8LTfwjJc4D3Be6qJ3kdcjgJljny8BFX19IKOCGyW2h+Oczx/XFgEVbR1a72hOm5HBNc6PQa5JYIU943uz9jJG43g833AO3Z0daKg/h46uJlMs4OV1u7XppgQYY4PikinIyMhUElvMJocWz/XGXiufD0pPUYZRUogEKpjcAKURk5QQ4drPdY8JDYJSbptk4AYwFBL4QmNrrt3dPX0CuPU8+o3skCrgBPgblgjXeibNrQQkP2uob9EaQ4CQjApta1g96XJLapEgejBI6Sc3Ghsb1Ze8xp4eesGEBVSQZWBYBV4xBL3eZD2HFy40obu7U/dM0k/yl/Ii7MiKKM0R4/X7BeIyEUTGEfuG0wf7ntcujEJVqB64NKfEBFRwbcnMSDca0KpCNMlCJems8TjjJ7HcXKg7d06/5bxF1g9BHRausJoxkfnCPlDlrqSfktDV2YWeBEYF4xIWnLS3tsblrsSoIFCRkmzmWEcawwIVBPGYDGDRg63gVUIlIVb/jwEqLrZn+qAk+G/ZrSVkQE2iauLvj01Ej6qMmqDk/OLYyQeBCxOd3HjhjNpmJBxi4uZOfI4POrNDqIyfxihUjfdYMOdzqtUTC5HIDeoAACAASURBVNic71+8t8dLGsU3PhP+aGSfOCrxbRNOzsdKgqupxpNOT5SeOSYhTaLJZLjH95RJZtlesRu+hF6y12f3ZCYnOvpe2Ir8Cc9gzz3+AiesHOezOvZe2yjMCi0k3kTJxZh9ztjX2Cs2fTjxawQkMd+w99gAVcwmXuyZMMldSc1KhsgyxkzC0MzZ9FgzUnimTeaOGdaKvYksvDL3T0lCh03AvY2V6jFFKua+xiuqnap+uxZbEFiFag4L0LZcoHhCxbwSowl+aAIJZKrr0T7NygsZHwYNqvgw0p6JCWptAg0wwb25KrQdKSH5QzkgiPqQiVpWoKti3AARcaaF00g7Juzcaav++bGK3By/Rf6eBTx2XRVg7jAYxFiwPesAIrxuk54xAI6RjDJyTYxFjdwq5VSNdJF9vvkZ4wwrd6RxkDAOzXNnxgjPYWN2w1QxhZb2Ze+dKvmd4gbTVtMnFlyXDJZ8Js0oNP3ogGascnd85rS+Cow0Ej0WPBBQIhZCWDENizZMMSuT9g6Twva3GKcsahyGz5+kIhkVPTiLAI/B8ymxz5wCK/FlaM04xKVCEAFgjgyTkbqi9JCVPjPMEsYL7R3tKryzMkN6Jlg2wvM7DBCzhpo8iXmWzDUydlDs5TWytmL9xpkEJlblfljjW/1r8gzGi8IwIZhrsf6iZvwxHonikcdGgIr77qO8sSmoNEbSBCIMABs3rU4yIILJtRD8M/EVv29Z8LYgVfc8RnDDMJt4PMNeHtJ94d7PyjXx9xw/KjxVDGfkz3gOjgnlNZwpQ2PITXAtrLiG16KSOpdbxT2G3WJ8JQwQZ/vT9JtmIubeHAaWWBSOzDCfZwPc2efZtNsytTRm/wBUjJZ++uXkB/D0P9yDFRlDOPHrh3D/F58ZBxqU3fgAnv72PViRPYQTL34HH/7CRsy20k/OAzl45k186fPfwIMHTaUOX/qdju288Qeg4iLL+L/t7W9db4AKvS4SBCeewabbzff/FT8QP0IZ14ufJnEDYWDrMRc19jyj/50YVI0HKyxQYWWQnGNrtfyg4479LDFoTGjexbrAou9OP1nQIV4hYyPvRIaEo7850lEJwenYvnZWe11CvA1OmBXvvzFgxTigwrnp8YA+UU7LOUECUGHLktSDDDyYunOCMy5WDIYGmQB3gAoBEyFWW44GKiYvqDQLc5jARkhJBlaW6nc9fdqscuJnwoV/CwQRUGGq45gUYVJm0aJF0jPW59GwKkzS09KNv0R/v0kOxoCD+/ajq71DQEVJaSncrJ6IxTB73nwt9GnBDLWHG2Im6Hl8TvxcwJVAd8ygzMJmqiu0IMQItgwoKchqfSYlaEbKhJ+tOCFQwSoBBn1coLTBl+SB2SRw4WPARX1RGhxnBoMKJnirWHWeLOkgGkx2o62tRW1KC6TjzIkzOv/M2XORmh5ETkE+MsnGCBi5DqM3bSpGpQ8ZGtR5sjKMPBYBJeotUhaCYJRNsLDdrOKmJBLbHh6iyS6DAR8KcoowHA5hYKANe/duRXdXG6qOnMS0kiLMnVyCnEAyktysaKVOvh9J3qgSQUwcGK1uytOw0oGG1T7RXjn0KLXFani20yMQiW0y2wRWm4par+N6BXoy6FP/KxlDCRRuHgyXnJWjNfWN2LBpC46ercaKK67E8suuhJsBntckwyg5xXPRn4KG5Qx0M4JZCA0NIMbg1wtVPhOoYHXxzu27kZOdj5tuvh3lFdMQ5rk8MaRnGAmtvt4+BVtM7jGhRaCCY0nVLj6/xpM7GkV7Wxsee+QRfOPrf4fZc2Yrt0xmhJKPTrUzgzf2HwEXml0z+GPfbXpvo8bNrNlzlNDp7OpCICUZITJ/CFT09JiZln0wHMbKVavw5ptvCrCgbj3NSt2uCGLRYRnQHz16HHPnzBXTg20mQ8bv9eDqq65SgMZ7nxJI0bUQSGSCiwbBne1tqnTlGCLNm+0LR4DkzHQcPXFcjIobr7lWAA07MpiWjqb2VgV3h/fvw/J581A6qRgRd4wkAAwMGOmnxYuXIC83TwlUyV25fNi5cxsKCjJQUlQEN1IAtx/N7U1obmnAvDmzTWAJFzZv3oryadMkI3T65Ank5QQlU0bPC7h9OEyPiuIpePGll/HjHz0cl36yQbKpeooiPcUnRsXH77tP88e0immqZOccxeCe8x3bZplatoLJSJQY3XYG+pREy87JRjAzw1TfRMIYcnT1Oddx/uAx6UGSkZmCs1VVOHnyOIqLCqXpzgo0JtqS/DQPNr4Hhnptgl1tHhzZmPSMdKN76lSscYzwOeMcwjmTMm8Ck4YcVofPg5a2FtTX12HGtOlirHGiOHu2Gjt2vI+GxrPa4DAJO2vWDEmBcR4+W1WNLVu2IyPoxdSKYuzfux/dHT2YM2sG8guzkJmVh+7eMCJRH+rrGuH3uXD4wHbkZKVg7brrEYkkoepMPXbt24XJZcVYtmwVEE1Be2cTli6rREpSPryedHR2tyE5LQnHjh3DmTMnUFychYK8AjGaUgOZQIwG8hE0NhIIqcKZqmNoaqlHBMOqRs/JLhRLIyczAwUlU9Db34vtW95Cqjeq9WIg4sarG96Sif3NN94oiaH6c7VobW5Bbk4WyirmwOXNQTSSgf7+MOrOn0Zj/Uk0NZ7D0GAv8vOSUFoaQHZODryeYnh9k+ALpIrw09cTwr69e+VNMWf2DBQX5aKpuV593dvViQx6UEybhZy8IqRl5GA44kJ9/Xl4k5OdXItJwnMu5D3nvCuWhoesrF5JyHE8cj41LDWXZOYSgYqZM2cK4LfJBCauOWblQ0MTbSaVlWwBenp7dFyOY85f9DdID6Yh2etGa2sb0tIoQcjKPYgtw2PSfNvj92ldsR5H8hDo7VXb+eJ/85wWMBFQ0dIhz4xgVhrS07IQQ5IYFC5vCGQIuIZ9ujbJjZ05hdMnjqKhoU4yYBGaMMqXwKwBBOoKCws1pkNMoGcRRCrC7NlzkZdXoLWBYLQAA23gycTqQWhoWABQcgr9W7jXGBbgYmQF3YaxEiH4lyIjaE4L5tkJC2xhMQXP393Tr3/zGaGHE2NbxhNiUshjxnjRiEEouUMjW1jf0KR5hP1IXxmTtDCJGZrA8vrF2nC5BDzxcz73XT2dYr2kUg4pmeC+kQdhtJacFEA4HBPYSRYU7yF9LVQV6fMKvDfxYQyuKNc+shgJEA4TizDSU5o/KKtA3x5TMOMmU4NLasyFC031ei+Ywes3SYZE/XceXeuxKncNy+1c3TklKSllR3NybvJZmCKPLyfRY6UulLQlUOEnKNOr9YjrBj1K2H8ce+1trRpzceknrwcpgWQBO0zM8BVuczng0P9jQMXFtmgXy8wm7n/+EwMVFwWDfkffDNNNE3SWCaJH9a7xOTD7GpOANclnm9S+uNzv7wZU2GObMN6p/NcW0+7ZbNLUVso6nlZMelppEMKBTMI6mvpjN+CcL81QcEA2R/s/8YINEOCANrIEGL0hTUzyT7hVvQhidbGhKQ+CCXbniZjQqI9HgS0jn4yBX+L7oYnOa9utggxHz16xnyOvwn3QRC/LiONnjKfYN/JDTGBWxJPOVoWac7LDBLCAKgFde7+Z+BX4oUp9ehCa5LI17rWyRZalYVIftq2OrwKlf53EqM3aK3Z0ZEZNMtYkT036wFFdcDpZ7H8l0J0kr+MhISaA47smXzWyFRwJJlaTK4Z0mBpWBknfcbw7VGjjyDNxTz0WqLBj3STGjU4+Y2HO49z7cp/DPR0VCSj/GGcPO5X+bK+KB5wxagF+9pX1jBMThCCSquON8bLJARg2glj1Tj+YwiwjKxUHFxKVMyyQaTbTcQlpm4xXMtspBhTg5DCetR4655N0q55PA8wbTwLxLQW+c6+sdd+R67KghFkTTZV+DxmmjPstwOQYQhvwxG8YHkxaOyCJ1CYIgDggBNsmBqoDmIi1wPccrw77t5XqYju5TnONNzJYJrfBvaV9JflV/q2cC+O2ltZmJCf7VdjImInnGgpZGS/uV0yhyP9l702g5DzLK+Fb+95dve+b1JJamyVZi3cbL2FLIBAgMyQZgsmEf5JzhhzmBMYEhpMAgWwznoQ/hGRCCAwEZiCYQPBuhI0X2ZItydq6pZbUi3rfu6u79qr/3Od536qvN0HyJzk5McVprK6u+tb3e9/nee5z77U+FwKCWMCC48F0/TN+kvtsZCEtaMZzFe8Iw14VUMU06Nnt2BjT+lBw9P/5n5drUv/p/1GZKWXB0/tEPSn4b+6TShSMaaxkmtRgBLR2Sz7LY2Q9gdeGY0ilvqjewGPRuowAbtmsxIXCLuH2RUKKEmTKmCGwwYHDxg5uh9ebeZ2NHzXmVEa7nWtYZ2GzoMxhZvzzeyXPH2FNEejS42M9S49JgS1txNZ6HmXK1PPEjk2VmbLPwE+AilUeFZ/CwLseVK+JyRP4+AcewGeeZrFk7asZ7/6jB/EXv9iJ4PBRfOBX/wDj7/qf+r3ZUYxHmtEYWMKpL/0h3vXAYxC3iupD+MjnPoFP3FUDLM5gPlyDONZLP/1jGBUf+eaT+MRt1/e3kDMYO4r33PgAvrbhEvhv581Pv2mHkfcxi30JkVYTLM1x7L/NE2NP/8cFKoSO6NzG6uK6BGKrUJINAg9buTRBqJP4sLYXY+PDWg1UrP6OE0Rx7tv5701Ctx8BVOhEZc+uTO/iNV3FmFgbMDpPohQFrgFoJIoxN8N5XUrDU/+4OmFYe8AmiJdNrQEqhENaJh/LxqzBG4EKIuGC4juln340UFG3bYdIRdiAg4tCOBKW4CS5rCZhnPgp3aKoucqpSH8D9daTSfT392PPnj3yNylY5DKIxStQFY+rfnWC3bdTIiMwPDiIXCpTAioo/cTle+fuPVJ89AX9WFikNjoXc5WOYADBRDgcrpDztFrVvBoW1adpKrvRmez7qJns94s2PY0vLbVWji2jjAoGbtL5ZgobHMNcDLlAjY+OCVjDgJryGqJv6CqKOSe3d214CNlsCoFQEAFvEBcvXBIz7Z279yIWr0J9YwPCVZViTK1AhSY5wlYQXe+MnEM1gYoQixsEKrLICaWUQZouivwMGRyzszMSdLLQQBAgmymgpqoO2VQKycQUnn/x+7g2dBWJiVn0dLaip6UZVSGCE+xqdYtmYsBHTf6gyFcEWFyjGbqYbeWle0cDY5q7+hAMRKTQKGwQKa4oQMGUgICE0FVZNDPMD+lgIGhBuShTeJPr6gaWkikcf/Usnnz2ebR2b8Pdb3gz3GQsmCILJaeikZjICE1OTkkQE6uIi9Ep2L3idSG9soRLFy9I1+pzP3wB8cpa/Nw7fh6dWyyjoohoRcR4mazIf9U0dk6Kv5TrUZDFKzr0BCrYbf1XBCo+9TvYtWuXnAu7ZIQWy+MzrBvpgF5KCFDhJ5PH48HR7z8lARHHrC8YFFCEHdBkVLDzOJlYMhJ3RQGgbr7lFjz66KO4/fbbBagQqRCfkLtx4cIFjI1NCFDB68+C5bXBYQHF7n7d62QMSEc/fTa4HFdVoaa6Ggvzc/LDcV5VWSH0X6EkuzwIVlXgQh+BirP46XtfL0lG0etGLBzFbGIB80vz6D1zBkd270FbawtyrjxclEVKpfD0089IQZxFRkqOiLYr3Dh27Hk0NsQEqPC6IsgXPZiam8LExDD27N6ldHu48exzz2NLdzdCoYgAFfW1MTk2moJzfJztu4y6lnZ869t/j89/9s/F3N4GkhI4mmk0FvIKUPHe975XwIwtXV0GqNBnhxwQBuo26LW6pCzg2Q5tBrT8qampBkEEmooXwTkxI2NEOr99PvH/OH/+AnIF9Y5gEsBCaCgQQjQcFSYErysTB6Wok3rN49BOpCIpytmcSJ/wHghQYYoyXpMM8NpSw53jxwKiLo9LmDrsWu+iMXw2iwvnL+DkyZMiQde1tUVYO5w8yDbisXZ0doj81vnzfejvP4WKSh/6LlxEU30zujo7cHXgEirjNWht24Yt22/AV770FQxc6cP8zDXcecdhHLn5dkxOLGNocBSXrvZj+65O3HjgCFyuMEZGB3HwxgOIRZrhdtFjgoVwFtaXcP7cKWzpqhZgLRyOifl2Raxaizt5CEuHsmJcC06ePIHR0UG43HlUVETQWFeHzu5dCFdUoO/cK0gvzuDwkcPwR+MYGJnHo489iWIujSMHb8ClvjNwI4vdO3ege9eNcIeasLhIY0I3VpKzcLmzINOv99XTuNJ/Ah7vNJqb6tDS3INYtA1B+g14chgZHkdf30U0NbWguroGI6PjGB0bE9bDFl7DllbU1DcCLh8yeYIFLgFcvMGQzLGcL5g00muF8nRMRulZxMSHRQAayXMM0IhRwDwU1wEV9G2ykksc105GBdcBWcJlGScYulgGKgoFKe5XVMYQ9ClQQX8MS4e3SSTNtwlUWINBjl3OE0zSyNbj+mYNFC1QQdmn2alZ0fatqCIgHUWxEJDue6+frKwicukiBq8O4MnHHsOV/j6kkgkxJOeaR7B4bfdmScogT/1lj7DzyACrr29AfUMjenbsRFt7O/z+kAAVcwuLyKQVqAgQWBQtbTIMFKjgM8L5m8UhyqCxr40v7d7Ly7PAa0mfrJWVNOYX5h1ABe+lFg7owc3jKTEqCNAL+0WBCn5Oi/ra+UjmIRNOC1RYM21KeVkPjMXlRWTyWVkfCVQok8ILSsZwzmOT6ejomMwpvGcqi8W10bMaqCgWxHycQIURplCdaK7vWdWZtowKAhRy/gQqJkdQyJFREZXijMyFhkFiJTI0obamrW4MDg5Kt+J1gQp2bRojSxZ6/IGQ+LCQJUsAjqw9yhuShbERUBEMUfopJkUyvn4CVDjyUsOoUjr5+tzlH8eo2Cjv3YDVYHvBNqV/bAIKbJJWb9pr7wAq1p6iCquWC71qeLw2z3TucONjKnWRr7mEzl9t17YtJOkca/ZVQgrIelQT1qzIr1Duh3Gt6qJv2CUoqdnGxWpn6mfPQuVhNs5T5djWnYPKD218Vze+GZsDFWY76za3WnLKbtU2aqkks4GbrsOqULkdBWWsKbamoxsbc/NvzKUkbzOygbaga9kUhkhQAgI4D0oRvWTUrPOKyASJhJSR8jEnIVIwwlpQNq0W0fVeWsDAmX/LfoVJo9rzNi+XNcH48umao8AGYzMBNITxvtakV9+zTAvGRDwG2zxj919iAphrYIu4sgZJB7nm77Jf05ltGR/2XpWGofmH5rBuYXzY3NY2w9jtyrm51INRivFG0oZFWGUpUCLIeBGskk8iaKFd+ozhZdyW2BoqaSXF4ZKcuFsactg0INdaQA7jRyJgpcoj8RylO17klJThobiHS46R/+Y6zfNRRQK9J9bnw0o1S5WEz3AmW27WMAbPcs/E0FkbE0TCyaeNTU4WhhbPFS2z94+AAnMD5l2W12NzDWEnGDki/tc2EsnYJKBkpJ8U8GEzmorAcR8c06KokOZ5KWOC22MOJN37cl0C8PnVGJr1CFu7sL6VYvZOMMKAMcpuVS8K3Yay6tS820htyZjWBinGQzwXMmgJVFjfEf6X+2bTlhbZeQ2CcqzC3PC48fnPl+tVv/ofjTSXMINU2UKeIwPGMV4mUMG/8RxE6cKrUrt8T2SfxKBeAQYdW6zJqVwVfydLM7mSKjFHFAw1fib6kMi9IMOFD2mZUcJGTG4/LxJWliUk/h4B+mMkjUxo2cRdfCOzGXkWhCll10s3RCJLx5rGnwpU6L8FLBI5trKEG2Mg8RjNZl4jjArvEgZOD2BcWd2rXxXN2N9TgyDNtH/9q6j6zd/DR26LYf65L+Ln3/95HJ3deHHr+fefwDd+7w3owQC++JsfwyP7/5sCFcNH8WcXduB++ltMnsBnPvAAPv50Gje//xP43791NzoDSzj29ecRf8sb0BNYD1SkxvpwarjMwtC9pzE3dAJ/9ukv4pGx9cfT+esP4ocfvhWNyrze5JVB79f/K/Z+8PnrfejfxN8+/SYroaGns5qR4Oh7sK0qptNZPvtjXgHb4bJq4XN6ctsiu/2AUM7XvEpSSQ4mhI1wSsX01R0lpeYWs9ibypaGkauitrVAxfpiPvkDG70sbW+jvymeqtdJggL+UgrkDIjguIqrAuk1TAvdjgWT9L9WwXQdEOHcR+kr9jvXu3NKyywPBLOHkmSlBnFa6FCqqQ0CaDLESVnNtFX6aTNGRfOuPbILLkgsuFodQQlyjO2G9afQTmKVMZG/MbBg0ai3F93d3aXCIfdPeRoW+1i8mhwbl+ICu8FXEglyllcBFexI3rajR9gO7BLlIk2NfBYKuDBJ52EoKBr3NnCyi58UHoxPBTsE2W3g97ul6MHiJIEFq+vJxdhKZFB2QhIfCUQ1gJcO7HwOo9dGsbOnR3SyFxcTJUaFq0h98GUkVxLCqKC8RiFbxKXefvjcXuzo2Y3KGhrMNiHIQkIwWDK+IhjGQMAyKpxABTsfec3E0swYADOoYLGG8kU8P0pNcPFLpelNkRFPg1wqicGBPvkZ6L+IxMwsdne1o7u5AfGAT4oL0hXg5VjKa0d4OCTa1CJFReNLdjW4IJIujC0YaBI4iFfGtTODnawi3cCAzyudoW6PT+mzpqvBAhUs5koRC+wioSyUBwz1Lo+M4W+/9yiClVV489veDln2HUBFRSwucigWqIhEK1Sv0kg/URv98sVeKeo8+8PnpED6rp//BXR0bQHVTVloEqAil5cuUWFWLC/LeKaPgHTtyLG6S0AFgYe/+su/xO9+6hPYtXuXTLZk8IiWpwEqRCbL45HCGscvi4v8/amnnpTz3LV7jxTaqJEuQEWKQMU8UomEFC5J1GKwcuTmmwSouOOOOwSo4HdDQTKSinjhhWNyD7q6qOufFzPewSsDCAV8uOfuu+VcJMA0WpqTk5NaRA8GBERkTtZYV4/qqrgwdTiWQvEKnL/Yh77TZ/Dme35Kgue8G4gEw0ikkxibmsCV3l4c3r0HLc2NKHiKzAwkgBOg4sAhKe4SoJAuGbcHL71ERoUBKtxR6UCfWZjB6MigeBxoV50Lx0+8jK3btwsQdrH3AlpbqiXws0DFub4rqGlqwbe+/T187o8JVNDAXpOXUvLociEcJFBzB37lvfcLo4Km0exy5vhkcMpEmfeJ8w/viQVyquKVUvjkc8QgmMlKVXUVYuyG97HkSfAiJ+fKezo2Oib75meiFWENrLMF1FbXIxqKijE2wbmMFD81+KXWK/fH+8WEIZ/JSSG3oqJSVgIWGqUznN3KPgXECVSw41iShFRKEwSR4pnFhfPnBQgbvDoorLD2llYcOnwYW7Zt1efITcmVNAYHBnDx4kUZh5GwD+cuvIxsdgnxijgO7DsixekTLx/D+PgUtm7bjZ96/dvw1BPfx8snXsC1wfP4+Xf9DHbtPoC+iyO40j+AiZlJ7LphK/bu2YdiIYjhkas4eHA/KmNtcLvCWFpOiOTTykoefb3nsXVrrciZXbrYJ4lQZ0enMAY4e4oYQ8GHxEISly9dxFNPPYyx8X6gmBQGkDsQQ1NrB4qZJJBL4NZbb0GsrhGTcz7MTC/iiUf/DvnUHIq5JdRWhXD44D507j6ItKsGmUwMmbxXfHhYuI6FYpidmMDx5x/GtbHjyGfmEfRVoKmhC13bWhCKsjO2gKWlFYyOT2NsnOa/cXR0bsfWrTvgdqvmdAEe9F8dwsjYJLZu24FCwYVwLK4+AXlK5YRlLiSrgutOLExdfnqJrBigIg2fR+WK2PXvZFRQrssyKmyXmgUqrDk2111JotwekX5ax6ioiCLgdYm0EccWk1VS8EtARWpF5mMmv5aJwXmPQAXnCL6scXdTE03aIWN+enIWHp8b8eoKAQ/cRfooQYAKgkszEzN46skn8crxl0TGLrWckGc4n2cix3GrUgRWykLlqwgdZuVtKXSLHrJLgBx6Or3xp9+MLVu2IRiOYmp6FtkstZOVUZGnfFGRjL8yUMH1gDFWJEzWk2HiGjFnAjc8Z0ny0zmRhqTmMpkAnHOlACX0f/0vjz0UCEqxhYwKvjcyOmUKDizAGF1mv56HE6jgNbs2PCxrINfL5WQC6WwascpKmfMDPt0+F9RIhJ4WPgwNDWNmZroEVEjn6hqgwl0kIEqpRWVz5Cj5xK7cgsoX5LIqAyVxqOkwJVAxMTUqXd+VMRpX+yVWsjGbLeQq+KJFC/YxDgwOSlzDOXAzRkWpC9PI4BBsIlBBac+KaEyeYTZ3UFpsZnpKrr94VAgQRI8Kv8Rb6tXxrxio2BwV2JAosCqXcDAqTLViwzzExpOlP1qgQqP19enUJn1XP/qA1iVmpYajUuqw6bbtJzb5wPWuk01L1u1+421Jyd5UokuNYtc5rrX5neRB1shZCqCrd/zjABWSaZlueAl+TRGa8RSZxgQVpat8E6BCUt5SV73J25wGxqbDXNNnsrq0ALfZa2PT6U2Aik22s5n0U2ncrGF9OLNO53GtBSrM5ZaPbHYOAhRYP4wSy8AwSjY46bKZu+asVqbOuY+ywoHGTPIcmX1YcFwAEin6KhtOjt10dYtHm+laL41/k7s7AazSyBfpFgU4bKHUggfCJrDG36ZuYAvcUnzf6GXGg2VwcD4XgEYAaC0kK4NHz43Hrv4PvlIuL8NMJ375m3bNs9BcauZ2TAs6Xng8IqfFcWd8K/gXey4y1oWNmJY5XGJcI/Fkr7+NUfi7sJuN1JA0J4ofBzv5y/U9OS7K6BivDltstsVwkWMqaPFYmglFU1LvPAv6UvjPGINosjnpiyC5RpmlIYVhyiDy2hk/ABkXpjFTb4FeA+5DvD+EUaCsPisFJUXknAIVHB8EhERVwEcZJGWhqGSVsnHkEeZ9Ej9OlXTiGm9lm2iSrA15em76Bb0PyvpQpocaUWs8xH8I2KUXXNgBjNWsR6VlfHB9ZQOTeDOwu1AkKXleWvjhfeZ29XoSHNGmDAVlFLCw912bd3CjCgAAIABJREFUETXGFMklh5cJ7x3rAjw/y2qwMk/cDtmUXMuFIW6Mtf/yC2UWyK/+qoIwIoclbCKVrFSWgQHtzD7svMrjZNOmAjUchypZpWOH41eBK95rxrhk6/JxF6BKwDB9Ju244ENBGTg9N2WO8EaoZ0dGGshkXBNMM2bYBE9kS8Z7UNgP0mylTSsWSNH8zHihGAlRC1SwWY331Taq2fhLARszyxKU47zympB+KkuCbTwx8l0CFR/6Bro+9Pv4tX1+DDxCSadv4tQmXhGNr/8AvvHZX8TN4Rk89MmP4mvtH1Sg4upRfOAzA3j7p+7H3fXAwCN/gv/w36fxvj/+GO7f7cf86W/iw3/tx3/51Fs3BCo2PcCrR/H+9z2AL/Zu/InrgxWvHZCCV+fTb9pm5jxb0d78tpem6HX+Ctf/Dlf+EqawWZeN8/117NLVBfp1EMkmQIWuKRZd1g4CScNKXUbOIM0AB3YRsKckH9lIjsp8YNPzWUPbLQWsdsNOpMa8p2uq42V/WX+ccmqOz5YZKc4NrAFcHPJb5Z3Yz6z9nnHlMgCN7Yux91E6MYyhtmVUZPIEKrR72PpRrKTTKqckPhUpJNNp9Nx8uxRzuY1ZMdqclUIHi2lsD7TFWtudweIgfxiAKSUvK8Uzyj/YojCLbVxAWOinFwATZnYTc1G+NjSM5cUlNDY1SZclGRUsrsaMOaYvFBD5CKL5fLFgzgIBgyw2KjNQ5QKgC6gGBDxGLoAsIEmHgU+Biso4i9QKVPBlgQrefsp5SIHUJFAS5OZycg3SyZToiycTNPFOwMdObMrN5LMif8HCyaVLfQIeUDOo71yfsBS6t+9EZXUN6urrEK2tlMIJWRQSUOTZAe6XAg7ZEww6YqGwMCqEJUIdSPEXoVGrAhSUYWLBiQUs6UApkh6awcriklyXhZlJvHryOJoaa/D0U08it7KMHe1t2NbcgMqgT7rtRX+RXd4Uzy4WJTBTQ2ntROE1oQlwVbwCdfWNCLN45A+iMlKBcCgkQZNoQLJz3DCxvD4FXETCyXQfSGGE3eaGUcHveAI+8bAYnZsXoGIxncFb3/XvZBTTUJvXn4Ezu5bJXGHSyAIwO22ZiFAayesqYmlxVsy0a6vj+MH3f4BIpArvfNe/R8eWrcgyOPAA4Yh2wLDwzWNggY6m45TvYBBKNgXPWYy18znMTE3ir7/wV/jUJ38HO3ftEuCEjAp+VrwpDPWX42tucREz0wpU8PcnnnhcZLN27d2DAKm6U1OS7BazWSwtzGNpfl4KV6Slcns33XwzHn/icdx+2+3o7OyUADBEuRFXEY888ggaGmhS3SyFb45hdjP7vW781H33yTkpgJaXwik7ogk8stAeCvgRr6xAW1uL/JfHSEmrps52XLp6GWeOvyKMCn8wiDwNcf1hLKVTmJ6fwuXeXhzY0YPWpkYUvOL/LMf6zNPPYu/efSIVI4bqAjy58OLxF9BQH0W7mGkHUSh6RPppYmIEN+zaKQE4x/iLx09g77598t2zZ06js61BgtH2tnYxaT/T24+axhZ86+++h//3wT8VAzf7PNsAW2RKQl7c+7q78L73vU/MyQmEklnBY2TRjZ/lvECwxhaPuZbEqGlv1jjpaqSMVCyCmpoauD1FMf9mEZkFW8rptLa2aPdNISdsI85/w0MjuPnIrYiEoiqPBjfSBUopaWcSxzyPm4kLn2dKTTF5iVfQ36Aox6h6yy54/ZTj4ryREoYXgVUCLbyn3NepUydx/KXjMkfs2bULr7vrLknYhGkk0nWaiEgxkwBNoYi+3gs4c5LSUJcQqwxh/76D2L37sHRJLSxM45mjT2NkdEYK87W19fLe4OWzuOd1N2Hrth6cPXsVgwMjGJ0cQ8+eLdjStQ3Xrs1geWUWd951BI0N3XAhLKBZMBJFLuvD8OAQvO4MurZ0iOH31SuXMTU9gfb2NpnLfcEo8lk3cski+vr6cPKVFzA4eB5btjRidOgiJuZWkMl7EAsF0FRXgcM3HURdWxfmFmOYnU0gGnLjr//XnyDoTaO1KY5DB/ciUN2K5RwNy9uQL4YwvzyPSDiGWLASC5MzOHX8MTQ15dDeVomnHj2KoatjCFd6sW1HO1qaW+V54fqSzXtRUdEAv5fF/gAmZ8Zw5eoA+q8OYmp6AbX1zTh05Ba5zwFKR0l3pEued4IUBCs4YUfDIZkXeC/JqGBS6fVQXoGSAQVUxmICuNLTgF3sllGhIF5R1j/+2xpca4GaAZYbS4mErLv2GQgFQ6isqgAdlMg241hlMsflamU5KUkUQX3xqKBBpkgLqNE25xCeu2VUcHwTUOL+2DgwNTUjQEVNbRUCgTAC3gpZF65cOYsLvacQCQZEfuvcmTOYnhhHKqkm9cJMk7yvrMVrE0dlHSolX2MGzqGM81gwB+oaG3Hw8BEcOnREwJFMJg9/KFzqLOR14VpAlgDHO8EcJsKxaMSYTeo+eQ5jY2OS6HI9pYwb50T6U9CDxilrSuknO4+HVwEV3pL0k2zHzw46wbFlruK6z9iFawf3R48HJrM8r5X0CpKZJGIVClRwnpbzlZiCLIcQBgcGMTU1iSg9TsRbxCeMvQybEKS4QbNKNW0l+C5eO2kyIxQgYwJMoMLWJ8kDk//lCpicHpNiFJlKjHFKxUrTach7Iyw4UdCjHCgwODwswC1jKrLDAvTqoV8XvU7MNbVJusRU4lEREilE8QOJRIwEnk/G/PTUpGxLWCjiJ0b5LD+qquIlRkVmGv8qpZ+ssenaLGltO9Sqv2+UVxgpo42yrY2BCn5yM6bAZjkbQaqN/7ZZt/7qpq9yUX/dMTlSn83OYaP3tRS0wct2fq2ttbOA5+AWKFBhMpdNMZL1kkaaP252ncrva0HclMINsOns1tfDVB1+fo5sKc7LbIySd+ShW3+GtnAuH7KsfKO3X87aNI80me26wy1lkGvMtEtHv0n+urb4rp+XMve6C2IyZ/OR1Qyb6wEndk5ff4U3A09YZdRmSru+2c74je6SFOqNzBw/Z2WZbF6p196cFw2PychmfmaKpPL0mGK/Kgdo8VK6rA0LQXwTjNl0+V6akoHtbLeeKWKybLvQFdC2xtQCFBi5aC2SaqFaCrLSUKPFYymem4KxAincnsofyfckblNmm/NlpaQYHzIHs2AJPyO5rAERrMeBGPc6RuWq+8jc0VFktTmxSmtRYofyvco+VsUAZQxb021bXOXntCBux5SOYo05aFStgIu95jxWiYelSVDZBMx3yVDiS5XPDMghhtDacS5eHVB2P9cgka00CgPCDDEeHioF5NE4xtY3zH0uNTSZbn4ns9oCWPb+WYBMiuTi82gACcMsoOQwn382dopptJGNZDGd3gjqFaXPEa8BXyK/S4lQid1UspE5nTW6tmoQ9rngftmIyKYNXjM2TTDfZK7K6055I8YbfJHxy2dKuv4l59cmLpGXdCugwlqHTENWmkuAGzUhFyUOMiPJysznTGMVPQVVvszpicFjssfoZOXascpYjDEZYzHGkF/4qzJQ8d73ZWQfliXC42IjppVQ4vVg3ULlk9SwWpke2oAh8soy1SqTSMcW62hFOW9hyItsFkEYZSzw3MQfhdea+za1Q8YrFshMraRkH4yNBBQThgQZDipztrC0ACphiOQv/TNkHPglJxM5c/H9Kkg+J+OYDCqvjGYjdVcGKSxQwbGq56jPv6xA0oD0WvGowCiOfvN5nFpcT6kItt2Gd7+pE3ECFb9hGBVHYvhREkydb/8QvvuH71Sw4YGP4aGd/7UEVLz/V/8E8+/+BP7iV/YivjyAhx5fwt1v34t4ehQPffIBfHj2nfjuH24MVMyfO4qvPTe6xoQbSE304VtffwynNmF4cDBsDFbQR+NTeMt/NhJUG61+/8bes0CFTEKljn0bdm0QQrBwaN7eNNBeFfwoBa0Uijn/ZqO5Nbthh9f6l1McavXfOdGUCRdr/lZiNVjpJwk/TFy4AVDBzFGn5PIhmI+tO+9V3U6OI7aACN9ydPXIJ0q7XIUyrNqX0vaum8aYTZXBDidQ4egfWX0ZnWyYVdtf9QfH+RvauOi+muPZyEzbSD8JoyJPRoUDqEilkGAhwwFUHLrvjabrn8bN1OhnscElRd7pyQmDPpPGpoVumYQdnS58j92g9HOorauTIs7M7IwU27kYUHqnrrZWFo6piQlJ+pMrydVABbWtq2sQraARdbWY+nIflLmhaSb/zYIkuw4ta0QYFWICpTQ/1e4mo4KFZo8U2aOxqHRrKuLPTuesdJ3z/FgIsl1e9sZwgaMeNTsIWThOLa9gYZEgAbfPLkf1iaCpNY2C49VVyKZyuNo/wBI9tu/YhcrqajS1NANBD6KxCpV6MvqSAlT4uSgS9Mgj7A8KgMNhmcykpYNZtRW1OMkiB4MoFjQtBZbF2nRyGflMCpd7LyDgIcMyj9MnTyKbTKGrqQHbW5sQM0AFHyECVdw2uycYGFErnwGg6CuKdwi9OTII+EMSmPg9ftRW1aAiEpXjJWCSzmbFS0MLulHZDrut+SOFVMpfuA1oRJYGixg0N/X5MbO8gv/73e9hMZ3Fm3727WKgTgCEAR4Bj1i0QsbexMSk3ENun8XoYiELVyGL6alxYVQ0N9Xjhz94FpGoAhWUfspKp10ekZgCTwz+eH95zfjD4gmfAbJBWHC3QMX05CS+8qUv4bd/+79h9+7djEhK0k+81raAI0DFgspICUDn8+Hxxx+T+Xnf/v3wkVExNaWal9mMgBQri4s6uRhGBYGKRx97FHfecSc6OjpkG8EAA68Cjh49isbGJvFwSKUycv6XL11CyO/HfffdW5J+YrDGe0Y/DEooXbl6GaMjI7jtlpvR1taKaCQkHTtXLvUjXB3HQmIJ/ecu4N7b7pRCat7tQjgQxXImhZn5WfT3nsf+7TvQ3tKMrCsPhtzcx7PPWqCiSbvMpDDvxYsnnkdDfQQtTU3wICzST5OzUxgfG8I+kX7Sbrbnj72IG/bvl+t99syr2NrRimIhj7a2Dnj8fvGoqG1sxUPfeQR/8j/+pJSkWFaFBbDJqLj3nrtw//33i1fOtq1b1duBSQ1BwxylY4IlXV52J0kxOBISk3mRHhODuax0Di0szIuMGrvBKWNXXV0tx6ym2B6R8YlWUtpoGlcvX8Hhw0dkjhAjYCYjYgbNrh0GszSJI9MlK88L2T8CVFRVSTLAAFi7N6lDoIEuPysSUoWiHMep06dw+tVXxZyXsk9kz9AwnAAwped4XNVV9WpoaKQMeBzKrnHj8b//G5w9/xL27NuB5uYuwBVFW3snTp46gaX5SQwMXMPSUk5YaJWxEDyuJO675xa0tnfgQu8AXj5+BonUCvbcsAs37D2I2dkULva/iq4tjWhr24aqeB3SuTR8gTBchTCmJmYxPjqEG27YK/svII/RkWFcvNgr8j4tzS2IxSoxcm0Mp06dQltbM86eO42p8RG8/nU7MZ8s4OgzJ6Tw3VpfiQOH96N9Rw8uXlxCNu1CNOxFLrOIR7/3DdTXxHDkyAFU1HcgkY3CH2xAwRXEPBkVAlRUY3ZsAsdf+C66tvhx44HtuHRhEC8+dxrXJq4ik0ugsaEF7R0taGyqExmlUCgGjyuGixcv48Spl5FMZVDb0Ipde27Ejp4b4PGGMTg0An8oIPeaDy+fN8r5EKgQ6RzxNGG3F72TkionsAlQMTQ0JEAFATL7IuhsgQrLCFCtaI/MzywK27WK0gOcu1zFHBYXFqXjl3EQARTrLbCwkpCEV9cYnfecQAX3y21yDnNKP5HRQC+Kmro4KqJVKGR9WFpM4Nvf/ir6L72Kxflp5DJZpFZWUMjyGcrJWiVrJ+du4/+iIZWR6JCwRaUWCERwTSCqwUdAEu1gQNayLVu7cfjwzahvaBKQhLR9Ne6mXKOyUzg/cr5lIYnrIwsItjhjgQqeM58RrumMN8gs8VJygoiBeVmggs8UiwP8rzIqvLh2bUKS4mAwIICyaJe7iuL1Q6CCMQqBCp7H8PCwJMKc/1dSy1hZC1SQGeHjDxmUEfDeT05OIBKOCPjJ7zFmI6tNDVI5i/C6QbSc2UyQzRUE5BTTUsY2OaOTzDnY1o7yRQEqWCCoqIgKOL4WqOCpq1wfmzoUqBgaHpa5kGbaFqggw4tjxRYPrwdUxHgewYAAD2R2TU1OOIAKFuMgv9MHyEo//asFKlQ/YsPM8cfLocxXZRubFHE3y8k2bqMvF2jXHtXGSlEm39hk32v2YX+1z8+6c3S+4bgum2ECGwIVtsC8KqcqXwRnOb2cS5U75teeNrlZa1+bXLrSx7SL3VTOTWHRFvJKqa1ZkwV0MJ4BBJXJhItGVbZR1tpVZWE9KaeUUzm/u455tAEXnbmjlH5NDuXe4AJvYu+wrtCtJ23H3+oNrbq/Nld23lfzb1ugtHO4vZDO49Uxs/n2BSCwrAqZbxSMcII6cl9sQ6KR2XFWD8omyhZU0b+K9BHBV9OoYYt/UtQ3bBUrOcTOaauAIPJ3JU1+IyVqGgXWSoBZBQYWo5UQY7woDMNO5lDTJc1jYnwsflTsIhd/CZWAkcK5yTGlq92Axvy3ldYpXVczGKW4aQrjthNePIes54GseVooFUNkO3ZMIV1kZ8y+5N9k9hoJJwFPBEHSrm8FdZRhFyALTzwvyBhQkMMCEvwcj1PYdQRjJA7S68LPSwOOKdbzfAlAsllImiMpHUSWBTvRjdyW04eDx28BFVt/4vboF2G9OuQam9yXx8BczRyAVoCMLwCPZxXbxHhlMlYQtrU5D+cY57/5N8b0vE6Uu6aHphT+i0XDAFVlCZXbUo8oK7HEeyyNETQp5+elmJ4yTRmUJiUIlJfGCwJE0tnv9wuT2s1cN09Fg6DcX7kvIkWl4AbjHGtezfvIRk82P0kMZc6bc1sqmS7tTxkaOh61JlKW5NSivD6HLMbxmaAKAxkKyi6hX4rWUlQiSfdl/2uBOisVxriP1+pzf1ael3/5vWzSUfCEABhBCokn3Nq4sby8AspBKpijgIGWrRS407HP/bMBstywnEwnBUizOY/mhUUF1wxbRO6PeE4oI8o5TnW60hoaAQpljGj8KHJsBQUVnP6m6m2jjCMeokhJlZqotXnFSmpZ82/LIrGMEsvi4b5tYyxrIK8NRkV6AF/80Afx/odG16zbfty9yqPiDzH+HxzeE7/2cfzZy2tlmLiJGrz9d34ff/H+vYjPnsBnfv1TOPlTv18GKt73AL7meSv+4vMfwru7VWeOL4If7/nPX8TVuz66KVDxowCSdZHHmjdWgxWvPZCCl+PTb+w2V8WEg9IZagMwGzOoGbYGAJYSa0r5a4r1dkGwi6QWZsu7ELqVCXpK1MxV5AJNjEtBjONfztjULmYyMdo6+6ra/3UK/URR1wWmthBf3nM5gNIuOdvZIJp4DnqnTULkVOU6leNO7WxQox65dDaAE8CnrGNqAxjRFzQ+BhKQCEq6/lxsE44tfEuBjxOy6TxU2Gnt90pE19I90eKW5lEazxj9RNsjZPat114/ZMNITUrLHhUq/URDbQUqxDzRAhXm32RYHLz3TdrxJ932STU4KxYxPT2FhdkZ0R3m4sMFXBb4ZYIBaaVFUoqFgYnpMGKCLMVEyqCw07u1VQoNLCLOiSFoFCPD16Tru8EwKsBgLpcXY2RKByRSSekwaGxoQDRGKQGaPCtdkGu87TCwQIV0wnBBL6iZ9lqgIidm2kpN5N9E+qnIxFq7YyXoMeOAAROT+u6uLVqcX0lhYXFRgjsBKjIsSCZF+mBo6Co6ujoxP7OAK5euiP7ijp5diFXG0dLeCm/ED790MFYIGFBiVPgDUjhnoEUPiaBZ4BMry8K0YLGFJuA8bxZrNPgsGNAlh9RKAguz05iZHMXC1AR2bt2C5YUFXDjfi/ExFgFrsWdrJyJ+anS7pAOWndGzC4sSDFXG44hGKwUc4P1ggR1FrhUFLC8tY2ZyGtlkFnU1tWhhMSlIVgY7PlOYmVvE7NwsFpeW5ZgqqqpEg50/FfE4YpVVUtyjDrk8e+xEEKAiiYceeQypogv3vflnkBfPCzWfYmDHY+G4GhsbVzpsrFIYIMV8FoVsCuOjwxi40i/Fz2fXABUMpQlURCuickzs4iBYxmCBXfMsSHNckGrLvMrJqPjql/83Pv7xj2HP3j1SKON14jMgJsuG+s0xPb+wKF0lFqh47LFH5Xm+Yd8+BKNRYYLwOlI7f3FuVgp80swH7cy46RYyKp7AnXfcgfb2dgkOKf1UyGdEaonSKCwkklHB8z/36hnEY7H1QEUkIowfmlIPDA5gbPQaDuzbh3icfioe1NfWYX5uBt6QH+FYFKMDw2iMV8tYzrldCPkiWM6kMUeGSm8v9m/bjtbmRgEqWG3inEEz7D179orGvCRILOwF/HjpxDE0NkTR1twsZtr5ohtTs1MYGRnAgT17SonQcy8cw779B6RAdv7cWXS2KlDR3tYBbyCIsxf7UdfUjm9/92F89sE/VuBPgnwW6Lg/nScjIQ/uved1AlQsLyVE+onFUyZC/GHx1BZo+fyzIMtXOER5F4IFWSwuLogECzumCU40NDQCbkrIkR7sRyQaEcNbBtrjE5MIx2rFD+bqlSs4dOhGkTsRZgSdLYSCrvRiAnz8XfxwpOuJgHBKfG04l0jAK2urGttx/uK45NiiMfWlS/1SVNm2YzsamhrkGd+6ZavcRxZkpiYm5bmoqa6V7ilJlsnOMDTr0ydP4Ngz30ZjU1QK/rm8H0ND02DuXHRlURHzor//CmprW3H16hBGR4ewpb0WRw7vQTgaRayiHi8eO4XB4VHs3kug4jD83hq8cvJF+PxFBIIxeQaCYT8amlsQClZhdmoRVy/3iqm3FNxFacCFRGIRF/t64XFRfi2Eq4OXpRhaU9OIyYl5/M1Xv4IDuyK47a77sLgCvPjcC8gk57F911bs3H8ALx67JEyIjvZmVFYGceyFZxDyu3HzzYfRtW0fkrkwZhfYghUUgI3yOrFQNWbGx/DKS3+PLVvC2NLVgu98+weYnc7A7XOhpjaOleUUZmZGUFMbRmdni0ijhYMVgMuLwdERRGNxdG/bi1C4FgWQjeXB0NAoPEGXYTmoRwWBChacObdEIkG5/5yrSE0vAxWU0KMcj2VUjAkgv6NnRwmo4P1jssdrRtaFBSpkTLlpCr0kILWVcOK4rK6Jo5BNCw2fMogETyxQwfG1lExIAZz3iuCFSqCR7bEs3ggcd1b6iYxHzmlkH0zPzMLtc6MyHkVlpArTE4s49vwxPP/ck/D60pgaH0aayTIlBgg2MAGnKTyTTq9fChTWhHNVIcbDzlQCDerlw7HL7jSl3mu3INlzO3ftxo03HkFtXYMk65mMyl8JUEHj+mBAQGZZ9wiW28K76agk0Mdnn0USC1QQKCerYi1QYRPnkBhTqkwTj3F0ZEpAd66BBG3EDDFPMD4NduWlHEAFi5m8T2y2IKOCP5ZRYaWfwsIA5TlEpEubQAW9TRSoUKaHAhWcQyiOqEk2v88ojsU3NkrynDkPynMvnddsj1QtcV7HqakxYXMpoyKgfdVkjpnYj+OrzKhgMQIYuuYEKvR4uJ5zDP84QEWUpvKUuWJxJpXG5MRqoIKm2uFIUMaoTdgFqCBDxqcm5gS7rZ8Yz8PZm+Msjq76gzNH3ARc+FF55T/J3zfc92achuvtcRNwYRNDa3oJbpY5/UMZFZsdVbnVzZSkf6zrrJI8q17XQTbWwg72nKSovGHBfv2b1wMqbP7B+EUyLeNPIJJ0JYaF7fzXpJkNDN5AANcGBqQZSoBgk8itGo8m1bLgyboszhb+1xyyE2yx2+N3JdcwjV5r70lxQ5a9MqM2fq0GEuyxlQCGja6tOV7bgVwCsBzGyDY3ltx3kwsvTDmHsTG/IxJBlCAyMsR8TwGH1X4Sax9rzgWWSSi5uSn0C3jq8JgoFZ7XoTxG9MWcA9dlAqaM0ZQRvNn1MzUAUyixTxvvHb9jDZuls9to6ysoYRg5ZhKzcjFyvYw0jfVd0zFojHxtCackRWMkfBgz0q/AzN0i+2MKuLZ4LNfUSCZxf4wVOB9zfeHab0ERYaiw4G9YIWXgSO8FQXFhmBuARdYLnpuA5KZznUVw0yXOvwtbQgraKi/E85Q1ij5LBqiwzJMSK5qgCHMiA4ow37VAA+8v121uy9YMdKwpSGJZMTxOu/3SeRlGhhyXUVaQ+oW5xsL4oIOdsA50jbV+JczDKWmooJPWLXge+nzq0yNgotTcNOa3bBcpdotsOce3ghj8sNPvguPCjnWCAbw3ySTlOX0CknCbAnwIqMU8Qr0gFAShBCTBAub7vA/lWp0W8vWpsVJIjH3I7LBMGMk12NXvkCuznxeJyCybltiIQVDLj1RGJa+knmUYQvy88/pbdo4FLr7gkH5636+oKoTISwrgYTxMhMmTNSCeyjRZsE/nHFW2sI9kaY6WW2C8Sgy4yTyejYz8rHxHwB8FLHj92CylTTNktlOZg8CNXlPWgwS8M2oaKv1EcE3vd3msKUtdgQk9LJUZ05WRQ4O1M61D6b2iSoacowPE0zlMZdiZD3JcyHh/TUg//dhAxQfxyLaP4hu/91b0RJZw7HO/i3d98ijG16xuwYPvxJc/+xt4e5ffgA/fRPy//OkqoOKLvX7c/YHfx5c/dCsa2ZgzewYP/ubH8eFHRtH59n8+oIKHqmDFIcx/97XFpLC36XffaD0qjGabY4G1PgT6cPDHFNtLlCRHwV4jjdKDZhdgnevM02g6CEpEVRtw2enaVPhLxXw7i1vi7pq1vwQWiOdEeeBtFmqvDh7WBhJm0TBAyurAUZcSOS4bYJgAZRVgYQ/BMCokyDHnL4uN5M929nc8KA62gg3YhMJlwBGrXbnq0TJGSaVLZxY+XXyt14STRWLuQ+kYzT8cF84CFabiaWZQs1jZ723GqDCG1+yzdZAlAAAgAElEQVSC5w8BCbIo+F9hVFigIpXCwZ/6aQNU0IgzVZJXoXRBJplCdVWlLM4snHGRYFC0ML9gzHznRUqKp6uUPzXW4rViEm2NJLng0AC4qaERp0+/KmaM7CKn9JObtLt8DrUNjVKkX5HO5LiyMMSMWqWTCFQwvVePCtWi1EBC5YZcRbcUpBmMsDCp0k/0OiBbQLtf+Dcm6Pwuiwg2WOfCwmCNhUT6DfTs2CELOiWgFkxASLNPFqJXlpfETHt6ekLOgd08589eQCgQxvYdPYjEKtDc2owaav+7tPOCBSYNMgPaiZHJIJNOiY46AyzpiPH7EQyHBM3n8bHTkkWeqclJ6aglGED5hnRyCVMTo0jMTMGdWoGf3SzpJJaTKQxfG0VdPI4dXe0I+zzaheMqYiWZwhIlc4RSTNM1Bk0uYVbQfJjKJVXxmHgYLM0vYHp0AvW19di+dSsqSIl3ucFOh4nxaSRWElJQ5z1lAsqAiYASNdQ7OregprZWC2quIgoMgrw+TMwt4qGHH0NVUyv2HDoMN3donhkWjJkkchwRaCFYEIvShJ3FaLJXVjA8cAUjI8PoaGvFD3/wDCriNfi5d/w7dHZ1i68HPSpoAE8QitIUwkopFAXoqamtkS5QFko4PsnMoaQZ2T1f/+pX8Vsf+Qhu2HcDipR+IsjhBCroz+Hxigb64uKSUE5ZdHnsscdkvOy94QaEYlFMTE7CL3JAaSzMziKbTmnwj6IADzfddDO+f/QpYVTQq0GKcX4XlhNzeOmlY9i6ZTuqa+plfM/Nz+Ll4y+iub4B95JRQRaLMdQWRgUL8p4ABgauYmlxEXfecbsEwyxI8l5SWicYDUsgRXZHTLqW/QIahYIxJHN5zCzO4XJfH/Zt60ZTQx3yrrxIyOTyRTx/7Dh27dyFmopoSTLLF47glVMvo6WxSqSi3PAjnS9idmEe14YHcOPe3RqQFl049tJx7DtwQPT+z509i86OdmYFaKeZtseL8xevoKqxFX/38OP47P/878ICIgDIJEkKocZokh4M9913N977y7+M5cQyttKPREAKXg+VfxI2g9GWJZBEA1sCQNlsQhIVJjkcjzU1tcog8gXhC7Dr11/SsVfZuDxS6QzyRRpHz+PK5Ss4sP8GBencmqwzKeeYEmM5obFrp4+ed167tUJkaSkAJ0BXUen3Y2OjAlBMTE4I6Ml59MiRw2hubcXc4pJ0YNMsvIrydyhianJKOr2rK+MyJnhdJfAt5sXc+MnHv4eKaAZ79u6gaC3aO3vg81Tg+EsncelSL6pqi5iZW0BtbTPqa2tx+pUXUV8bRUNjDS71X8Vtt92F8fEZXLx0Bbv27MfOnhsRDjfi5RMvIRT2yHPFazkxNSaMqaaGDhn3IyNXQQ+QlpZW9SkoqrH44vwCXnnpGWRyS6hrrEQ4yq41DybGl/Dcsy9iuP8Z3H7XHTh46CaMDg/j3Kun0NLRiD03HsC5V0fw9NMvSAJRV1MFD3IIh7w4cGg/Gpu7EI41ILFSxPxSDjPzCZFiCodiGB++jNOvPIGenfVobKjHY4+8iEi4CV3dWxCJBjEzNY1XXnkR83OjCIbcqK2Nq8FzXR3C0TDCkQqEwlUIBGkIHkc250d//xC8EQ/yUpxR83QWsmmaTKCa8yWTSWr3E6woARV8vqAyRQS2KU00PDiMHTt7lLnDhJlAhWFUcF5ioZ3rpowhjw+LiSX5rnRjFYsiCVhdUyXPBmUAad5ckn6SNdeNpdSKPC8cd2SkWaCCzwtBAcZYZBLxmOlRwTmJUgdTM3NiLB+NsfgcwamXzuKhbz6ElZVppNMzyOXI6ssJS5B6RMV8AV4X5YuALKnwpmtOPGCMISTXfEoBMlFkpyePj4bQLMCIrjiZTWQ6hsPY2r1dwMyenXtE0iqd5UrCIn9Q5RH9fnkOCSBWxKLwiYyUkQIpFDA+Pq5AWigoTQ7TM9MlBp9T+sknsgNqHhmkFKEFKtw+jI1NS6xTGY/JteC9YKzA5guuIZxTCeoT2OD+mCgLIERGRXoFlZVx8YAie5PFed57siA87oCYaU9NTyEajkrHKKWWJBU25o+MYFnPY2GBTAyRsyxmZS3jvGXZFLavqJin+a5qLU9Nj0scUxELq8eU4BfGpJTmpJbdWJJ+Ksr8ws9Y6SdqX7NQIUaV4vGk91TnNWpXU/opIHKMXFeiobDEc5TryKRSwggLhQgqqVQCfyLRkNzLEqNiivOv3s9/EFCxJmf9l/t182LmZgyMfwxUsdH5lOVWVv/1ekDFRsekMuarz8NZvN4Q9Ch/wGaHP+KS6/bXbksNsjfwjzDH5DyqVce00WXflHli9r0297QSKPmCSKawaMYmIXamlBrapBBmG8G0mOQNBjF0+bIwIdksY9lOIp/iOENtQFt/txV4MDCM45hKgMRmbPzNgIpSjrr6FqzKwUt/ssyg8o7L92SDvNYCLqaYbot12nVt8kqbD5dAC+YLGz8XUgxkl7KVczLFa45BstZKghCGpaCMlA1eBoy14IptCBT2oLl/tpFOpJ+MlO2qLUl9U8/eGglbk1t+RzTzN9q1g6VgwS79nN5TLchTXtgnNVSOD9ssok2FppFRGq8UTLYNdDwc618ghWbTCGnZJZwTBeQ3Ej5SyDdeEsKot14J5qbaRjuRYMrlpMnm1Csn0dzSIvky41MBwU0Tq5yFo8lStq2FI1lXecVKjBRTS9HGyrKUF4+ReTevIYvd1shZO+EVsLBAilwP3msC7cJCYc9AeU3h59UfUtmL7DaXYxS/D42reT2cXhYWwNLai20aVekdBU+0EE0WJo/Fgh8CROaMzwbNukVSMS/rF6WcGYPzTWV4qCwVc0Ruh7GH+Fz6LMjCTnsel9Msulw7sk2tMl6M/yrvnTBMAtxWRpoURFrImKyzzsIcmWul4pbq5aESY1QmIONCGz6VDaDHz1yUY5n5tx5nWuWKvLo/OU5ugwbx4h2ijaNSvBcWg8pA265/GbNklZtGVQUDrEy1shBEmsrI7X7pS1qL4YvSTzx35joqPapy3IwJeZwcW0uJJQFmePyMH6SGU6TsE/MvMiy0nsNGINYTJI4pZoWlLDKbKysqZ2XYMDpmVVrNzFjCpOV+KdPFbch1Eha8MjdE/ozHQ+YFAY2APnfi2ykG48qgsWCLlUdj7UrkVAvqEclcQMaryHCpV6v+bozATSwvzAs2mNua5E+Aigfx5Q8fQiOln+7/IB4c3ouPPPgJfOL1zQBlm/70j/GBB58vgRXB3W/AH3z6N/BrR2qAxT782QMP4AMPLeHtn1oLVABouhWf+OzHxJy79+t/iHd98DugxcQ/N1Cx0Tr2Wnrvk68nUCGt9GCQCtM5wMBJbfF01ZLJhn/Xmr28JNlwBjoWqDCo36qF2lHgl4BAqvZmRVxj17BReFZic5ibI4dhbBTKwfIaiKK0eWUvaCRg/m9V1Fv+RbtS7XZUj1LPVQ2V9BeDvVja74YDRpFwBSuMlJMFKhxo+tqvyqZLrAhTVBBXq/Uhv4GFFJ23AbFFUsyBOr+ll9sZZErIopel1NljT9CcpGWOlA7UXEnjT1E202a3r4IUIv3EAjvBCQdQIR4VqRT23ftGSXi5h6QUX7JILC1hcmJSEkwWCngfuDCGw9SWzkoheGF+RvTeuTjYwgWLvOXOGKUAskjKcckFix0WE+Pj0tXOopF4VLh9IM5dWVMLb5DdmrqQMullB6oFFAQBZ/CQL8gxyqIoVG1j4JxX5FuMmoKU1gkYjwoWNWlixUUrJ0AFF5NoWJkiyrZgMOoRWR0uTux65/Z5nOymp+SBGImmU0guJ6STnV4VxTwEgDl37rwsrlu7u6WAUVtTh5rWZkRiMel6sLRcFk4ZrLDAvLK8LIsnix9cFGXxM+ZkTAK8LAB4vVI0YQFfu0NcSCwvILm8iAAprlMzGLnYB6/XJZ4YLOQFfX60NTUhSJNVCbAL0iE6sbKCmbl5kTdi0ELpEz5CHe1taG2qweLsNCKhAEJevxTaO9vbsXP7dlTVNYB1JPofsPii9GePdDBQQz8QUmkLamszQGFBLBSMCEiTY23F7cfQ6CT+z7f/HofvfB1qWjvgZRLpVmkLBgkEOcg8YOeqMCpCMZFFyuYowbGIK1cuYWJ8UpguR598AlV1jXjb296Fjq6tqlvrZbDlUcqs6b5YXEgIUFFXV6+GaCLtAaXu5vOYGB3D//363+DDv/kh7L9xP4oejwRGHM/qj6ITIY9vZnZOCoEMLBm4PfH44xIwstgWrohgbGIcDI3y2QzmZ2aQSa7A56e6vFsKmoeP3ITvf//7wpBQ7wd2lxZw7dpFXO7vxc7tu+D1s2gawdzSDF5+6Xl0NLfgnnvukWIfn2WCaHz+EstJFOHDyNiYBFm33367PKcryRXp4o4EvCIZI4AMDdPZWZbNSdE+HK1E3ufFPOWl+i7ixp4eNNZVoeAiFZxdWB6cPHMRW9rbURX2CABW8HjhjVTg1bNn0dbUgLrKSjn3VK6AueVljI+O4Iad26VwzYL6qVfPYtfuvfD6Azh1+jRa21pQTKfQ1dwo092V4TFEaurx948fxR/80e8hn1gCVpLIFNI6Xkh3z7sQDHnw5je9Ab/4C78gz8q27m4FKYRNkRVwgeOOOrcMwEfHxvDyyyewtasJ3d3NUtB2gSZ2HtRUN6C6tkEKwpRCsh1KFlS102m+4BI/gKtXBrB7905hotBcmGNRp2oFYZUtp901WkC1FHkawalfDsfc2NgkhoYHMTZBTX0fOjra0dLSjLHxa+ju3gqvL4i5+WUx6+XfmHDypiV4TTgnxkIogF1SPikYz0xeww+e+h6SS9Po2b1VGBSRSDWqa1rQ0b4dy4kUHn7kYYxNnUaoIoLa2kZkluYxNzaA7u2dKPh8OPbcy2hubEYwHJC5tGfnQezZczMCwRqcPHkShWIS+/btk/FC+b+JiXFdO1FEKqPmf52dW+D1sJs7gMWFZYyOTGJi+AIWFicQq/Shuo5FdQ/On7ks5zc1MYalxWu4565D6O5sx5nTZ4WCvf/QPkxOFfDwE88gGI1gfmoS/kIOLS11OHjrAaSzLOL70d3dg4WFIkbGkkimC5hfmMXY8DnMTvbhppv3oaOjC4ODc8hlQ5iem8PI6BDmZ2cFEGpuahYmxOj4NfHqCIf8aG2Io7auBpFYpYAVkUgd/P5qDA1NAuEA0sxBPJyr/eqtFPRLoT0ciYp2P+cVelQIKO7VQiwb9/h8EtCcnJzCwOAwenbtRFVVtURv9NohO5HrLKWKCESZEQW32ydSbQT+uBa6KHkUior0YS6fEQBVOv8NhZ1zJDeUSKVLQEVyRYsAXC84V9GXhZ8he4PrHBkV4v2wsICZqVm5p7F4GLRLOnHsNEYGrmF2ehiX+l8WwMLGVSyQy4+cBVDw2qBTixoEYLh28pkIRWISsorWc45+O0lhdEoXsTwjBYkH6hubsGPnLpkX29o7kCtwdHkR8EVEPonHu7xCqcKkAC5elzGcpmSiASqE7UJwmqDz9FRJAtLZ1OLzaIcmfzhXyLxrGBXjwwQqUqiqroDPrwk8QYpcriCgJddJ9ahwiRwc51qCDslkAivJZZG0FOadR+WjeO+5BmYzBUyMTWFubkHil0CI0ons+MyL3400WVhjVQOiqFxqGWxQ+SdHF2WOZQ0FaqZnJrRQRYk7AmQe1QGXrkcOW6dnlOn+HRockqItv0MQ0eNXn5zksspgCshkgArOaYxL6CfE+0fAiJJn7PClsTmv0eQEgaKgASl4jd0IhUMCxIn2NKXyyKj4FwAqNi7ibpgEXPdNE3lvkj1s9LZAT5tsc0NIYNPPb3YOmwIVm7AeNgIqSinSpkyJ6wA0G572xkCISVzWfUOv0vp92FlkQ0ziHwhU2KIjnwfmLozRApGwNBapebFN2cpzl1wXnxcXL1wQ/x7G7WX/Ei2Gai5ml/6Nz+G6QIVBGktFK7M9e0+cF2tj+Mcew0b3SAu8a8fgqpG35ms23bZvW1acZXnY90tXqcjYZ/XL/i5FccP6FxaFLewLMKAxFucl+1rdbFjeJiW45HqIn5EqCHDcc8xIEdBIHWnMpjdynQKDYR7x77Z7W+SLHIbSG41BGweulYTiNbVSOnJeAsCZQrkpTlqfibJ0ldZg+JLiu8kdtPHAphPaqS9xY8nkWOde+YhRJrDNCiJ5Y/zypODMfI4Ci9kcqmtr8Nwzz6C1rQ0VlXEjA1VwFOhtEVzjVAcGpU0ExstD/2aBhzJIoQVZn+RD9lra4nKpaZM+C+m05IK8L+oHYAvrOZEo1DVTPbN43OpxoYwMGz+LDwAZ3dKEpHJGZTNz7U4XqR7TBCHm5JRSCoVKkpfchi2EU6pZ2AniY6BghBbdaZ6dLDUssImCOZ1lVdgiNIEEqhrws0QNLABij1difhv/W2kzMgsEKCqbsFu/Eeb1wr4g40EYCCqHZK+DxI8EF6T5yYJNOk6skTWPXdUudI23voVcY/kdbdhiw4VKD/G7BFt4Te3zpc+pPt0iT2a8Rax6gAVLFNzTfVjWB5/LL36x7FHxy+/VAr9tFlWJJfWC4H4Yo0ZiEXmGCQIxXuB/ea52Pyqhq7Ucjn9RuKVccka9MziPM7akLK8+o+r7Z03LdT6wwIoCEBwrPG+JiVgrEh9Tn9RTBFxl3cGYntv5QRpYCKSJv4qOE5EjlVqssm8sY0QlrNS3Ra9lWUuf11+k2mRsmNrhT4CKNUDFaYCMib/4o/+Ed/fQ/C+D8f6rGJjNAB4/GrftQCfZ47kZHP3cp/CezxDEiG0MVGwSfl0PqEiN9eHU8EZyU2kkJ/rwxf/xeXytd6O/b7Kz1+Dbv33fVnPWuuDZYEn10ZTGpsguOUY2iDE6jA4kfe2lsxJPNhiyD7iTgVAKJGTXZZBhFYW1HHZoYGIW11Iwsi4oXR+w22BEA5vSVja426aL1LFPG9CrqoahU5rOhrLM0vpuH9vpL912Qtnj5KITtgILVgLLGUmWJabszVhl1GZPrQQelKIRxxGrfqV+X/dhv6aBk5nszDa0k8cJVFga8+qIs3Tdr8eoyFmggowKyj6l5b8JSkOkDKsinUbXkdsEEedPNpUWtHp+bh7TU1OojFVIMu5MgtlhR/+JbDYlpsQsPPAzDPYptcMffkYon0zEvV7xWpBgjIn29DSy6bQUTtpb2+DyEKgoIlZdIzrWLKDpAuUT41pN2JUaGQ5rAUy0PIU+yUVbuza4bQYWDKw2AyosE4CBTiyiBVcWEAqFrHRTkE3B/TQ3t8g5s0BKoIKB2ML8HJbmZ0Xblt4JNOkuZFWbkx2UPM7t23egsrJKrkWwsgL1jY0lk1P7fEnRmdJAHo9KJkmnLLtcuE01YZMFl4abPu1ooQEqryf17LPpZaCYQyifx3TfRSTGxhGPR8UTI1Nwyz1sa2kWQ9RIMCSd/vQ+GJ2fE6CCIIVLdF4J9gFV1VWojUdETorn5me0kM+je8sW7Nm5ExU1dUims1IIHhweksJXOkutUg/q6hvQ0tQixXfq09tO8nhlNdx+DzLcVNGDc31X8OQPX8Bdb/ppBOPVKNL8isUZua8+KXDwvrFzlUW5WCgm7JFMllrwcyItw2uwc3sPvv/4Y6gUoOIdwuAQgMTH56SoGuomKJ2ZnpOCYn19oxpzma4qC1SMj4zi/3ztq/itBz6CfQf2EZEoARXa7axPqgAVc/MCztmi1xOPPyEBFD0qCFRMzUyLxga7nwlUpFeWhX0Bt1eAikOHD+Po0e/jLW95q7BH+F23O4feCyexMD+FrvatyOUDYkicLaRw8pXj2NragbvuvEu6nxjgUc6FWvssQhbdOlY5Vu64444SvVbuTWpZgDApboYjYvAspqlwoTJehbzPw5YWXDzfi4M9PaivrULRw+7pAnJFL85eGEBHawuqQ+yYzyBL5l4ghAu9F9HSUI8ajleGES4X5peXMTk+hp6tXRKg54sunD3fi+5t2wWoOH3mDBqam1FIpdDZ1CDFtpHxGURq43j4yRfw6c/8DrIL8yiurCBbSCNDMXZ26edRAip+6Zd+CYvz89i+bbvMTdLlklf5J847FihlF/u1a8Oor60QKSANLFlADqCquh7xqlqJhEskOpMAO9dAxrG8hpf7B7B7z04Jrl08Jv6YnNsW9koJpwEqpMDnZqCufjkL84s4c6YXuUIGTc31Ij1FSSQ+XlcHKMtUI/JDi4srGB4eEqYNgQoGwGLkViwiFPQJ2EWwZXlxASdeehaDl8+hZ3snquuacObsBezffxiMr3ds3y0SQj985ocYHT+HSEUELW0dePw730TQlcSttx9BwedHf99VjF4bkQJnW0cHdu2mEfdN8HhiGB4eQSabQltbW8m3iM8AAby5uVnMLcwKWKrPux77+Pg0/F4yDhaFdXDy1MvIF7Joam7QoJ0+Iaksnnn6e2ioDWNPz3YsLSxjKbGAGw/vhS9QjwtXRqS7dWRgCMnZOXjceRy89SBGR6dw5sxZ3HHXzeIjMTaWwtM/OIHpuVmgsIBcegy333EYTS1tOPb8eVy+PIFULisSWq1tHdiypVu8KthRNTE5jqsDlzA00I/EwjX4/W40NTehpqYKlRVViITiSGXY7lWDXNGHvItyNQSRK8XfgGtdOOJDMMRu/wUsJ1ZMYm4K4G4y1EJYWlrGxNQUBoeGsaNnJ+IEKli8dymjgsv+7NyMmkZL16R2Ni4kFjHDZ4HvFMpABU0SOfdYdiLHGe8Hx+EyO9QMoyKVzMi2mWQrUEFGRUHGM+fqMlAxj6mpOYl94rUV0r0/fHUChVQGjz7yt+jrPY5cjtrQJp4xQEWpicLDhNEUybj+Ut1POuu9qIhFxFuHIEs+k8dyMikADFmc6sXBbN0NXyCI+qYm7D9wI47cfLM8B3D5SkAF95VMryCbSckzY4EKq4XNjn4CNwQqeL8tUGGL9DYAI1Bhk1ACb6uAiqEpec4IVHh96mfD9Zc1hFRGgYrKykpZN8hwYsMBmTgrywmkMoZRwWK9V7Wo6f/A+C2ZzGB8bArz80uoiFYgEPYhEOC8ALgLZbkKHiOPTRiXDEsFqGABxvpUOIxwCVSIKXkBM7OTsiZwbpLOUOYDIoVgonur420YfdzeNQIVZOlEgnIOHq7NuRySCTXT1uKCFjm0a5nyW2FhOXINZRzBAhQloJi0s9lEgQotSnh96ufC8W2LWtlpMipC/+yMin8qoEJygQ2ykM3L+P8SQMV6hsL10mIFKlZ3rv8obwdZrJzJpnMHG5z8ZqDDuoK5zU//EUDFeilgU16zx7PuuIraLRsMILGocRqB75w0UXGO1bmsDD4Y2RafVyQw6xsahC1XZqk45YQVaFlnUm6ukzVKXjt2ZFxaSpS9po58d+190ca1jfgLm3mq2PmhfDE2AxVKu9fEsWROLCCOKayzAOicQ/TfyppY+7JAhqnGmeGjDRzM5UTuyUrRmQZBk9iu25YyXpSZqsVba3SuqhGUr7Wd3iXAx+FDpNvVeoUTqLDzqxZBN+E+mQK+1AekDqD5v5gfi+4+WXgqiepze03RUoEHkRSSj+vzI14PfF86+MuAyWpJbePXYZosLcNBWPWGhcB5ngVVBdjITDBFUcpPSeNaUkF3nw8vnziBrVu3akONBToMK46/c+xbfX1nb6UMTcNOsfUGYdOJd4EWXxlnMxe20j6aC3F7RrrMNGzaIj6vM79DQJvXi2sTQW3uh8ctDYHi+eCVcaLyU2pGTtYKX2r4rZJQ/BvzNvHEMOCOaP7TBNl0+AvrwXhs2C59xbKUgSH+blIf0H1QtpC1CGUbUFmAMZOaHkuBmp4G4i9XNv+2oA476m3dhV325dqVATON3wM/U/IoYM4pMmjKluD7/JGGRcPwZy0vn+M10iYGkYiW89Q4QJsIeD4qraYSWFauWj0otJ6nBXbL6LFeFNIMSCaGAB1piS84dtSjwsp9qQSW1hi1ZsV7oQwN3T7/+4UvKPjHFxkVHKti9C7sAX2fY1bluoqgnLU0U9A8PRwW8IL3RRsbdcyzPsR4luoZsnYZw22t0akviLIctP5pJcusz4TOy+pZwnsoOZgBKC2rQmMcI0lXVLDMjnuRKDXX1Y43jvsy+0PNsW3d0jLp7ZxlPTZY+5DbIM12hkH1E+mntR4VH8SDp3WgBPe9FX/wkftx/13NKBN19G+psTN46C8/jw9/7oRhWvzTARXrViDnG7Mn8PFffwCfeZqdgj95bXYFPvq6LvnT6oZ9g4CSGiZAhWqtiY5aSXLI0o/KwYY+iFYmyiD9BgHUIGR14KYdDfbIDFDByVKYCo5gaEMGggFWSuwM3Y7dnnNitd1b9vj0cw4D6dLFUfRUEUvdf/n/NUlYWzQqHb3DdEmCBkHjy0i3nbhKgZkjRdFYUhkYvMYql6OLPl+CjjsAGkv9k8nJghbWgMt8x8x05qJYTNuZ6FhgSoM928WjHS/lSbUEcpiu3tIVMYwKTrg8Xho3MVhgx4AyKixQkRYPCEoB2fea9x+SYl9NdY3II7CQS9kMFkeoec+Fz5pUWwkaBizhEKWdVMufkzqTei5EBCK4X7I0+Lf5uTl5X0ALFvxFezovxS4LVOSKBdQ2NiEr1D9qKHql4B+LUCs9ogAEPTIKaoZJ3WqLpDPgYDGBCzs7N3gulH4izbMyXimLnOhRirFxXo6Vx6dABYuxZaCCxXh2UtAUXApCBCoWl4SlsLyyhKmxUSQosVMZRXIlgYpIBa5cuSK631wgd+zokWJwa3MLlgt5tLS2SgJvfRO42LL7kteB++Y1sxRDBl8aqNC8VLX6ef14PvT0YEBAoCLscyOVTMC9soKhk6fgTabQ3NKARDaJHLVO0xm0NjchGgxKoSRqTMOnVxJYTCSkcM4AReJNl1uCIq+ngHAwAK/LjTQNVNNZdHV0YEf3NgGQ6HUyPj2FK0PcsmkAACAASURBVANXcb6vV7t/5+dRGatEZ2s7tm3bhu6t3WhtbZd7TTPVSGUUaQ+QyQHHTpzGmUtXcO/PvBWuUBRZdkuYtIzjhNeA50mvBymwBwlUcOyuIJGYRV/vBTF73dXTgycffRRxA1S0d3QpoZoMK5HfocSXJpnjY5MyFmniLECFKdw4gYqv/81X8LGPfhR7990g4A0LM/ysE6jgfaKZNp8HW/R68gkCFV7sP3AAoVgYc+yEzmSRSSXF1yWdTMoYJluI1+OgASre8Y53yrb5/BDsOn/+ZeQyy2hubEMy5YbHF4I36MbpU6+gu60Ld9x2h4AUlDOg+ZtQlxPLcqwEBPm67bbb5L989pcSCbh9XizMz6Ovt1ck2m656SbTGEI5Nj/maCJXXY3hK1exf/t21FZVoOBh8kWaqxcX+ofR3tyEqpAHPg/tcd3Iun242H8ZTfQjqaxUYzQ+y8mkdNd2t7dob5/Lg4uXLqOjq0s6cl89ex41TU3Ip5LobGyQTrmx6TlEqmN48pmT+N1PfhTp2RkUDFCRIkXJMCpYFH7TG1+P97znPZidnsaO7Tsk6dEOnJyYanPcWAM3Md8ljTjoRzQSFPYV5WTcnoCAFPF4tSYkApBpcilBv2OxpfQVO4gv91/F7t27RHednydYQYk3O+/bhNmuN7ZDSren2vxkb3EsE8jldmzAzxO8NnINoWAYVdU1IiM0MDAghuhV1dWmYKqeHZSvE7mdTBpnT7+Cvt7TaKqPiyzVQsKDl46/jFtuuQXziwnwWaB/wzOURou5cW1kRJhGfWdeQkUgi8NH9iORK2BpcVlAVxoEkwG2c9d+dHfvRTBYhQwL9cYsnJdFOhpl2VQdWMoT9fdfxMrKElpamqQo29TYLKBZrrAijI7JiTk57kIhCY8vjbqGGHx5Hx5+5G8Rj/ogpfkir1EaBw/vRX1TNwYnZhGIxOCHF9cu9mNg4DIO3XIIoyNzeOrJxxCuKOAtP/sz2LplH148dgG9fVfQ2lKLsZE+7N7bDW8ghEcffg5VVW1oaW9HXUMdqmrrEAlXirlxLleUJJVd+mRojQz3ou/Cq1hcnBJfjObGOtTXkVkRRaEYRyAUR5FeJu4wgqEqBALcRgGRMBCNBASM4DzKa8JERRpIXGS3RAQkIFAxNHQN23t0PeC497q94lfERI1jjGNROhHF/NgtQMVGjAr673Du4Tpix6qYaZN1kM5IWZL7TafINMqLnI90s7E5wOOSpgGuZWuBCo6NyqqoJO4LU8t45DvfxfPPPorlpUnDEFJ/BE2Ly514LvrZmGiMZtWUKAwF/SJV1VhXifqaOlTHq+B1s2BRkLmzf2AAQ2OT0iwh/hb0h6GHVUcXbrn1Fmzp3o5gMIKAPwq/L6zPTzYlRYNYJCxMBBu/EYwm25MAP4GK5XRqU0aFX+j9Cvhz3lU2hYIqY4NTyGRSqKqKCdDNQoYaaLqQyqTluRRGhQEqCBRHY/TbWpLvURaKXhpkM2oTRQher1+8UQhULMwnJE4JRihjwIYNjxiTS4xmQBuRAKR8k7DZOP9uDFS4choLcJ6ZnpmUeIb7E/kMdhSazmUbD9sYW1L3fAHXhoYlMieYEo6F4fWzIJPFigOosMUh6WiV4wojQaBidhbhUAg+jxeRcFgaO8bHxtYBFRxvtumCwyM3Q0bFPx1Q8U8HSJQSjDX/2ByS2KhYq/nIetNnXSMcjU+OvWwm8bTZEUnH+nUOa+33/v8CFc5C92bXW9f51QdV+nVNUduZrziPtfT+JhJIP9JMe801EX8Z0/3LeZnPRYhzuZG4cQIVeojGiNXrxdXLl6WhiEVPLQ7zA+sZFVJEMwfuPH3ndVoNFKw+SAUudNTIGFlzDnLvNnPT3pC58w8HKqTwaWWypPCncr3SCW7Md60U3PWACo0I9FRsw0bp/jqkg2yMJWPGwa5YNW5lG+XnSP0fbG3CsA1MIVEa0tiNzzjR+TJAhbOhTpu99PMSr21wDeW4DFihOIXWWoTNIXLAlMwxAITZlgUebOxowQTJ20T2hjmlSvVY/f+1caMCy2o8bkeEBRrk/NgwZiRzbBE/Q1Y0zZh5LVwuWXtOvnISLa0tqIhVlOT/xHRYTMhZ/Nd6kF0XZMYqSdUYdofeRO1yN/LN2kWv3+cY0Q59SIGZaw/fl65zfqaEWuk9LsfT6ieQXKE5skrvcA216wy3pzExr5UyALhf5sEq1eNoKjJ+G+KLYlQHRIKr1Pmv35HzZKNaQf0oef25b21q1BHA38km5L3WIjWlDj1S97AFdGV3WBkqBcosE0D6XO30rjetBKTYppOyLJDWnRRI0DFtn3H11yB7kXWmch5C0ELYl2RKikm6MmOs+oAFO1QGyiv5Prdr61IcT3L9jPk541N9FpT1yudfQSLRAiuBhBqXGJk0cy8sA0YkylwufPnL5YoyGRU6jvUZYhyjTNByfMjcnkCS5N/mHLXZj7JOVN+gzyCZqDqm2dEjoESxaHIIwp6U+TISXQZUUEBNTcS116dcf7SAC+dzPTaN6WwjgkhSm2dIWC4GxLK1Uhtn2uc8SzUOI4nGGo/MD/K7ASrZRG6ky+S7UjNU8Eae+3/LjIrg7rvxa2/di6b8KI5+6zt4pH89E6Hxtrfi/js7EVruw8NfeQzHZlfP3fGDb8CvvfkQDvQ0A7MD6D3xHP7qm89jYHn15zrveSfed1szMNOHb339MZxasx3np4Pdt+L+nzuELs8MXvjON/DQuRju/sW34k3byeC4zmt+AI98/Ts4Onb9j73W//qROzvL0kQluqpquskCodCePOCaHDtokBZJdgRDFl1etZiYiVVWGLPI8EErFcWdilKiy6mghn2V6jo20HIUemRzZv/OApAsxtLBzcKHopvrwRiHobWh01mdxjJ7xB4Pd0IARQMZ7YLgZK5UVQEZDDChE4suioK8CvCgplIy0RqGhR6vdpnbc+Z3VIdcFzVBxanjZ7ovSryTEs6ii5YaKlG7V7UT7fWz06kGJ2WzJOf7emEMOCNglAGZSh06ZVBDL7YGwCWT6Q2BCjXUXsk4PSqUYbH99ru169LtFmNn7m96ckoKx/zd6v7xPNjBzIIJFyUW7/w+RaNZGOF/uR0pxPsDkihQ0kcYGvPzIusjbAx2jeayaGpqRkd7u3SdE6jo3rlLunEyubQCGyzsRGKor6tHIBiSQlMmy+pZuZtFWRvs6PNKx2sqrWba7PCjfn1FZUylYgoq/cTuezXlziMS0u4/eiGwY5oL2jTNl6uqUF1TI8EZmQ8LBCr8AeRyaSQTS5LY0M+Bsle1VbW4evWqSDPRAHrbtu2orq5Ba0srlnJZNDQ2yrVi4ZjXh6Z9TOZttxG7QvkjJt/GrNwZbPMY+D7NKxcWF0QrPeBzYX52CpnZOYyeOYtAOoMtWzuQyFE7OyvXu76mBtFQCFWVcVSEwtINuZjheRfk3FncJWjDoU+Nx0DQLYalNIFOJVLwuTzoam9HZ1sHwpUVIhk2v7SIqdlZnL/Yi2RGgS4ySmorq+U61tbVo2fHTpH0YlwZq4kj73djbnEFjz75NGaX07j3LT8LBCNgqCt9CibAsdeAxeapqSkBKlzuAtKpBFLpJVy5fAlzs/Po2b4Djz/8MGLVdfi5d/w82tu7tEjDblQGuzInaNA3ODAs2+ru3q46oaagQ0kSjpWxayMi/USPin0H9ovWP6WjeG0YsPJZt5JdBKs4Jrld/u2pJ5+Uvx84eBDhirAY4dJrIZVcwfzMtOh4M0j3+AIiBXPjwYN45pmn8ba3vV0KZgpCFXH21ePweoqor2nAYqIAlzcAf8iLs2dOobOpA3fdcZfQUQlUsADKZ28psSjd8ByrfCZvve1WSaj4nBKUzLs9In/Q39+PocFB3HLTzaJvH49VoJDOYIlATGUES7Pz2NbSgkjQixzhCDcTLS96+6+hjZ3mES+dVZBze5Bx+dB/+Srqq6rEA0W6XrifdBrTU5PY0tao8i4uL/ou9QtQwQ6kU+d6Ud/ShvTKEjoaG6SzfGRiFtGaGJ5+4Rw++TsPIDk1iWIyiUw+jTQImLjhLboRjQXwlp95M9797ndjfHQUu3fvFiq5SqfQp6bMqOB9YTGX/6U8CcFMCczd7CSiBBzlkao1cJR5tww62CRSnsmiSzqICVTs3bsHofD/x957Bkl2nVeCJ21lpaks7137brSDdyQIiKREEoYAIXIkShSlXYVidndGs7OhnY0RSWmk2fm3fzYYExsbIRMyI1GUSEo0okiRIECAsA20993o7vLeZLn0mRvnfPdmZjeqIVE7owjuoiIQ6K6uynx53333fvc7jvY8/PlyTVHxD9UoLGCtKeG7GrVtW7/Kop+5AbQOGhwa1vrCvBEqKniNyqERKEtmUrMC169fu4xTJ48h2RzFkcMHMTw0hOtj63jrxEl86MM/haXVFTVJBweH8J2/+z4O7B7B+OQ4Tp85gZX5a9gz3I79B3ZjbHZJ85dhvwwa379vP/bsO4iuzn60tnYjFKbNH/1j6xYA/iBekvdqABcvXcDM9ATa21tkddbe2oHVtQyuTV5HV9cg9u85LMXE1tYCpmcvYmVlAvt37sfrr7+EfC6Dwf4hnD19Fq2pOB584AgGRg/gpTdOyGJuuHcI4xcuY2pqHHc/dC/mptfxwx98H9NLF9E/0IVPfvIz6O3ZhbevjGs/mBi/jl17h5Bu7cTYDQIknUi0tCgQO0TLnSYGDqfAfhUbyPRI5j5XKBCsWcB6ZgFnT72Ohbkx9HSlMDjUJ0ufRLIV4WgckXALEi3dCEWSWNvIIbuxjNWVRUxNzSCToaqwhOYYLW9apI7r7+/XfeOzyjVjZGQUcQZoIyTgjD7onBorK2tq/htjk2AakFlfU3aMclqKZaTiSXR2dIixz/2Te6+31JCiIhjAZi4v0FIs9qodrhuBCs68tfU1HR4HBgZ0IKcaZH5+CaFIEMkW7mtlnHj9OL7+V3+F9cw0Qigo4JnWifyPkvliviB1FlWE5VJeDQnaOKaSceXiENxvaUmiI51AZ2s7WhJp7d98ngqVKibn5vDGiXO49PYNbOS3ZJ8VZgZLdw+GR0e0jtK+KxZLIhblnk2v+Zw+TzIRF0ziGf/8HgFtgghNzTGsbW1gaXm5Bv431p3hoP0e1/FbrZ9mxua13re2JhBtsqBQq/XCyObyWtP5Hnw97iMkQXAd3djI6DCdakmp1uH94R5PMIKkikK+jMmJaawsZ1S/NCcJkLCGD6GqLA4DlfnF3+N1sTFbrBBo4tpmNSprlRpbu2TgO7+vjAqOS5LAlS0zdixwtbADYFWruvqW1nJcjRLxGJpp/RQJCajIyS7MAFtf31pGBedrc01REXekk1Q8oTqK6zFBD+VThDm+IZFWCPT9t1JU3K5xfus54x9an7d/nXdDA+oe/je9tlOE2qbSsN7/VwYqtu1R33Qiq18V58KtTf5bG+I3N9MbmsTOdsY+j7Hub/3yoySgwv2l/no3j9NN73NL9kIjUNFwDKq9Xc1OqfEC3Pm29sY1r2H122pe+ayXOCfYyFVDy593XSPaLtvOjzyjXb16BX0Dg2KC01Oe9bO3HLa3t/NjGbc0x/21NUydW8e2dq3u/LsdUOFPh3aSe+cr+GtoVHvUrsvoITdPy9rnc99ueAPW/3UlgDWGeZ+Nle4IegqB9b9rpA4bwsZzrJ23fehs7Xzu/O1rBEVXi6t5eYul9E231tuoKOOAjGfz4ue9sOapXae3bKG3vl2kt1+x+0SbVJ51xAbPF4zUKWvf+ln7HXP6FqBCM0ONYgNxSIhhHg/nBGsOvWutn2Cv5seH6y33S686YFPcLGQsB8hIiHXipOU5GEDAc6wIkk4xIAslRzxkw5frLPcrI40U1cg9feaMzppUsrE+yOZM5Wm9IXPe8PuCGruOCCeVgmP++wBvXhcJVObfz3OxEb94zWYBla31VHymAc8bVIayuc7r5bmGNZGfY2TkU/3Ms8D6+gY6O9ul+KxZ6bC/wmeUoASb1Y4xzzEmScEHVXPP4RnH1B1UerBG5VmeYcu0FDL7aX4uXifH0AARn5FR0lqgTCvaAKs5TauiiLIg1OdhfmEuVyNcqvfk+i+8R8yX9PknbETbfbfGv2ZfhUpoU+Gov1UDT1kH1a2ZfLB1433h79Oyk5+LageCJuGQzRfWrPy/1BJOzSIgjLkhUis45YmUPGaFzX8zqzDOIQtGFyFCIIsHKqzfph6KA1PMaszyGnyvjHPPQLgS/ugP69ZPn/3vSP4zQigJfnzEzDa5WePiM0LstWmHZqoSs30yhY3lAxpYQ9tunt9NxU6gyXo2sWhzLVeUYJE9n/Y5FVgfoJLHAB2evcrOpsmcOLhmuD3AKZc5jnQUMctwjo9lmXgQzNuEMQeRGR/KL3PKJG/5y/luIeBehWKvJRCJvVkqYrxC6f/LQMU7KoT3vvH/ixH4d++jZ78xcvQwOnmhNdetMKibMnHDJCprDzwXJnr2ccOp+w8aumqyRJPdWUPGFSnOK7BeWFhD3m+Q1uy3Qk29+QZ0wVBn8/avW1O5TbrhbtV/pY7e+sMC30syOdcAVJNQeQkBLXps9jWCJDW7JyLBrkjRYkSJGJkEriixTcAWbl80eMmcykGxR6xI9/Y63gvSy+08kkJJsb8P/FjGbLNQL94TLohkLnrU3NBWWgrVmRxc8PzGZvI858/oczOcVFTllw811AbiPO9obxOm4YKhuTXiDVF5MTPMM9EYgRU1O6iqIAsjVygiy4wKp6rwYdpscvD79z3xjBpjbMSuLi3rtdjoJBPCx4CzkcwGuw8D5cbHkGPeW/4um4T8YiOVhQsDLmPNCXR0dDjvP1rXbGmOnjpxHGvLS/IOHxkZqQEV+w4dVuBvPNGse85Nn4USlQ82r9nks7moYk++jCw2rCixQsEyKm4CKkpWLHkFBl+Xz0M8Zodq2pVwbMn2YJhpazqNru5uvQ7nIMO3mqM89BSwuZ7BzNQkdowO4+TJ4wgF6P9fxNiNcSQSKezeuxfpllb09HQzZVonKLE5m5u1gbOw4Dh6VgTHk2PWCFT4eeKfaYI/Y2M3VJjKWmRlEWuZJWBjCwsXL6ElGERXdzsyuTUF8xJwIFCRisfFbG1JJBGSjJShVUn5nLLAzBP4dOsM8wHYiNnIbKCSL6E1aUoJFsFNySS2ijkVI2RUX7hyWYHPiZY0urt70J5uU3HHRimLUX6+ZDKNZGsLAs0RzC2s4stf+4ZyCR79yOMoRZpQYiHnWFEcE44Dx4QNOdp6JJrYMK0gm2Modg7X376ChYUl7N29B3//d99Gur0bn3j2UxgZpU9/mZ4auscqKKPmyzk9NatQ2337DtykqFCzu5BXqO9fffkv8IXPfR533XMXKi5MnfPUpLnWANR1ra2LHc9nn9f7g+ee079TUZFsTQlEYvB6jnPIhWkzkyAQsjHhz7300ot49tmfdYUsG2gBnDvzFmLRANrSHVhZKSIYjSHaHMHpk29ixwCtnx5Tkcl1kUzBRCKuOQoCFYuLWoeYUaFDzFZW95Vjy0Dya1ffxsT4BJ742EdlnzI5PoV0PInmdAvW8zkkojF0JuJoClcRjAZkt1MsBXHhygSGB/rRmWK+SRGlYBhFARU30NXWik4FPkNB6eu5AhYX5rBruM8AoyCBircxMjqqgvvMhcvoGRpGbn0NIz09+r2JmUW0dKbx4uvn8B9/598ju7hAbyHkHVBBP/wwQkgmo3j640/iX/zcz6kxdvjQIR0yxI5yQEXjIYUgKNd9ZtqQvS6ggvka4Sha2lqlGBMgfxugQq/LMPOVFVy9cg1Hjx5GrNkDFSV6s/zTahAHattpxgp1rrVzcwvYvWePrOXqioo2ARUWVF9FU3Mz5qbHcOy1F1EqZHHk4CHs2bMP0aYkrlydxcmTJ/EzH/0wlleXteYODu3ED773Inbv6MXE1DjmF6cx8fZpHN7Tr4bwuavjylngYe+1117H7l17sG/vftm2tbV3orm5DS1pAhYRB7hbE0RNg2oQG9kCjr35BmLREA4e2ItXXnpR63QPwcloCL09Q+jp7JcCbHFhHItL13D58knMjE9jZvY6+gf7cNed92BlfgULsxN48P7D2LHnKGZWNvDSK6/i6B2HkF1exdLCLO566F5cujCFM6fPoLu/GRcuHEdHRy8++bOfVs7H9bcncenCNQwM9yKZbFU+RbkcR4AH1GgV0VSTsfQjCeTzHFNa61kAYK7APIIcujvbkVmZx6Xzx3Hm1BvYWF/A0GBKADpBguZYCxaWNjE2uYC3r09gdWVJh33PD+CU5yGc7C2u76l0i9ZY2nUNjwzjyNE71XyiUicWTyDVkhajbnkpg0DVchNUd3igYnVZoH21WEaLAyq4l90KVJhCMYj1rSzCtA5yqgcD16mosLXCAxVcJwiESeG4uoqF+WWpbXKFNbz4wxfwxosvI7exhnB1C6l4GLsGe9He1opkImHWF/m8QAnaTuSzW1r7UmTQpxJaW+JOJRaPRZCIURXBQ3FIlrOhphi2CmWcvzGNF19+FRcuX5L1HK32mlNJpFpbse/APjzygUfQ1tqNpmgKlRL3Y8u7IlBBf3APVHA+MpS+tbVNa/3KRgbLyiMx0KexRuW+54EKEhdY/3pFxdT1We35LWkCFcYgNXJJVAdZAswErfjlgQoSDdbXV7Ume6BCtYZspYICKogzjY9PKwfEAxUEpUXqKBrjVPV8IKAmC39XDN6g1TNstpmq0qwfVIOLuFoHKnifCVQYbceK80Z1GP+s8EgXRjs5NqFajUBFjGozKipIgthiuKXZrvj/5OmsbDE2ILJSxFJRwWBU/p9zar7B+om1rxS2ccvaskZNAPn5iggebPAoTFu5THagv7Ul23jP3g0y2HYBvoXFb4W2+8kfS47wzqbvuy/4DdZct5C57PcaCUUuxJkWgtt8+fOQV2f7GtAA75t/QRiBs5ZQI8/9s50LbrEouqWJrrlSQxvcH5wNRiPpSluVzwC85Xrt3FV/Yb3/Ntfof82iFLffO43T5hEPx/B2xLCbzn3+M+qa6g1z/2eRD1xGIQE4AuiJdBrFXE7ztnFK1K/LbGeOv/UW9uzdp/lrTNvt1TByFnB31asPPIO8kZVvII8DQtxHaxwea3S79+Fa4JwSbA5sPz9kB8R9xzVseR2sdfXc3KYs8dkJjfPDN8r9EPrnzgOnBurYudg3W/m+nklvzG7LM/D2Nh4HMha+bwr6Ua67Nhjouv3Tzfe1MbRxMZUH/2wjriwxkfcMiDPMxDHU/Rxynvsa3wYFhjHXec3WvGcNUGO518AvNw/d69qqagBDbb54ZQbXbrHT6+9D1rW5SptKhbWiX+N53WL+c+1zigCNowOAbno2XO/GADPLK+CXAp9DMCWAyJJl2cCePn0aw8OjAsztnpjfP6ewNYXZuzCypM9GiDbFUMxbaLJI7M4q1/YBsx5TD8OFcftnQg1Y2hWpEWvqBQ+KNNpD+XspRr8DDbnvqo9ChaObuwRESPKQJaS7GDatOdf4bwacWL9K85EgCLMLgtbT4lnHwBHrOdXwyADU2CZIJOVHhJkIRk41Sy+SS2KmkohGdbZSD8sVdXb9dm89WEsliwiQVGMwJyJgOU6ajwTSRBQxFw6CWb6XZIoJHwRuDfWacpHjGLT8BX4G1gH8fDZ3yZsLGqlGges2hxQQr5wPKk8sX0NjL8cQm6ucN9azs7qA48Czuyke2AOgpeOms4BygeYaP5fh6npRVD1wbdKzwCD5Ugl/+iesNe3rFz6b1X0wMM+sswXc1BxBmFFj4fP8Esio/YrqN4JNlmsiQIXqIdZATqFjzyvtoVk7e2sp6/FxHKT6lG0d56xTNrh+nu6J5rvloQn0cT03/d/9m9Y1l+/htyABlHwepEpxgA8zT5tjNWUSP4eRORwJ2WfOOCcHv8Lxbuh5fQ+ouKWCeO+vP/Ej8G8f7NfhhQdNHgAl0aqVeS7Is6EwYVOjJl+Sp2DEFn6pDBxzy1lc6iAStiY7H1JJzhqsL/g+fLBsY+SixYXSe+HVWWA+LMkWMGvGm4TOB/rdDKb4vd5vlibpq/+eBR4ZKGMyQ8eAcCy67W6qbaMuWEvv6wqEW3/Y2WMZU8FqYm0e/HUxrLn4WdHVCEb4zcrv5mYBZcyHRkaWMQCsyJLdkdgFtgDaZmse9z5cS4uqNhBbZH3lK2BFcld7rZqSxDWJWGRIsubAGbOlMhTfgiotWNpvrkWxZAykoN9ylv/R+iKfw2Y2BwZpU2GRzRdw7+NPuw2ujJmpKfnbczMmIk5JKTd1hWJHImqq+yZ7uZxHdmtT7EZugjt37tR8ZaO3WK6gKU6gorNW1LIByNc4+dabWJyZugmoqAQC2HPgAEJNESSScY2fjjcBMjub9Z7mS2mbJjcUFh8GyBGoCMleg+ACWSceqEi3tqhYkxrJeT56AMQDFeRKsWlMhjHtpbiR9/T2aB4SgKEFhHmUF7G0MI/lxXncsX8vTp85hXLRArcnJiYRicSwf/9+haeSXYummJ4xPs+0ifBMQx7mPZjYCFTY57Oi2rP5OZYMSGYxxSwJekzOzU0hhDJipSImTp1GNzNEykUsbjGDgpkM3QIqEtEmtLe2GlBBZgI9ppsTYkXr+bFqVoXbanZVapfNtU01U3raujE6OCJbl1grgQoDbXhtZO3Q1oQs1uZEAn2Dg5bJESPDk7ZUZKW0IZaIoxIJYnJmHt/+++ex59BR7Dp0FOvFCoJkuzl5pJpeqZRem9dAoCIWNhbqVnZdDfSxsWuycto5ugPf/dtvorWzF8984pPYuWuvnjs+VrzHPDAwXMxAjzVcuXwFBw4c1JxkIcUih/O6mMtilmHaX/ozfP43Pyeggg3OLQECmzWmqwqsSkVABa/NPwceqLjr7ruR7mjFamZVQfQEKtZWp+O9FAAAIABJREFUlqWoIFCBYETz58iRI3jl5ZfxiWefrRWxBGIunDuB5lgI6WQ7MmslNfboaX7y+BvYOTiCxx59VJ+FY0rGCZuPK6ursuyiLzvnywc+8AG9Jq9bQAUqavK9ffUqJicm8fGnnlLgO5uMW5ktjM3MoqOvG12tbUiRucYuWJiHAgINEZy5eAM7hgbRkWBwXyNQMSY1BYEKrlXlILAmoGIWu0fqQMXlq9cwPDIqpc7Z85fRPzKM3Noahnq6xYwem5pHa3cbXnzjHH73dz5XAypy5Rzy1ZKCe3lViUQEn3jm4/jkpz6lxhjHkMxujgcb7VxnG4EKAnr8Yog2g+3J2hHLKhxBuq0VbR0dFswo1Y1ber081x26/ulAhduPbtp/Gry/9X5Kltf6pfvz9ts4fPgIVtduD1QUy3m89srzWJwdx+ED+3Fg/yHEEx0oV6K4cW0MJ0+dxEce/5DWh+WVdfT1juDVl99Cb28cY5PXEApXcOrNF/HoA0cFHr5x8rIAi4nxMXzlK1/FkJtjPLw/+uijWM5sIRRJYMeOXZpr5nFsNhnrmwVcvDKOUKgq+6RCltZ3Kdx1+E7ZQ758/LiAQe5FzdGQ1Ac3blzG+PglhINVvP/RBzG/uIDmWAoH996BsyePoa87haP3PopMjm2BKr7zzb9FrFpBa1sz7nzgLszP53Dj+hSu3TgnJcPWVgFDw734+Z//OFpS7Xj++6/i0tUL6OsbxuDgPrS3DmvfCUaDCDeTrR5HJBJHIU+rMFrJUVVWRFaeOCG0t3QgT6ZggAz+DF55+QVcOvUiYmGgk4BeJoOJyWmsbRZQDUVRLDHM0HJUdBjSqd6H/kUUKMz1n0oCKigOHz2Kvv4BpNvbEUum0N7eKSVFJrMplUU0GkOEc5XWT1RUbANU0MaQAdjch72iQuquYBAZrlUxk+Nrb6zw3jQAFYGq9jDuNwQqWF9wH16cX9Eh9K3jP8J3//YbyGfzCJXzaGku49CuPuwa6EdLKimrOLLl2X1vTjSj4HIwuIPw3xha2RSJChxnPRaNNSMUbELQ4sOlEAvH4qiGm7CaLePNU2fw3Es/xMLyCirhIGKpFkSbqb5swkd+5iM4cOAoYk0tqJZDUqXwS2CJe159M517BNUOXNOX1laxvLJSA5e3AyrY/LhVUTF5fRabtBlMxQRU8PqVa4MQNrJbGjeqI/nFGodMTYLwa2urmkMEKmT3FDHwmuPEWoXB6GNjU1iYW5L1ExUVBCr475WCNZ78Hs/fEygeDqEcMNYlm1CsHWk1xvm1HVDBOUjQoMJmmjGIarV8DXhwB23+feIGMyosTJuKikiTnRMYpt3Y1JMKYxugwu5BEE3OqowqOjbHuO8aoB8QUEdCyz8MVHjmcP0g8/8KqNjmgFAzevlnAyr8RbjPpNK+hpbUwYR3ASpuali+CyYuoMLbTTRAAB6osMPNLUACL+cWgGLblnHj+94GMTKbnpv/sfHXthtyb4n7jlvl7Fh8o9KfEX9clYyAL3qul+j3bs9YjOH2DJJtALIar9Maf1HtwwP9/WqEUkHmG/B6kYaukz61a+D6w6RZI3rrl7rVsRH4PUpRHyv+yZ8l9ZwaK9HY+wzSvdXSyA0Yr4lgOMdFeQ2edMjzwjZzxQMSYgq72Vf7swe/GoiHjWdaA8dc41LBtZ4J7W1s6rkJBi7Yf+bV7kCEWxU/Dpzd7izv1Qi+sWrNTu/AIHuDmhrB3Aqc34FrzOo2uXvsm+d1hrjrK2hdM/sab3FUW4cbXAs8IdMTAo3UaANs72FKI16Bei2lkpE12dMQjmLAuBjvDDyrESitQc7rIonGWyapDeEeV42jGzcROItmh2Tvbw1v1mlqkErxGlR+F3MROY8t04BAEX/a+gH8fc/wl21qgX0Oa+x7b30qGsTiZ8OYTfWGm8Tf5/7A1+DZWquas1I0m2IbX9/7aQS+fJC0/30D33lep1qCihCqVJzVkzIZjCxgzHTOOQN7+MV7ZyQE9qwsP8Nfi59/nqTA37F8EXuWra9jhFtTDzhyLOPIBGJQ0eEyDJyaxn8ejrW3lBNg5vJhBdbq92kvZOPO6eHnBO9dI+HUckscQThoqhV+FuZ48LOyJvQ5LFKrOMCy5pziAQ2GoDvbdz/2Olnw3wu0G7ZGvvXoLMyeTxPvrXIjZINkagvecwO3rOdgvSOz9zI1Rth9HrtvBEX+4Pfqk+PTBCp8YL2Ua5alUsedWSMbCVmTys+5igWEWwZnFEX2ZxxY658Hr/IwEMpsn7z9lAevauCmXFDqwIzcCtw4cRz42qY4NiCJlrwCkxsyCj2oWAMw3Tz3NlacQ+yJGThqa4D/Wa1XTlVTB0Xt7Km59R5Qsd2y/973fpJH4N8+NFjbGIRSKmDHGuQ11YOajG5LE2PMZRo4CyMuMvJnc6igIcWumKLc1R1GOE7ctAyttYXWFwWGKtrCyrdS4BEZHPqzO8yEiIiaF6C8ltn4p7qAhAK5azi2Bz2+2aDh6ynYh+i1FTseteQCS0ZwU8zYgWqEuc2AF2ZFlhsDsRJuzqfwC40t2s7HUmiwU6HIZ9wFDwmFtYMdF3v5xdN/nNetjZdIqV2rLWY2vj7kyR+W/SLmFRbc7DgW8WaGBvGzNOn1/IJo0nrbQKwosfwP3luxMJyvJQtDzw7k4mj3wgo0HkIkISXDogZUeEWFochio1BtICukgvIFaPmUzRGw8NZPTmGRz+Pohz6mcGwFhLKp4Ta3dEsaLQxHlJzSpJUEKuwQXcTG+hq2tja0obGJwuY+P//mxqbekwzSjs7OWjHgFRUEKpbnZgRUDI+MKEy7Ggxg9779CDdF1BAhEs4bQiUKPQz5DOh9XSNfSL8ronhCsfEjm8FscqiQYCHEjAreJ8r4zPrJNmkWSjVFBZujAfP3503gz7BJwo3ZyyXpv00P/6mJcdn7DA0O4MyZkygVqwIlzp05q8YorZ/YqKKSpJkN3bBZ8nCO0QaLc4CvaWFTbBwkauAPr8sX3Jy3LJDImifwwjnA383ntjA2cR2J5ijaohFcf+s4upuasLAwiyzyiJDxWK2is61Nlk9pMlbjcURDEaSiYUTD1hgJ6lARcIqbElY2lrCwuIRiNq/g0p6OHowODEkx0ZROoRKyAwsVK5ToVkpkJBewurWBcjCAVtmlpCSlZQHEjIogrS7CIYyPT+HK1esYHNmNVO8gMmRnsNiGHYC40bMBxM9O1cLM9AwiATbsGUS9ilCgjOmJcUxNTWNoeBh//+2/Q2d3H55++lns3ENbp6KsLFicao3iYUChcwWcOHGiBlQoTKxY0PWX8k5R8Zdfxm9/4QsCKnyYNkNUOXdkyeGep8z6umzNzOIjCmVUBIO497770dbdrkYinx1agzGjwls/sZNDNsuhQ4fx+quv4uNPP63nxZ554PKls4g3R5BsbsHGZhXFSgCxZBNOnTiG0YEBPPboYzp4sxGdLxCoSCgPpRIIYWF+Xs8DG8xcf9m8JChZrJT0DNDSgPZWTz35JHq6urG1SYUUsJDZwHoup+yS3pYWxKKK0RZQEQg14czFa9gxPIT2eARB5n6QUR2I4O2r4+hqS6Mz3SoAuxwIILOVw+LiHHaPEqgw6yfLqBhFOBrBydMXMLxzFNkMgYouvf+1yRm093bgpTcu4nekqFgkIoV8OYdc1dhDtH6KJ6J49pmnBVQsLizgyKEjCrS1Aw/XgpKY3MzwMKb4mp7xeDyBSDhaA+KDoYiamm2dHqhoaOK8C1Bx5Aitn9gE/sdYP/GTNbIh/Z+d5YBYmrZGcU4xI+j8uQu45577sLZBoOK61pS2DioqmKdQEOvp4tUTuHT+NPbsGMbRgwfR0dGPSjWGSjWK69eu4tTpE/jo4z+t+XT92jQ6O3tw8vgFZDI3MD03hkNH9uH1l5/D0x/7MCqlEE6eu657s7S8gOe+97ysyEZHdmAzu4WpyUns2rsbFy5fVrbD3Xffj2SSWTFVZHObuHz1OhLpbqwsL+HKpYu4/567sGvHTjSpgV/G2NwcCvksTp96E5NjVzA/O47sRgY93V145NEHFED86rFjCKAJh/cfwvz0NaRbgjh61yNIdw7g1TeP4aUfPIdYoILDh/bg0N1HcPLMNXz/ez+SVRbXVs7hSKSEkZ3t+NjHfhrVchjf/ObXFQ6diPWhq2sIvQO96OrvRjLVg1gsJbCCQAVzB+R/G6hgg6BmMYDOtl7kt4pa20KhCuZnJ5FdHMcPvvNtzE2PI7fJgHA+l1U9c6UqyQeOGcbARSl2Io7VRaKHvQ/XiM6uHq3tZHDt2b8f+w4ewK5de9HcnHRABWXlzZqrPMhyjaGFlykqSmb91NmuDAiqIHzGAu+Ht35aXd8E2V78KhbME1tAxcamiC58HjY211Vv0XKLNdfK8gqWF1eRy27i63/zJWWfVAp5JKLAvXeM4sDOPiQIIkQjYMaDLAiCAQUp88AajcRcswcCKKJi0tk6HozEEQpSIUKmHbvYTYjE4whGYtgsMTA8i5deew0nzp2VqovqLwbgBkJVqc4efOD9siFDNYL1zLpCnfm+viel9wgGBRxwb+f4M4B8dW11W6CC1y4rEAIVLhdKjfVQGFM35vTsJZNUNdAijmsyWYTA+tam9iKqsPietHbk3kfFTCazrPqqJd0ioIJAEgkqBE2oJImEYxgbm8T87DwS8RQSKYIXZqtREpPVAmN5H1n3So1BhUM579RiZp9BwIJ7NPezgPJx7IA8vzirWjpBoEIdq7oFha9FvaLCasGKARWVirJyEqmE6ix5R2/lNWc9ScgfrrlHhXnPtrakqCBQwZrcWKrA8uKCgArW1Prc0bAsG24K015gk8wUFbTV4RmC90vAS60BZ6e1f06gorEp23hWdO3IH+P46NQsvrvYmC/gu8fextU1IE39sg1r/jagwHZseR39nKrC96h9k5NkJsv1ux1Q8U6Fhs0he6VGsKRGpLp1RPxBseH7/1SgwjfF1QByV+2V6D/GjRDITYsO2YWI6OUV7W5+eXWL54Y1XPDY+JhsaLlO8ODqmcnWnXZXYUiKNfr8vfRMWjef603lBkDj5rZvzQ6StYuRKJjVZPbDJO40kuUaP7/OtyJu+XvkCFu3USjo0msdQ/ud2vVtA1TYp3NMZN/018JiZDh/Zm0kNvJ3/LnbzrjWjL3pyw+WftZN3DpsV1sL7bPbXqqsINfI1DVrDXRXWPHWZm6mCiQyNQTvDK+H955nEI6pb3gy48usNA3s8WRF3zD2a5JNbesF+C/fd/HnTd8vEagtRwE2xZkLYZkDfj3zyhwDMuohxATxmUdkX47sWctLN2CJz7DIpI4tbjkKpgaxvg6Jg1G89dZx1UU+9Fuf3xFBeT3+HMkbSVW/VxcZ2GVDRyU4/80IKfX71wjQeDCbV+wbxkaaqDduda/cs+DVPj7jk/eEY2NNY7f+O2cKvqXsLl2finu+BXA7hQ4rZ2VQWg6Net4ET5wNUP3M7O+3ARxN0ZjOezbMAfes0X0kKkKXV5iQ2MYzE0lMOsK4vhhZ/nw/bzfGM7hsZ7V3GTHVW1uopohENJasZ6QYYHZZ2EKZSTDlVDWHDMv05Mf1PSIqSXjN3lKLSk/OKXtU3RwBbYebrPZjtqRIA/ysdNUwIq4H4zg3Nzc3dF85j8w6vh7kLecRFwDPNZP9GykwmYPS1KSzJOct5xXfg/e8KRbBH/9hfR7/8q+SMMZc0KzqXFsP6laCtPNi/6oWVF8xq0s+27w+Eud4FSI6qx/A+1QHvvz8MyUL54LNTblg1Gpwr5IhkGXAivUpGMIesgwvp5oyULEopw/WPKplqbJ1bhwiKJL045Q8vM8CUBpcTzw4IntA932FeDuwU3NTNlkOLOLovQdU/Dhb+Xs/+5MwAv/6gX41Y7jAbG5sIZVMOMa8C/BxC6n2fwEDZTHtuRHU0WY2uq0RyofOo6pq4KvgqkuWlXHR8ECqKU75sLwAjTlABoCBEER+bcE38MByH7hgc1G26zFJu9UnDYwpX4Q6tYBnjnBxMRmXbQKSBrpF2FBq2/g9G8TYFkTUTXXgFzP/nlxAtPCo4WzXa1fKJpztzLciqRagZu/B3+GBVj6LNT8973PIzY+2RlZ4sLjyIBI/KuWaLFrMSsoVL65wMeTePDa9ZMykpfb55FHpw74ZoETrDefT6EOiBFa4kVVuhYpI+64VAna/fEFApFo+xPStzhfM/omKB6opZAVl1k+DR+7CVnZLd4ufx0scec30mpbM0rEp2CyRD7YyDkpiFZKJzkZXX3+fbIN4sCXjkOxSZj14hJ4Hf17jW6+/jrWlBfT09RrzOkyPZqiZQ9uoREtCjQ4DsniQN0WFFCrkfxctcJqblfw0XUAmR5MyPzYUyHChVVJbW1qbt5RJ7n7ydygNTSV9RgVZWCV9Jr4WixtaSSwtLev7qWQSvd2daIqGceP6dQUmc9Omh3Xf0A6U8iUcf+OY/PcPHLgDyZYWjO4cRaqzXUAUWZsMLOUYav7KniYuRiQZiN72SAWN7qFJBqXmWF8X6EE2Pz/zxvoGZmfnEI9H0deawsSJ44hubWBmcgzprjaUwiEVGb2dnUg1x2XPwVyLZgZWN0XEpCTww4QI+YDnS8o6mF+cUYM3pIe4iu62Dgz29Qt0iRKoIKOBY8i1Ip+zIprcdEpgabnBJlAkhiCLJ/o6xuJqhvCEsTQ7iVCugPx6AZH2PizH01hviiAs9pgxkAhU8Iugzvj4uLIdwjGGr60gXC5heXoak9NT6OjtwfPfeQ4DAyP4+NPPYHh0FPlSWe+vQswVFmJAFIs4c+YMRvkzsgOLCJhh8UlLgLmpaXzlr76M//Bbv42DRw4hEKkrKlh4mdzdpLgMuiWQF+P3I1G88P3nEKwGcd+996Glq1W+5RvLGSwvLGBuchwrK8scYhU+LM7Ierp86ZKacVxrzCYmgenpSbS1tEmNs7lZQIkKrFgMl86fx0BPFz78wQ/LsoZFJ3NW6JW7TPuZQARz8/Mqth599LFa8ct5XixT1USg4irmZ2bx1BNPoKO9zZgzKGNtY0sKgxNvncTQQB96OloRj9oaX6hWMTk9i+72DrSKHVxFMVRBKRTG+PUJdKRb0Z5Mmow6HBLTfH5+BntHBy2cPRiURdTg8KByas6cu4j+kUFsrGYw2tcjNuG1iRmkezrw+snL+A+f/w1sLSwhkM0jW9xCrsrDGRAsl+UH/8STT+Izv/gZNSYPHzwkAIifg3kxPLQx3JaAFJ8pWmzpQBbjddczhTgXCFTwObK19magonYg4/pRrmB1ZRVXLl/F0cMHtf8aKYBz9WZLiMaGl2fq2SHY2bW4guPmJpyB6LTdu3jxIo4cOYqN9U28/fYV7Bjtl91OpRJCIVfGsTfewIVLL6J/sF92SX19QwiHeaAMIZsv4vKVa7hy+TSeeOJjaG5K4fKFcTUUL126gKWFywiGcugb6MCbb74Ohrhvrpfw+msn0dvfJgb58bfO4YEHHkNP7zAisSTGxm8AgWV0dDThzOkxhEId2Lv3ENLpFly4dFwgYK7Ag3lRGSAHDhzArtGdClLe3Mzh5NlzyOc38daxl7G8MIF4LIhDB3cjFuVa3oxkOonmRBpT00uYn53D+voU4ok8Hrr3HrR3jiCzVcKLz/0A2cwSBgZ6sf/oXbh87Qbefps2OhvIrObwvofejx07B/Gtv/sKBoda8aEP36f190fPv4WluazUS7GWANo7WjDYfweGhvcg2dKFCqLIMVCbh8tgAFtlAhUVtKc7UNjIg6UBykXlgLz83DcwPTmmNY77hA6rrg7h80MAmwdO1lhsyvPQJesA1+jh2k3bIK7DVLdxDWlOxLB77048+MCDOHDgkLJgGNQdjaVRZfM2AtV7S4vMMuKBuSSQrLurHRFEtO5771/OLwXIM3doa0Ofh/uyt6ajBzTXUdp58VqyuQ2tf0NDw4iEYlhaWsXi/BKqpQK++ld/jtOnXkO4vInDO/vxvrvuQKhaAkOym6lubAojRmBV4G8E4WBUNlW+NuPrcz0kgCpLg2CT1F7VID9fBEGu401xAeP5ShW5Qgkzi8t44eVXMD47jyqbDcoG2kR3Vyc++MEPYd++w4QqsbqyhnCwCfFE3JobDdkOBG64Z7C2pfUTSQbers83ilQTBqw24lpOGyKBFVIKhzA1taR1Ot3GzC0L7xTbsljFFjOY1jbQ1kJQ1oLptd60WkYFfZC5PhGoYL4Fmwps1FcqVNI0S2E5NzuDVDyFVCqp1+B7ck+y9UFtQWNx07YjEkaeTSixM9lwofKPwITPKjOGLCfZ3MK0fpf1i5pRZBzyAO9CN7XGucwJ7ic830+NT0p1yVrGZ1Rwr2RGRSN7Uc0g1rdR2lXGVRcSGGc2BRu5HDs2OZaXFrUXaZ0N81mwMHHWMv6983N2DvHWT6rTXKPG3yN/JvtvA1Rs70v/TwEqbvc7te66WKM+LMRciOrHn5vb/+8GVGwHDtyktODLurOKxtBtZdbkcbZPtwEqvJXTrQT8Wh5E3aO34dy0zalZa+HNDenalsr69hbQ5XYYjF2ysxWWtY/rOTsS2o9zXi8FqojEnAc7m0Yk9bCh55vpOvi6BIgq/92awXwWlxYXZV0q8gjPUS6v4dZx0h7v1Ab+2jwD37YHd+qt5Tnw/fynd+dYf7/YkJN6yyxV6uzghmnTMABeNc9/1VnfIbe1bIlbBkvzyINZHuX1Nke3ASrEw2+w+/JnZ69u8Nfo+wx+D/AMZ78+N0wjO7vXPvP2QAUnDBv3IQH/xqpn47ZGzFSjwc0P7Y0uj6dhdH0/whjZQXOGYC1NEJ1Nf2cJzXO1zyKKOLa17I8EQnkHiqoY9vZVv6c1lr3sjyw42xqjMqPSOVyNaHfh/D7PqroGNfTJhmcGERu2UZ2R/fPeaLNGIpWx0y0vQP2ZkhEk5EYhAqVZTh4/fhK7d++ukd8EZDgQXM1xOS/U2frq3zgXCFoEsW6gityyIKzJ7Od0I1ChRjUtCp01lcBAntHd/TWAyl7bzwMfxm1ET1Po1HpPDnDj9fKNZU8uwNysGUnS9a/DPokRFAjqUf1BIIN9LVMCiNjqnUEcAZRnBGuK0zmE+671DDhXOQfY7Gc9xX2We6i3Z7I+l9ms82fVNwjArK4c2OatwmX95Nj8PveB18XXJYmPXzxzcgoxf8rUivUzrzpkTiHF4fMgBT8S5wYVq5y76guweU4LXrl2RJ3lltlieZcADq+RYW2sWH/6Z1OfhXNDqgazNNK1uZ6PD43nv/MecGzZezGVh9UjkaYw/vgP6megz/6qgW0GspiKzc9bs7wyhxS+FsEJPg8kOogUrL4jnxrrz0n94hQ3Prxd4+csxmzsjOThz1qaa04hpZqnZr1k65i35fN9Nd//yRcMjOGX+j26x5YBwrWVtbP2+wbwXCCSsxIzkMT2DoGXDXPfMoMNrPCqu/eAih9nJ3/vZ38iRuDXHxzSA0CfO+9RZxdel0P6D6Kmp4otC7/jIiPlg/IoLGyHi7IhkI6Rr42FPmwywKjV0jXLGZdPwUWZnrI1IMNL7bTxcUMyP0RtZu6B9guIX0xqA+6KV48M671d9SKAQl59dpi0JpQMeXVttln6EtYXD2R38wDawFJoUFF4ewR+Zo++cjPiAZvj4v1BfZHgf942xqoOjrTzYTPG/7z34tPCK+/MxsRxk6bKhzJkQUX0SSegoQ1aGzhzKdhIJWruGIgKpDArGh1eG4LBfVHI9/ebv+61Kz4NwfW1lH0SLy3ka/G9TVJXUXNmK0eQIi+2p8+mEFBRyGP4zru1cLPZsLS0pCY9VQL8+9rKhootk3naRs+F32wUGD7XJAYoGYgMjq4WSlhbzcgiIxaPqTnIDZgbHpvu/IzHXn8NmYV5AypGDajg9e/Zf0DMwmRLUsHGvO9km3qgQooDuCLRKStqQAU3X9pvMVcin0OUnsnNzWqy8WdUEDkGAf9OCxABFSokqshns/qMvFaOdyKZ1AFmdm4OS/Nz2nOaImFkMit6jz17dmF+bh59wzuxtbGJY6+8BrqWHjx0SA2MkZ2jaOnq0NRlU8mY+DYO/Dsl6WyGs5FFZqj3PRQgUyrK3ocFChus/OLYsbii6ogFZiBQRmeyGfPnzyE7M4nM0rwCkjNkMJTK6O3ukpKiORpVqHZSAcNQwHhTU1zFYT5fwuz8POYZnF7MSf3C61pbySgQdaCvD92dXega6EcskcDW+gaKhZxUF7Emsu2rau4HxQiNIBSNIRhloyqMEO0sCM4V88ivr6KwvIoTb5xC5+heJA7ciZWmEMKOYdUIVPAzT0xMMOEb4aYgNjeXES4VsTwzg/GJcXT09eLF7/1QljVPEagYGUFOVhVNmu/GKDIAk38+d+6cQmT5umTVUmHE541gy/TEJL72lb/Eb33+Czh85xEgEnZZEJsqNuVHSlspWqysZxR6HGmKSm3xwveeYywG3vfQw2jrbcPs9BRuXLmKS2fP4drVK1hbz7gGDlU9bbIWGBsfVzORr8l52T9ABngXDuy/QxZbJRc8G4k14/y5s+jv6sIHf+rDasQL5GPzsjmqPIJSNSSAifOF1k+epSO1UKmgz0FLAwIVTz5uQAVBy0qA+QhZARWnT50VAJemb3nEGq9lMpciYSkawkWOJVAJV1AMBjF+YxIdLWm0MxyYnsnBADayRczOTmPfjqHbAhV9w4PYXF3FjoFerYVvT8ygtbcDr524hN/9wr/DxuwCkM1LUZFXzHoVwUoZqWQaTzz1JH7pF39JHvGHDh4UUCHrriKZwPkaUMGD1trahg5ZFnBrfsDcQ3kfPVChfe0mtly9HcE16J8KVOhI6z2MnaS4seCoA+52WOMafP78Ba0XbBZS/bJjZAjt7QzvBS6ev4DnX3gOHe0h3HXPvRjdwcMoLeMI6Fcxv7iMs+cuYS2zgMcqWJ2lAAAgAElEQVQf/xk0heO4fPGG1rKl5Wlcv/IWhke6MTV9g0dwPPbYB5HLVnHh7BWUA1mtzRcvXMeTT/4c0u29mJ1f1vVfu3ocwwNptLR249KlCZw5dxXd3b3KgEm3tWFoZFR2NrTHYy4Pc0O41l64eBmvvH4M2ewGIqEyertSaG+NIRqpIp1KIBHv1LrMHJhMJouzZ85ifv4K2tsDeODeuzE0fBDTi+uIIogXv/8ddPd0Ys/BI7hyfQanTl1UMPGRI3eit6cPw8PDOHfuDN5660c4dJA5Lg+jlKvi3NkxXLo8jvXcKvLFNTX6mbvR0zOAzs4BJFJdCAYTCDKDoJKXBLw12Ypyvozs2jounj+D55/7LmYnr2BrY13PlMBxd1+Vl6XDIPdzU1GwBuGzwLqBdocMtub6wDVoYXFReyn3vGgsjESqSSHoDz34Phy4404kW7sRT3UKBA5Fg9jYyAmo8Oxast97utsRKHId3BTwb4GStHbb0vWtZTfVxOFe4sPk+ewbUNFq+Tb5TVkGDg0NIRJqxsICMyoWQWjlq3/5Zzh98hW0xqr40IN3ozsVBUp57cOJWBQJWjv5Z0lARQQULwqoZJ1azAuoUDZVOAoEowIqeJ+pzgozNDvazBO7nq18sYL1bA5nLl3B8TPnsUkGND+TFF0hKc8++FM/g6Yoa5EVAStUhpDA4p8x/p/2VWyKs+Za3VwTaWA7oILsAdUrzBDhHszDaANQsaqspZiAfzsUs34rI1csYDNDoCKt3+GeJAVXOoX1tVVr+t8EVHAMYmAfoloNY2pqCgvzc0in0gIH+J5erWDWI1A9yu/RIpB1e4H+4swZK1mzpBGocHxh1aMEKljrUe2q5iKbMQHPNLSuIA/lnIM3AxWWa0Gggvu1V1R4oMI3OcQAppqmKSY15+LCkmzAaPFFIgN/j/aXpvCxfAqqSrz1k71OEPn5MpoiMVOzeEUF7fgUhHuziqIGVNQavv/445pvhL7jN25j+3RboOJdbKJuC1TYKaVRwOBY4r5BfXOGgNoY76KoqAEV79Ldf8dl1r02hFy408A7hsOU0v4sWd/3jBrjzoINXWb7zLe5kFsGvfZqXuzf8O7vBlSoocT9vsHfW4qK7aQkjrB26wdTYygUQJBz1lmxBMjM39qSQkIMcPdLHDudJp1NT5R5eHZ4QoFnPpeZ6Me4EaywH/MkP5eP4LIbG4EKrVNswUmp4hUsDqhw48x1q9bQds1Dbvw8rzW+Z+26nbe7t7xVjcQG8K1oSu1IyEad6xw0gED1I6O75w22RrrfvqHswRaXDWSKQ8ui5Pt6djPXIe//bkCH5SPYYu1nz7vNAPf4eHV8Qw6nZoZXKLgJ6pv0JEk1riGNz6e/Tj9P5HGv7AUDHWTlo4a1nSX9mJivveu8q2nv5r8fI0ciE+FT6gDrW6iJSi9+10D3tjZeRcDzmlQeUovU/fW5N6kPUlOwGPuUanU/gN42mvddgchSsdG5wayDzpw+i3379unPBIqpFKjNDZvYeiljeJtSgdfn6wjV/FKwuPyV2jhZT8ODXfw95Ux4lQfzOGRZ5Nw82Lx1QIVv8nrwwt7T1EJsWnubM7NDMhUE64dc1oh8dcVDwzXJbtOeK3+OVk/GkTOtNrBcAcuhYH4DFfEknlpmoVRMygszKyt+EVAwS2Bruvt+kd1DU3FwfHjvlLchu6J6xqhlOJgFFK/FgCkCkM5izPelqmXtqbX5zHvo1iXribOWNIBNYE2Q+WEM1LYx4nVw/EjGIgHTmuPMreFcZk0WlOKee61Ipaw5CaK5fA8pWZyi0c607Fc5Yq4j5Fl/h8ogU3iZurQsAi5Vujx/fum/kORoX7R+4jySkkREVoKo3nKK9zksm2her87kUuOUNL/9+LNnIwKnU0FxjgvMcHk1Ave8Tb3bIzyZU8QPZ1WvNUjPiJGIlffhSCFaVwnwuDBxfm6RkR0Jkb/Dml19UxEO6jWU1jPZqtp8qL+39TA57t5GygMXWk+UGevW0/cUFbdu2e/9/Sd9BP77o912wCALT/YwXExMZiTWgCvkzfnJJJFsuhrKWtGirEXM/bskdHo9Ay8ojxVa6h7sxjrU+83Zw2kgSE3tII86O5yTsa5FXfJ+Q+0bbZEsj2H7UpMLkGVU2EHFe8jJB5PNLw+6MDxabAK7Fr+A+EJRFlTu0M5/l3egsifcdTt/RzL0tRlqDOuHI1NgGKrrWQHGcgso4GmDwZJqRBiQwgVc8lJ3PVJV0CogaGFCvkjzIeViGzh0Xr6LgZA2OG4uYlLoPpIhgVoehd/YrWg30MQXQvK3dAiyNjsy2QNsyLq0DodQe4Sd941hiQxTFFCRZx4FgYmChWrn7f/KqPjIR2u2CNevX5fNBJtBbO4RqFhaXJLtDeeHz1SwYsGuiVtmZnNdQAWKZaxn1lAo5hVEy+a3R/WpCuCf33jlZazMz9WACjaZ+Sl279tniop0UtZWHCM2P8iQ5nvZhubseGTnZOCJZ/BRvaAAbAdUsKGWTqfM6qlgm7dAijx9yqmUSGnz4jNCL3Kb30Ft9mRr8mfXMquYn5vD7OwMMqvLqJbL2tR27dypZkTP4DA21tZx4o1jCFUDOHj4sFQmIzt3INmeRsSxUNho5nhyA+XcW1lexuryit6/t7dXoJBH91fXMmpMtbe36/DP6+A9YQMqs0qv8jgq1SK6EjGsvH0VYyffRFd7Gmu5TcyurekZ6GpvF0ARo3UG7aXI7A+yYdYssIIZJiur61haXFZmSSa7qfnCe0ewYqC3Tw1+Zhv0dnXJAqMtnZba69rVq0jFY0inUmhKNCPUHNPnZEMqwOKI5SCLJ641+SwKa6tYnZrB5fNXkR7cidThO5Gh1NT5/fIZY9OHX/ysU1OTKFeC1rzbXEKwmMfa/DzGJsbR1t2Nl3/wo5uAiiz9QF2BytfwDAquDwQq+vr6NHYeqFDhnM9jamwcf/21r+Bz//43cfTuO3XQbcyoUIHvbNiWV5cwPjGpZ7ct3Yq3XnsdzeEoHnn4YZSDebz+yis4+eZxTN0YA2XmbKwF2fAPk7lhzBI+R4vLS3qmqbRguCobQAxUPnr0bimK4q2tCMViOH/2LPo6u/DYYx9CbqugApVgK5thKxnawzCjYlHr5Qce+YDmFOc15zqbh2xUXiNQMTuHJz72uAMqCuDhaHPLLEzOnb2Awf4e9LS3yrJKklwyo+PNqJaqiJaraGKmUZhtxADGblBRUQcqSgFgk2DXzD8EVAxIUbFrsF/3+OrYFNr7OvDK8cv433/7f0Nmao5SGhQrBRQClDGXEGKIbjKNJz/+lIAKWqAJqMjS+onqqrzWGCkqtuitG0ImY178lHJzvMUmczZgDMUlaHoTUNHg0axDEBUl76aoqKpD68+QNTacrzm0tzkU5CaGcK25oSOk1nZmBF1R6PgOjfvVy9ewY3QIHR1tWFmew7e/8zWUyjncdfgo9u0/gFicKhZaABIoJvu6ghdfeh2Z1Tk88fhPIxJuxvmzF5FZW0Ihv4LZ8cvYv28HXnjhB7j7njtl4TZ2fRrr6zmEolWsrK2ikA/giSd/Dn0Do8jmygr1HrtyHuvL0zh46IBk2X//g+eRbuvFxlYF7Z1daGtvwejIMHp7evHqK6+gq7MDmdVVXLp0BU2JFIaHB9DelkQxu4pqaQuJOAHjGNZWclhYXpD3//T0goLe84UF9PXF8f6HHsbIjkN4/cRFjPYP4MKpY4g1x7Bj30G8/Op5nD17EXfdcxgH7tiNleVV7Nl1EJOTC7h07izGr5/GPffux8MPPYhKNY6Z2S0x9idnxrG4PIXNjWWEBZa0obtzEG0tQ+igtVA8jHKpimQsKYuhN15+BcdefwUTEzdQyNLuyddNRjbwewwtBaNUisGB9SF6FOtkos6z7m+DXy0b6sySYRpyNBZEazqFHaO7cN99D+HQ0XvR2TeMABvATVRE5LC0sFJTVMQTzejt6UA5a8CE3yO4x3v1xHpuS/OW+zL3V37dBFSUqR7cElA/ODCovI6FuWXMzS0iUCnjK3/xR7hw9nUc2j2Auw/sRDC/iQCfv0gQDMZONhnQLZaeDtARRF2wqbEcDQg0cJjPB1mAtPwLIxCKOaAiJtVIoUhFThnr2Swm5hZx8vxFLKyuSatE2yM+HZ2dXXj2E/8C7W3dWFnJOEUFQeM6U5OfkeNKNSL3/PXsJjJrazeFaYvEw/8cGMC6OMYciQagYmZmRcSDWCIi+yc2LDiY+VwR+XIJm6vraG1JoykaxcTkpBFQ0kmFaVcaFBXMqGDTniBAoUhryYpUj0uLC2htaRVQ4e1TfdOG1SdzScyn2Zr3BVcXkqEopmeZDTE7OJuNhzU35xZm1IBJa8+soioSEa1vrEZVY+M2QAUzKuKpuOoskViyVKaZKtUaMwaScO9mmDZrqYX5Bb0XzyNc/mhJtbK8aIAwQTsCFRECFbFamDavoUCgoqlZTZw6UBGyOvZ2QAX/4bbIA/DJz3wMbR1pfPfrL2L8BpUl3lKmfvL71C99DH0D3XjuOy/j/Omr7zgS3i4kWtaw2zR+rYH7zpPlHUf24sOPvw+Xzl3Hd7/5Eu57+Aj2HhjF6eMXcfr4pToNrNb8r2JkRx8efvRuzM8t4QffeRn3PXwUe/fv0O+cOXHR9hT3Xr5Bdes7e0WF/t2d89wKpP1dNiDbHIR9MGy9+W3nnRo4UrN/sl+uKS1ufS2npm/8tqeT6dx3y1jZ6Wj7ZrXP2vjHAhWe4Dayawjv/+ADmJ9dxPe+9QIqbLyBRJwoSgVjHStENejsY+zIVG9KE9Dh2StsYbb8Pba+Wbs1ikVuHcdG+yKvavDPnGeia0zVSOTZsg5QaLzcs/npX/s59A/14++//j2cefOMMYPFDr9ZtenHlTVC/bm2QGI1xt4FqPD9Ap1rfQPOOSh42nytSe886v2aXmMMax80ZjnPR/7nZffsmd2u4a+PV7vP9SZ5I462zbRUw7DRrozvRw+Zf/W5X9eP/+f/9MXar/lncTug4pf/51/BwOggvvnn38TpN05qPfNjRmshX5Nx3AwAKDuPavtU/rV19hZIUsEjH/kADt19CG+8dAxv/ugNDZvPUTDCZQWPfeyncMedd+C1H76KYz86pteResyRGsmEl32kcgvY8zDSokF0TlHk1kNv7cX3ETjkXABsvSRr0WfGG2Hh1KkzOHL4sFN4UimQVZ/Drs2CkK3JbudfNbwdUM+zjZwjZMfn2P1EyW+5YRwHb5vlsxcEmJXM+UFNeWUUmEW4ehBOlaTMBn5uOk5Em5DNMivQSLVs1HPP4DXI85/kV9dQbrTMZvNaje1AQFl9HuDw1ynLMbL+mUdD9YPLkWCjnba8n/6Xv4DsZhZ//MU/ku0vARE2362P7BrRJAioz+OCn6V6tH2K75+IJ5QRaPPEyKY3BWMzG0dWQgwqp6qFqghrmrOPJfUHOGb1fBeuZaxLfL6Fz3gQCYxEzCqZ/2bryXO3KS7s9ujPFZ7lDFwVqc4FUfMHuL9z/jPrlv9uNSmJnAxjtznIpYbnRLM4tjnL+cE5pF5IwBSgpixh8HgIf/KHNib8+uVfM/tn1pZUTZrFk+VUmKU6s1ioqmRuq1l7mWOJvR/Pq5wTtMfm/PIB2LQSlUrEzf9bFeoCVJivEQzKHUQOL85pxe9bskAXqGoWWXLZcIHaysUgAcmFbat/WSiY9ZWAOFONejCPr2muMVRnGQFEygvnMmKOLOZc4+soZdD4Z/o9oGK7Zf+97/0kj8BnD3W5gsWKLp8PIPTfBQtxYaE0zqRTZPGRXW++i3qQaoHPRI950KbUkGHAFWxmN3XAUFFF9JzBl2wEE11UEFNArGELZ7bQGxZbbKjKG5wLslBxMgdjAklqkj4uhfKI5KGUiDab9dzETGkgJULIArrJbBZD0W3I1ni3RhA3P0OW7Xe4EfIQ6VnnfF0u3GQQcHEoOPUJr0OhT2wU+sAkMU+4kUEsQW2obB1q0TLwRpkPrmCvH0rUcqgxs30BZ4wRQ461+cg72GSIagA7Vj5fzx8AvbJFShF+ljC987jRUdJnQUEqotyByA6vDLdiSDDvp3kW+6AkZWho4EyCxoVamzS/p3ta1fgViTAzMDFfkHe9gAkpKgy0UG5FvoCHnnxKCy+Lz2vXrume9w/0a2HObbLJz+Z+TiqflnRajW8dRAsGoLFYXt1YFzucPgP06icwEEs0qznoF/6tTXorBvDGq69idW4Wvf19GBodRfgd1k9UVEhuornEucu5zeuj77U/7FsRYeFgLMZYjLJJQ4ljJBQU45C2C2reap5ahgj/80AFm9dlqT3Wasg/5zobP/w5WvOM3biOrc1NzRcWLJw/nHOc4129PXquTh8/gUgghH379yOZIlAxglRHG8IuxFOe2hy7ZFJNDRaOHI+52VmNKecVQQm+x/rmBthY5X8cZ957Bn2zEcVDGIGdQmEL3ak4NsfHMHnmJAb7uzGzMIfLU9NaN9rTabQwDLdaRUsiobnZEm9GU6xZjaSVzBpWVteQK5Y0B5bX1zG3sCDwhLZUPV1davC3ptOIVKvIbW5h966d2LtrFxbn5gS0tCQT6O7rRqK1Bc3xBKKxpNj4tP0QS5i2cJtrKG9tYGFsHJfOXcHAgaOI7j2AZWfB4Q8PHG+TRpfFnieDIxJjoOoSAvk8NpYWMT45jmR7O159/mUMD43i6U88q8yKHBVJrtFszRZXaITCuHjxggAfPT/RCPKUFHNMc3Wg4guf+zwOHz0sZQgZpASJfD6FP7BduHgBi0uLiMcZFAsce/U1DHV1Y7CvD2fOvYUL589ha20dlYKBZ1yTLbSc67apovh93sP1jXWt67FYRLY5LNzYSD5w6DDuevB+DI6O4szZM+jv6ceHfuqnsbmRQyZjQAUbTQyOJXBARQXnDRUV9jyyaCSDOqvG5tjYGBZm5/D4Rz+K9jaOQQEIQ4qKRKoFly5exEBvN/q6Otl90pjTu78Siai5hmwRLc1RVENVxm3jxti48ik6aPdGwBUBbBZKmJ2ext4ddeunK1ev6b7E4k04ceoCegZ6NTa7Rwa1RF2mhVR/F149YUDF2sy8MioKlQKKAirKCFXKSKbSePLJp/DZX/qsAtaPHj6MHBVFNaCioMBnevPzyxQVNwMVdmAM6Vnq7OywJfLdFBWVKjIrK7h86SqOHDqIltTtrZ8a6wwPoDeq87arQ6yFFBBje2x8UmsCJdZXrlzHztEhWdC8+OJ3ce3GGRw+vB/3HX0/Uuk2sdR5sqD1HX2Bq4EQzp67jAvnT+JDH3oUHa2dGBubwLVr5xh7ja3VBXS2t+KFF17AM5/4ODKrazh75iJaUm2IxAKy6ltbK+AjH3kWIzv3o1yhrQWwODWD1374A6Rbw9h/cBc2c1m0d+/AydPXcf7iFbS2xjAw0IeOjnZcuXwJY9evy2bv7nvuRd/ILgSqZRRyG9haX0IqHpHig03OteUs3jr5JsamJlCpcJ+OoVJaQ1OsgEceegAHDt+Hb33nRQTLFRQ3VjAw2I+BHXtx7K1ryKxl0d7RhAOHd2rN7O0axeZ6FQvTs3jtR3+LXGEG7//AA7jn/kdRqbZgbonN+yasrmYxPz+GqelLWFqYQghBNDel1QTvGR5GS6oVTeEYTrx5HC889xympyZQyG/psOwPGfU9hs3YCMJRHgr5nwO1w0YmkR1GyLIZdEhVHcBsp7xAhbn5aQSCbC4nlBezd+8B3HP/g7jjyD2IJVqApgQ2NvNYJFAhKwl71glUFDdLyishsO6bLwrTDgSwkc/qgEoFpLcH9EBFMtmiRspWliquAgYIVISasbhI8H0JlVIeX/nSH2L8ykk8ev9htCcjqGQ3EQqSJBJAorkJ6UQzWlMMp6c1XEj2A2Gy990h3tdFdkBjnUV1gKnsqK7w1k+0A2SQZzZfsr1mJYPL18cwMTsv677NwpZIGy0trfjUJ38evb1DWF5aFVDBZ5zTv8Zoq1ZFnKDChESMzdyWgAqvqPB7iq4tbExE3rtY5GagYm4ug/X1DJoTESSSxvpj7UNrANZxVBZ2tLaLxDE9Pa29IdHWIkVFuVioKSp4gOd7E6golwPYyha1XtEeqSWZkgIponlhzEhT6ZChajYNJLzIlqDK2rqqmtKC0YOolo2gVFaOltokyqjgGsjnSsBoxTd6rDYSQCN7GDJ92bgOYHJ8gh02EPyKJ+NWC5PEkrU9w7NHfc3dCFQsLixqPyDZgXUia02CMLKsYoaJ6tmgwEX+nLewKCxU0MTMDo27y6hw1k+eqOTXyEZg993ObwQh2jtb8Xd/80OMXzegwkpnY0vzzwQz+ga68P1vE6i4ss3L3aa7e4ud0T90jvRAxcVz1/Ddb7yED370Idx57wGcfPMCfvCdVzG8YwCPf+JR5cH85Z/8ne7dnv0j+MjHPyBbs//ye1/DBz/6MO689yBOHDsn4OIdX7VMAv8Zb7F+ukV7INtehbYaG9kDACJ7NQDm+kcHONyu2a2xddL2m85H7zKitxtZ49fVWfz+77fDpDwhj782umsYT3zyZ0Sq+dLvf033eN/B3fjoMx/C6koGf/R//YXVWk4NsL62pjOKzks6o7Dz7Hde+7kKfVpDAVlqmg1sUnOUa6/PqPBUO/+ZzNbYRsV/8bV801JnQ/2AB2Vc6LhDMLTzu6bWp3/t59E/1Ifv/s3f48xbZ+3l2AS/6dUbBtoFqDe+Pp8rMqobM0Z+8V9+Gp09nfj6n38D16/ceOedagi/9ixtXq1+r7sDf/1nX8f4tYl6LoUjLUoh4pqB9mdPnLRmoNT+VIEpLHkbWY27En+P+Fcfkst1z4wZjLGsXka1il93QMUX/+P/aRZLDkzRnGbmpSc9uizJz/6bX8HgjkF860vfxMnXT1qjtFi0BmJNDWDAum+mm3rH+1XYRSqz0p3pH//UE3jgsQfx2vOv4ltf/ibuefhefPzTT+P0m6fw1T/+qn7+qZ9/Sj/z6vOv4m//6lu1sfPzRIRCB0j4Z86IMaZl4ue49+F78cxnPoHTx07hy7//F/qeqQyyNfIL4ROeqy0kmn2WEM6fv4g9e/bUXRfc/OP5loQKswarygLJyKcW2m4poC7zhD0EETLZL6hbKet3HTnT21kLENdzYrkIfBXLT7Veic+kECgaIPBnSknte2KuU3VYdNZF9f6OzWt7rnhveC6XgoFk1kjIxsG5fVi/xJYTnvUFmDkg73/5T7+BnsFe/OkX/whn3zqLnft34ld/49e0SfzB//F7uHHlRs2aVa4gUlpQlWDkWU+I0BrhFP/WKLe9ujZv9NxHHbDiGt9lghMG3qjnI2DBZZ267CBlRvFnHOjA96dzCZ0SeL/NfYH9DrpsNOYjcE23NUJjQjtuNtddfqr2P1cjecUQz4PevcQDYH7p4lpWhxLdwykLNJ4xbGx19nX3WXkbkRD+8P+2sxa/fv6Xtkx1IdsnI3iyr+HPzAJe1H8j4YI2SaQwWl/HnA+sBhGg46zR+QFJKOGabMoUWs2aG0JN+VCpKINRIBnJ1MqBtXskxUs4rPOvyMVSu9AZwfpj1t8z4NbXSuzFqbfqgucJQAioaKjZOJZS5rrcStvObO0wa7GCI4pTkWIApAdE37N+2qZgeO9bP9kj8JlDPRY4Tc9jWvgw/IV2Kg6l1IPXgPpKbgjLFfDZDvZ7JrWzLAV7CHmAVBnlUGQ+rDyYCNFWiI0pGAy1rVrhpr9b0ev98fi6Otw4BYRvtNv3KT00Homkhq4w4jULNXVSPM8k0EaoRcsa7N7/zW98fuMyFYYFHYstS+YXZV9O8s6fEzLt0pD43pLaOx85FUEq9kwBUjsY+QXLL/j+oOd2Qt8Y8AuTWA6OjcGx4WIo1gMZG07ux0WVskjPYOD91PeoNKkBRCqFdDg3oMe+VCS76l0bp0O5JWlzKphGYEMLrw4n9bwKfo9Ne44VfY+pqCgSsCgUsJHNCqwgaEHwgt8jUMEvWkcwH4CHbt+oRzmoQzab9wSHuDlysWZT3WTb6lqAKoDOjk4EKxaIzM0lmYqbL7zb8LgJcxE/9sorUlT0DfRjeMeoNjtKAPcduEOAVDKdstMnvTULJQXL0qeaEkc2uTjX19bX1HznmPA/zi9+5s0tZmfka0AFbSNMRZFTkeYVFQId3KE6t7UFhlcxOJZfzIfhc8JG77Ub1zQ32binhzgZklRUECgk+MDsAt49svObozHs3rULydY0evt7EUsm0BRvlpKCllosTthQkiyR0l1ASgkWKLIKWVjABu2xQiGNjVdTcLzZmKGyI51ulRVQPr+BnpYEyvNzWJ8cQywSwMziHC5OTGmO0VO6Pd2CSCAgRiyzVagS4WtmC0XMLixiZW0D61tbUlQwDJfMMhZ+nHPJeFJjzjFOce7m8xqDe+++R57zkxMTssYaGOiXh35rezuaEkllS1BNweBZ9lA2VpZRyW5geWoaly+8jf33vw/ZngEsUW2gQHgrWgRUuMMOG25rq+sIN4Wwtr6AanYLuUwGk9OTiCQTeOOHr2FkeAeeefZn1RDP8jCiBjTDCR04Kql6EG+/fU3zlc87VQy5vAXnUlExeWMMf/PXX8Vvf+G3cODQHQjR8i1rQIX3sORcO3/+vKTBLS0ptLQkEKxW8PLzz2NxegYrCwuYnRuXT3i5UBZoZQUafUn5/HFttgA4Bpbx/i8tL2nuVColNEVCKsxamf3Q2Ymd+/bg0J1H9bwODAzhQx/+KDbWclhdNbUAFRUeqFhaZqhrBY888ohbG01ltL5pNmET4+NYmJ3HRz/yEbS3t5kFQgjy8U+lWx1Q0SOgIiDVF7BRKOH82A10tHchVCxipL8XgWAFxWoVK6sZJJtiaGF4bzWIslNUzDQAFbzpFy9fxcjoMJoTzTh+8gK6+rqQ29jC7mEDKi5dH0d7f5cyKn738/8rNjrUBE4AACAASURBVBeWUN3MolAuoBAk06wiRQWta5hR4YGKO48ckc0a9xDuM7SXE1hdsj3EKyoIBHpmlLeqI1jV1dVpbLeaZ97NtYLds6oydi5dtIyK//pAhTGbCBDSOo4NFjYy3756HV2dbbhy+TxOn3kDg8OdeOihBzDSt08B5bJp1LxioyWASiCIs2cv4ML5M3jg/vvQ3tql+3vu/DEEI1sobmWUw3Lu3Hl86lOfwuTkNCYnpjE4OKT5ygPV/FwGd971PnT1DGNkx27tB1cvXcHM+BhWlsaxe3c/RnfuQGv7IM5fmVG2yfXrl7C5sQZUS1KZxWNR7Nw5ij179yPYxPWlCVvrKxi/fhm9XW2YnryB5cVFXL06jWIlr7WxtbULXZ192NpYwdjYOTx03wEcuft+XLw6hee//320NkVw5OghARULSxWsrGxgcXkCxcoa7r//AYQCcZQKISzOzuHC2dfQHM9heu4aHnzoUTzw4IexsLqFXD6CQJU5KWxGLWBi7AIuXjyNhblpWdgkW9rRmm5HZmUNx15/U2A0QYpqhYQNmxc1JhfXFq/QIQuXNmlc53RgtLBBrtkG2ru8q2pV9lisC/jv165dRaGYQzIeU+N/cGgQd951D+6670HlHJWb0tjczGNhfsXlTllTubeXQAWzida1ft8EVJBRJvJBDj09PS4A0awFTYHRotpgc8uIA7z3BCqWljKYn1/GemYJX/3z30dudRLvu3s/wpU8yrm8spia41G0JGJoTcbRwnwCKSS4XocQcgoTL3Xnv1mYJ5UBTQI0AjxYVkJSUkRjtG4iuaaEXK6EpfV1LGbWcX1yWv9lNrewkd/QuLakW/Gzz/4chgZHsbS4glCQAEBCQIUx4swm04eLU1HBPInVTEYEgJtqOxJSIsaA2w6oWFzckEVfMhXT52XJwT2Q1mqFcgmZpRV0tnWotuDeTHupZFsLNtYzKBXzNwEVJN1wLZKtWLaImekZNfPTiRSaacGo5oM1MmtABRUVIlk4+4CAsfK4njUCFXboJdPPgiMXl+a0/pFEwP1OQIUjGWnOOnUEPxCBCq4X42Pjypci+BVLxGRDwZ/dDqhQSRkKSFFBggeBimSc9m3NNWuchbk5PesCKfhshAICjkgO8czM/ByD17cHKvh8NYIT/3ig4nEHVLxQAyp8be5f81O/9HgdqDi1DVBxWxb6NiHX73KcPHiUior34+LZa/jON37Y8JP2BiMEKp59TEDFl//4266B7ZrX277udqqDxouts6+9DYpx612PT1jNO62faq/gX95Qgrpy4zbj4dUL1qC2HzdA6J1ftTajzk23/rvP1rOGsFcieDXF7YbCv9Xo7mE8SaBiYRlf+oOv2cf16g8H5NgZl0eRIFgXSeEUT9QaUGoqKSfAPgP5zUJcA5CtW29vn7MccW4EbkxtaFwD1YW5eoGMvz5zMPBqSrNiNmUlB6JusOzP1nzFz/wPn5ai4jt//V0HVNiZebvhtTO73S+//vu1hCQBroG6ndUqPvM//sK7AhWyTHY+9gRl1ewPBu33HFBx48pYDUSoTS0HsnLcPRPd3wdPoLTzdt1K6db7qv3CNS59M1P9VXf8teux8z2tcP715/6Vfv6L//GLIkPoLC+WtNnIiKXtA4oDAXz23/wyBqmoEFBxwllDm8bDhzt71rpIk1ID+jBzZ4DmQA+zWfb5B3ZG4X/3vO8ePP0Lz+D0sdP46p8YUMFrUUqFG8uacsmf610+ir9H7umr4V28wnseugfP/OIzOHXsFP7y97+sDAvuE74xbYQ8qm5KConms1nIsd47jzvuOOiyf9xsVUOdbgdBkRj4zPnmtexyCgZGEBAXiKB/L5k7hvk6mh2Us0jivaKqQPZRagYb41/NeweA2r5stmDK2GLYNQmvJLnlcjpPsSezlWX9bk189kSk1mCfgqom5nZIFcFmszX7rbdiBE8989qcoB6AzuHOkpxjz/f7n77w6+jp78Gf/uc/xsWT53XvvfLBVBq2dnj3An8t6uXI8YKvnddnU73hsjEZkM1sBa8Y4nwkCcXPY54tSwRlnIKE94dnZ5Ib+EXVAIEpzQERijlONi9FzC2WRBjme6uPxuY9SQGyljISr88/oKLRSMbMdmDWidVEXHdEunVKV5+tprFx6icpHBzox37JzUu1I+x65xb1xqy5b3VVFX/aoKj4hV8pCPAycNL6iOrHOFKxrsmB/x4QlEpFy6XZ1Nuz4J9RqkhNgeH7l77vSVIEnwepLFyWhPUT6/ZgfC3OPX4+n/vD665ZYTmwQ7ZWjgjLdxd453qtvnbha+kZcdZPIk47QrEIyK7PYO/j3WUMuBCBmbbzobDqrPeAim13+Pe++ZM8Ap8+0C2EkQ1FPihsmtVDo827Uw+5KxgYnOoZ/nUpqo2Aih7XGPchWSwCtDQ4j0Ui3DzY8jDlEUYtjtpMTBnBxUh/FivdZN5kfgkldYoF+TBHI8jlzIbDAxS8DtkvlenhzCahNfetaKsKYZcMksoCbnsh2zS54XETMmmcMfe9L7KFVhmo4dF8Sf5cWKHyIuTJZ7ZMXDx4ULaFzDM5LGSKi4oPsvZAiv3dXkMya4WVG+hjog8DOnifTAppFlYqS12OAzcTbpz8u6kszLLIVAIuoyNgfp5G0qkrKrSx1RQFVnyQQSFWobc0kK2JC/Thhi5U2G9YzKhgYWFjznwKHryNfZiT/QYVFWT1Eqh4+MmntLDTXoUyfx44LYMijFgkbgwM11DmZ9CcDIUsfJmLeTCANacCoP0RmyqFfE6Nyk6qLFzTh7/Hz/XGy7R+mlUzfmTHTgQEVFS2BSqIfjNslmGZba2tiETjGkey0i0LJK5DiTZH2l5sbZmiJoCaooJFlvdBbAQq5KsdIes3o0KsJdWi12TTg8ACAZdEMo6u7g7d+9mZWfR09+rPqXgLMuurmJyawNLCAqbHJnQwoiUU/f8HhgYRbIqokUSFBYsGFmb9/f2yRyBbhN/juBKE4GdYy6zpc5BNoM+WSNRUGFNT01hdWUZXV49sgIr5TfS0JlGcmUFleQGVUg5zS/O4MDGtokHZFLEYUrRjaG5Gc7QJyba0GqOz8wsYn5rGysYGsgVaksQQoZqBIAVBHydHFSsnEsFI3wDakinJdPt6etDGz1Mo4saNawiHAti1Yyf6BgcQT7UiwmYRM0dcQbsyP48Cg6YXFrE4v4Kddz2ApZZ2LISAZudbyecslWITzhgcVFtlllbF/l9dnUWVAFd2S0BFJRLGmy+9gR2jO/HUM5/A6OgO0PqJQAutNMg24pc/iNy4cV3zhYUy17itbF4gYqmQx8T1G/j633wVn//Nz+HQ0SMIN9ta6BUVvP+0jiK4wOwAMm9o1xQoF/HS97+P1196EVtrGVQCJcl9o+EmHYb53OWLJbHRM8qWYIMoIcCKTTfe+/mFeWxt0W6pKMswNnx7e3owODyEzq5OtPV045EPfhgPv+8xrGeyai5ypSC7eHllGcUKsLSyrOf24YcfrlmwcN7w+5RYT05OCqj42Ed+RooCsUIiASkP0m3tuHD+Agb76kAFlXj5ahUvnzktZnNTFRju6UYq1ayQbB1UKDu20vu2QMWFS1cwOjqCaHOzWP+dfV3Ibmxi12Cf1vCL1wyoePXEJfzO534D2cVlYCsn+5d8gI3dssK0qaj4+MefVpg2G4VUVNSAihIbiiYdZy/YAxW878b0NcDK/5+AKRVfBlRsXyH88wIVZWTWMlhdXUN3VxfOnz+L6alrmJy8jtZ0EocOH8TePfvRlupR01IMILFbrSVER5jTZ85hYnwMj7z/EYSq9D8OYGLyEkoVsuU3cPLkSXkuf/JnP4UzZ89heXEZe/ftxYXzx7WXs1H72E89iZm5FXR19WMpsyrAcfj/Ye8tw+PKrm3RUaqSqsTMLNkyySDbMjPJzGx3281pDnU6yUlD0knOyUmnk9OMbrvNzMwkg4yyZVtgy2JWiUtQUt1vzLW37CSdd7733r0/zv26+nOLCvZee+255ppjjjEiw1Gcl4Xrl89hUPJAePsGwcXdV8yRz5w6gevXr8JicUGAvw/8/byVz4m/P9y8g2V+3rpxFTWVpWiorUZOdiYIBPsGRSEgyA+BoSEICoqGm9kXjfV1SD17BPHRFvQfNAgdTu7IysjAvfRr6NO3lwAVtfUG1NWTcm9HbV0Fampr0Kd3X5HBKistR9bddIwY1Qf3s2/j2vVbmDp1Nnr27Ym6Rjuamv3h6uoDI0zCmKPfTVnZQ2Teu4U68WKqwcMH+SgsKFJylo422O2tcHKoJge9KKTWYm2JFgNkdmkpHwongzLW1unn/KqbGutSjmTRlZaWoqysVFhoPgTw/XzRo2cv9E8ejIRefQH3IDQ0tQqjQtWd2uHqZkZQkD8cLQC7hHWjYs5hAhHMiVTTgU1ilM4W5N8Yw/4RqBAzbZMrqipqUVFhxcPcTOzZsgZ+rm1IjA+Fo9UGR5sdnu6u8HS3wNfHA4HeXnCXTnrRUJKiN284PR+Q/M7ZWfIF8Xei2bsy8kBrO70qjHA2u8FE7Xi7QfLD6voGVNc3oqCsAnnFpaiqq0dNUw2xT5F5nDF9Drp36yVd5wY4C2CjWJO6sahd1mcBkw0G2Oxcs2vk5/83QEV1dSNqa2vg7ecuTCbGEILKbCTVgQoyKghUMDdiXuDl74OmRuY3NmFCKiNs1WlHQ2mLqwfa2hwoLCxCeVkpvD08JU9ys9C4U3UbSwGKebPm78DXSUOQyL+0i5k341hHOwsFqkFH8mOteFZBoKK1Fb4+3kruSQMq1LqniqQ6cMbQwbQzLzdPgGgCFczLTGYFVLQ2K8asXtxgMUyaYY3skDT/E1DBphXm42yaYGFJ5E81oIKMEjZ76DHXVqKaWnRGhRhpyz3zqANXj8R64flfFcLVfsaBRSumwz/QV7xcwiOC5b5rarDh0vkbuHIhXc5j4ZPTFVCx/zwybmbJ88dOHorI6NBOGYu7t3Nw8nCqSGGMGJuMwSP64UFOvjzX189b9kcFeSU4tv+MyLHxMXBYXwwangR3D1fJ+wvzSxAeGYp7t3NwcPcpTJk1BgQvLp67AU9PN/Tp36NzoeF14e+tVTWYOH0kSgrLsWnNHnlNYt9uuHjuOs6euCxd0OMmDUP33l2kEMdrVFZaiZOHLyA/t0jmjSpcq//1TuqOiTNGoaSwDP5B/nJszNfpJ3Xi4FlUllejV18+ZwxKi8oRFOIvcevo3lOor2nA6MnDERwaKHsYSqJcv5SOs8cuaPtHB3r1647h4wbDx89bfmetrMHJI+eRdee+/JzQMx6jxg9BQLC/jD3f4/b1Ozi+/0znuScP749BI/vDw9NdxrWkqAzH959GYV4RRk0ajqGjkvEg6yH8g/zg6++jxv5hEQ7vPimv6zcw8e/G8cLpNFRXWpEyezxKCkqx6ZsdWPz0XIRGhuDorhO4cPqSNBuNmzIKA0f2x5WzV3H2cCqmLJiEHv26IT+nAFFdImVu2mzNOHvivDCl+w/uK95NLIA/yH6I3Rv3d5ri6nuYwSOTMWbyCGTfycHO9ftk/8t971OvPSH3A39XWlyGafNS0C2xq+a7aEfegwIc3XNMpKr4WP7CEoRHheLgjiPy85S5k1CUX4K1X2zsPNeX3nhOvv/sP79C74GJmDp3EorzSxAYEgB3T3eJEXk5D3F451GERYVhyryUzgYbvu5Bdi7WfbpBnj9p9kREx0fJPpHrxO1rGTiy6yh69u2OyXNTlH679sjNzsXNy+mYOn+yfN7qj75Tm1QH8PKvX5RnffLHz5A0pJ98ZkFuIYJCA+Hp7SnHxK719CvpGDlpJPwD/eT5VeVVOLzrKDJvZ3YqP3SyDAxAbNdopMxOEZYJHyUFJYoxZ7fjo/c+lg8PCAnEtPlTEdOVvoZG6UK/fOYyTu4/KffJSjIqYiKwb/M+XLt4XeoTIyaMwIiJZKV6ynMKHxbiwLaDyL+fjwkzxmP0lNHIyshGUEig3D98Tl52HvZs3I3iwhLMXzkf/Yf2x5lDZxAVH4X47vGd48TYuXvjbsR2jUXS0CScOngSR/cc1RiW3KurpgU+Rk4cKePh5eMlcayyrBIHth3A7esZeOHnz6NLjy6d70vlgh1rdyD98k3MWjZbPl/5BNhQ+LAAUXHROHPoFHau24Xnf/ECevTpgZ3f7cL1i1cFhJgyfwpGTR6tjmf3ETmGUSmjMHbqOPl8nmPBgwLsXLsDD7MeqlqDeGFqJuQGAxISEzBt4XQZTxVjm3DpzCXsWb9b5dAmI5Y8vxR9kvvIsTEe5tzJxu51u1FaWCK1kBd//ZLMS2ulFZGxkci+k43qiio5n7z7eYjrFo+K0goc330U859eiIc5D/HX33ygZH2MRvzyL7+Sz/rDj99D8uhBWPzcYnkOAT5PHy+5T+/duocdq7cjpksMFjy7UFh9+iPz1j0c3n4IT766UiSjfv/6e+Il4rAryTe96SEiNhLLX14m15FATXlxuYArXt5e+PbDb2XuPPHiE3iQ9QD/9e6H0khF5sAfPv+jxLw3n31T6nXBYSFY+OxCdOudoOSGmltw/eINfPfRWuXP5mhH0pD+mPfEHIRFhct63ljfiPPHU7Hmk3UaA0A1DCsFCJ6JktfU632qeYY5hFI2YQxTDa1sBKYXp1rL+TydkSD1J0pDUQpclDnY3Kyk/TSOW+eYsbal1+40bFT9TWuI3bBa7f74WP608jbRQSmCTbqSiTTwmjifFADG+h/rXkpOSbFKFPNAA1+1pmkdFNFzJamZseivgSu6OTrH5JFiic5+UMeiN6mx5iN5q9bMrBpEIE0dihGtg/wK3OGc43WXxlrNPFvGW1NDkPxTcsTWTrBEV6JhXNU9ZgXg1/B6kVT7Qfqpc8788M3/JSOwNDFMbgSdYqc3u0ixWPZ/JkWJ04x/BG2m9BNpcCxOi0+FQqtZLFe6ear7TyG5SpaAEaKVPgKUb2ppEUNf0f+TgrtDBRZK/5CCZTRKIsPgrAqAvLFVL48KNarI7mIh9UvJJvChSzmJ7IlQ6mkQTs1qNymk8/XcxDQ1NihTPunIo0GQ2mwpSjrNkdTPyjxJyRk5GchSoBxVm3Tcc+HhOfLcuYHXaW8SCAVhNgobgOi16BmKoZQqvgnCrlFyxWNCk1MSqQGhyCkkXG0Aae6jPD74S6GUafRfZZKoNmH8vdJB5FiSesruAW7wlXSE6j4A7LK4qK4HkQDQTNNYrWC8U1rr3NypTawOaHAR47iqNUQBEywiSM5BEKqDZtodoqvITkhbS7N0z7fY2xSTgn4VbZR+asHwGTOlsMEub3azc2PNoir/2Vs6BHjgXBB2j4Xd1A7ZuBM88fX3k24BAiCUWaL8ET0bqIvNRFMHKjg2eqf6hXNnYS0tUUBFXLxortOQ+/sYFaRBsiuPXX0sFLi5qY0/j6WBBYNWdhb6SIGDO3Ele2GTTbku/cR7QFB1TYtQl8hhAYkPFrHYKcp5wYJSTU0tokWHPRjNzU2wtbJ43SSbTAIVLiYXYRw02myob6hGQ10dbl+/CZPBSaSfmNhEx8bCzcdL6a8aDOKBwXlJEIPd3UKZ1fS9yWShVAQLqZSC4ZxsaGwQhktjQwP8/P1FIooMEI5HY0Mj2lqbEOLjhZbiYjSVFsHgaENRWQlyyytkjhOo4Bl5ubnBy91DtPwp0UTt7LzCIlRYa1AjeqZGMcl1JhjILhiLWQAh6tUTDCILIMgvCAG+fkqyqtkGN7NZzKGp52utqhDwIjYmBj7+QbC4ucPJ2YWZoJxvRUkpmmpr0ChSUT7wiOyCMosbSmhGqnWwMB7xWkiCJV0vDlSWV4recm1tGRzNTeiw2cRMu81gwI2L1xAf1xXTZs5CbFyc+K2QgSDSLI9TxJ2ckJ2dLe/HcaXsFTU9CT6y2zwv9wH27t6FX735S/RO6isgC+8XzlMW+zIzMyVxGT1qNFpabTLf0NGGjOvXcOLwQTknJwH/GqRwz2IUYxEb7+oaGlHX1IgWu9L25cb5cfo64yoN0WnKauwALDSqNTghOCgAsbHKiH3UpMkYN2EKmm0szNVLiYLjZLVWo7WjQzoHOXaDBw+RjjMWiZksllaUyX1QxOtcVoYpKSlyjzDeOzkbZX6TvXEnQwcq/BWjgnJOJiPO30yXv0f6+8PMxIyGuTTyNTnDhbFRGHlG0KOiqUV1D3fVpJ+EUZGZjWgCFTQFz8xGQEgQmusbEBMWInM+80E+fEMDcOFaJt751c9gq6oSM+1WGhxTZIpSAB0d8HD3wuw5c7Bs6TKJN30SEzuBCoIUBI5ELq2TUVEn6xMNB/+OUWEwSCE3KEgBFf+CUKGxYMioqNEYFT01RoXeBfsvWk+1Ipps4DSQ/l+lI7yG0lloMEo8KykpR2RkOM6cOYKM22nw9fXEsCHDERQUDg8PX3i4Ur5HsSnIOlNJdLuw5K5eu4GrV9Lg6+OPtmaHdEc3NFaitb0aEZG+sp4n9uqD7t174tat2xLnIiPCkHH7CtzdLCgoKMfYMdNx/uJVmN280S+pP2IT4mGklA0cKL6fjSOHDmDqtKnim3Ip7ZqwMnr16oXKynLcz8kUEHfE0EFyPtduZ8s6npuTidrqCtgaauHv64O42BhExCbCi0CpAAAecHK4o6m+CadPHkCAby2GjhgEs5s/Lp67gJKC+0hKSkREbAKqa1jsdId/QBAamxqQlZ0tslM0ICaTJyc7C2NGDxJg+uL5y7h24zqWPzkXcd1jUGvjjPaD0RAAWxPNCykBSFC6HoX3M7B18xZkZ+YIEM48il2IVDp3cVJFG13CRi/+Sg4lRrhK/oCFcbML/RuUvBi7900uqoNf3yy6uqribVW1VQzEKcdHoMLXxwthYeFIGjgQPfolwyusGxob21BZUa2aQBwaUBHoA7QZBagg4K0bsFIKip9rs7dITOOawnnFdY7x6/uAiqioaJiMFinyVlbUIu3yOZw+vANR/mbEhHjC0N4K9leyuO7lZoafryeCfLwF8BbdZ5Eh1Dr8dB8OAf5MIhcqWsyUKuJml1JPHQYBrF3dPGVdMMFZfCoYr+ta2gSkyCsqkbWovKZCGFWMneMI0A4bhbraRjg6jI+ZNj9iyxG41IGK1g47rLU1smn/J6BCCulGKSaSSfO4R0VVVQNqaq3w8/eGi1nJUIjZYwdk3a6pssLPx1fyXzYTUPrPk34+9HNqtknOzPc1OCkgmkPi7uENg8EZ+fkF4t3j6e4pzBoyKnR5CqVfzPyafidmmcuM4+w+pIyBYlTQmJO5nCbZI805qsu3orJUwAU/X2/J8wlUiKmnSK8oEEmKFIwVBJQ7gIe5ucL89PR0h6vGqBDpjOYWtDBnl85kBTqobkcnYUf+I6OCXhP8jLLSkk6PCmmUMhrg5eUhc126Ddk0Utqi/CmcCWiQefwYUKHJrT4iBKjY+t8DFTMQExchUnbp1+/JHEjslyDnemT/WWTevq+AioggHNt3Dtn3cjF/+TSEhAUgIz0bZcUVSOzXDcGhAUi7kI7TRy9ixLhkDBmRJPE/734BcnMKQFmnkPBA3LxyB0f2nhbQYezkYZLzXr98S8YqaVCisGhuXs3AwV0nMGX2eHnvi2ev4f69PIRFhmDI6P6oqa7FtUsZKC+pRHB4ICbNIFBRho2r92Dq7LECVFw4e02AijETh2LQsL4oKSpH+rW7Ih9FCb6K8mpsWLVL7f00U1mOV+9+3TFx5mi1rt7OQWF+MZKSE6Xwei8jG7s3H0IinzNjjNwHpUVlqCyrQkFuEYaPHyyNONcu3kRTow1Jg/sImHDq8Hn5XVxCDCbPGS9r6bWL6TL/+g/tK0XLrd/tkXizcMUsuHu449rFG9p79IWXjyfOHbuIi6fT5D3HTB4uspIEQSjblZjUU8CK9V9vxfCxgzFs9CDJvXOz80WuqFe/HgiNCMb1S7eQfuU2wqPDMGzsIMm/eRw8h5DwIEyePQHFBSVY/+VWLHt+gYz30Z3HkXbuijSljJo8EgOGJ+Hy2Ss4c+g8pi1MQb9BfVBf1yAFRD5YbHd1o05+G7Lv3BfZo+QRAwR44fEfP6iYMjLmHR1SeF/y3EK5X1d9uFbuH77npNkTQCbC5lXbsPiZBejaIx55D/Jx69odxHeLFdCC773l250So5/40WKER4XhwHYFVEydR6CiGGs+26jfEnjpTQVUfPofX6FvciKmzkuR63w3PVMK7v2H9JPu8Tvp93Bsz3FExITLsfv6++Lc8VRUlFSgKK8Yy4S9EYr0K7dkvPoO6oPQiFBcPHUJV1OvITw6HINGDoBvgB9ST1xAWXG5ACHTF0wRMGndZxslLrDI+dKvXpBj+ugPn6Jvch/MWDRNjunOzbvIy8lH/6FJCIsKlT1ycX6xXL+4brHo0acbCnOL8PXfvlWSKY/JBHFMFz+7QJggd2/eQ/4Dvk9/hEaESCH7w999LLWFpc8vloI0i9M59+5j+Lhh8Pb1xpE9R3Hu2Hk895NnpLC+e+Me3ExLx8DhAzF5ziTxJ0g7fwV+Ab7oN7gfSvJLsO6z9Rg2bihGTBohe/ucuznIzsiWv4fHhCPtbBp2rd+FuU/MFRCCQAUBnKi4KCn6Z97KxO3rtwWUmTBzghzvqYOncGT3EY05pzFgOxwClkyeNxm1VbU4d+wcAkMCMXDEQPHG+vrDVfD180Fcl1iMmTIGd9PvIeP6bWRlZAm4wd+x0J964jx8/HyQPHKQrHOnD57E9u924NmfPYue/Xph++rtuHHhhuz7p86fipEpI3H60Gkc2LYPw8ePxIxFM2TfmHr8PEIiQpE0JAkFuQX47N8/FSaADqBTEtAvwA9P/+QZAW44DgSNho0fiqDQYBzfewwHtu7Hcz9/Ab3698L9u/dxNfUquvXuht4De+P+vfv4+v2vJKd6/Z3X0K13dzTUNQhAVZhbKO9Juic52AAAIABJREFUwMbW2ITsuzkoLShBeUkFFjy1QECID97+QBPiMuCdD9+RdfL3P3kPyaOSseS5pbIu8fMeZD6Q68C5e+3CNexauxMEHHgtOL5Hdx2Re4QxnQBWc1Mz3n75bY2ZpFhdIh1kMOLVd15CQq8E3LrGeHMLfQf2kXOrtdbiiz9/iYCgACx/cZl85gdv/1VYElzL/vTVf8i98NZLb8Hi5oqf//5nAshcv3QdN9NuYeiYIeiWmIBLpy/j8/e/lHvwx++8Dm9fL7lfOS5jp42VmLL9u13Yt/WAKuaLn1erpj6i6llc33XWmHT5a3UmpWJiV/LfduZPShLscZN7KdibjCIJreQtlbG4KIxoGxX9nmRjqK5C0tlQILUxpWCy8btHQMXSlarWx/ufew2u8SK3JuofzqLmITmIZs5NhogOVIgChgZWCHAhDUCUrtRYXlqTmUi7a/LyCpRRRyyAQVubygGZf0jTsaodcH+kmFeKKcEHm4eU3wYbO5SHLh+dEmYaC4UelTJOWqObNLhqiiDMqZh/q/xNvV5vUGbjCF8jsvysbRpYg6Sn6g9Axb/aC//w+//BIzA73rezc4w3mQQdYS4wUNBcR1GgZCOtGUUrjTi9SEImAOUz+Ct1M+m6gfIcTWtPZAq4qWGxnrRCasRxZ6TpFjIeiMYn28s0eSQxVNJkVFSwVEUXeS/NSEZR0FQw0V/P4qMU7bVAIgAITXB0EyB2m2sbJBWIVCKja9kp/TlVsNeDFI+JHWlMiHh+3LAJmqwRbhX4wCCpQgoTrYaGRtlYMJjy8//eOEl1UD46f904W5l2i9YgN4NiRqWCuWzsOr0qKONEQIESWapoylPg+DmLdrWiXKqgqbT3WBxhgq4vTgSRBKSRRYjPJLikpCPElMpOuS32oSjfDqFp6oGb+1ktKBPQYBBnQGVHHTfdlEewcVNqp050M2xtyreCHZmDpk4VKYXKymoJ5JRwcnV1l6BLmRjxhuBAUuPY1U0oiRxrajCz+MUiIBcjLy9vKRxWVlTIe/OaB4cEdxbvhDlgNiNVAyrCIsIREx+vdNcNQJeuCVLwoH6+yJRRroed8K6kRLaKJEslCxLOzvBw9xRvCWpTs+hPLWgWRrmxZpGfY8zCsfJ/aBeGh1Ba7ZSfaJZ5q3tCsIhEtU3KKXCRjYyMVOdEw+nqajQ21omxJxMCSmyw45VARUtrMxoaa1BbYxWgwslhQELXrvDy8UZ0lzh4+fjJfOGc4zzVC+C8smYXFk9cpMDBghvNpHk8LDhxXnBul5dXyKaGm/ImWxP8/YLEI6HF1ghbQwMCfX1RW1aB4twH0oH+8GEOOhw2kYqj8SV1tM0mI3y9vUTf3N3dGw/y81FeY0VeSYno0vt6+iDQ3x+ezoCHhWPtDn+/AFg0UzBqTDtZLKi00pTWWXQwc+/fl47u0OAQ+Pt6w9vNggA/P3mdm7sHLNQUp49GWzNKRBub5S8zTO5+cPj6oMbZgOq2Zri5sDivjOYIIvAC6Z0UpVXlMFOmqLocbU316GhrFvPy5tY26daKj0vA1FlzERIVIyakHe30oDCJaSc1uXkf8T5NT0+X+5bAisXNDTSfJZOFBqQ0vt69a4cAFT0Su8Pi6SayWBUV7LyuQICvL25cvYJxY0ajyd4KW30t8rLuYP/O7aguK4eLBm7SE4KJIO97xgSCPA2NNuWzY1bFMz6okS4anlpyR91xZeClmFvu7AZqbUaX2ChERUcjICwMs+cvRly3RJRXN8LW2g5PLz9U17DDs0N00zkZBw0cIPGCxU/qaxaWVcocp6RBVXkZJqdMkg5uJmE0O6+pq0NgoD8ybt9BREggwgIC4Cy05A7YjS64nJElnbddI4LhJgQ8A2qbWkTSy8vdFQ5Nh7it3SFmZgS/EuJjZJ1gvKFHRWxcNPVykFtQDD8/f9RVWREXxW65DqRn5iA4KgKXr2fivTd+iYbaCtjbaPjbJMegkmYajrtj3ty5WPHkChSXlKBvYm8B7vh3MsU4vgQoCchz7jCGEawlUKH7NjG2EgAO8qf0U6DqOH7M7ZMxprObl8Czw47aahuyMnPRu3cCvDxZtBa4+1+pR//32YZookparEQCOoDWFod4hRSWlMHb3x0nj+5Hc305BicPQO++yWhodqDD4KIk0eh3ZLejoqIKd+5k4ebNdOTlPURubq5I16j5o86jtbUZ9vZW2B0NAlzNmzsPM2fMRGEBfXZqYDB0oDA3FyFBgTh55iSiohNgcQ1Cv/5D0NTahB6JvQQUQJsdpUV5OHZoJywubZg8ZSRKS6zw9kpAbWMLrPUNcr2vXL4ATzczJo4bIx3yR44eQGODFS4uRiT26olAv2C4WTzgHx4D9kdQ+oeGzrxOZL9dungWpvYCjB6ZCC/PUHy3eg9cXFuQPCwecXHsSGa8IwBjwMMCKxxOFnRL6InWtiYUFdxG7v1rGD1uAuztrrC3WnDk8EFUlmdj0aLJIj9Gz4o2uy8aGp3RxEK0ww6brRYXj+7D5o3r5RjoqSQ5kHReEd5tfyRtKIxMAqiaRrdRfRX/IE0KhPGFeZHZTLYpWaFsrjCA94eXAP5+4jGUee+ubGyCAwJFPo4eIkOTk9GzX3/4dxmAxlagrLxaitX0+vB0c0FAgC8MTs4CnrFbWsWSDgW4woAW+yOjbb25g3+jpxLXFt4rjAUEMCPCI+FschEWT3FxKc6dPYULpw4g2t8VMaE+MBpULuXj5gY/VzN8vbzg48t1wwUWbtKcmNu0SvFcsXxMaHUY0OpkQnOHQ7yC4DCLDxrXRIK9zAECggIRFhKK4IAwmAz0H7ODAiEVNfXIzC3A/fwiVFRbUddQC4urCfFd4zBz1mzUNlD31wR3V3cYhRlMrzXllVatgbQskjKXYUwUoFrbYOo3pbMOVGh/E0CJ/0xG1FTVS8zw8fWWnILru26C2GJrFoYjzbQ5rmzgoGm8u6cHGmz1Aqp4entJsZ4MYyU7BVjMbjCbPQQkJtvJ28NLjsvbU8VmylvxmqjPUUw/i6vKXe3C9u2QYjhzDNGR1ioJDi0v1IEK5gVkVDDWkeEiG27NwLQzpmn5LOdTfkGB5LCeHu5w9bDArOX2LTbFNlU5qBoXXcLDSfNcY9MAWZnU/WduwWMtKS0RkIZ5Nc+fr+X8FMN3slsZo8sI0n8/UCHkMPU/eeh+AN8vLKSew3FbsnImgsMCcXTfGQEe+BgzcYgU92/fzMKBXSflOQQqju47K/Oe8kyVZdXYum6/PJ+gA39XXFiGTav3YOS4QRgyMkkAim1r98lzuid2QcqsMSgrqcCmVbsxb/k0RMdH4MyRi7hy4aY8h0bYoyYOwZ30LBzceRxT5hCo6I6LZ67i7LFL0sE+ff54YWRsWrVHXtOrfwImzRgtn71x1S5MnTNOwIbUM1dx5vhFLH16DsIignF47ykx1+Zj9sIUYRWdOnpBmBgyZBpYwddOmjUG9+89xK6NB6WiHhjsj3nLp8u827vtiMhVTpw5FgUPCrF1zW517MOTpPifmZGDQzuPywo3etIwDBk1ELeu38WB7Ucxb/kMxHWLwbnjF3Hh1GV5HX0heg/oiQunr0gBtRMs+GqrXMPe/Xti4PAk5Nx9IMyMp15dJiyJI3tOCNOC82LxU3MRFRuBw3tOyL1HsIIMhk2rlKxTzz7dMHXeRGGArP1iC2K7RmHW4qnCDtn49TaZn/ycKXMUULH2i8144gWaU4fgyK7jOHvsnBSmpsxJwaBRA3HpTBpOHjqDmYumCUhy4uAZKdKbHAakzJuE/sOTcO9mJrat3iFzt/+wJIyfNga52XnY+O02lY9IcUx9nf/kHHTpGY9DO47ixuWbAiAQrDh16KyAIAQdKkorsf6rrcJY4n239LkFiO0ag5OHzuL88YtY8dISAWD2bzss5zxtfgoK8whUrO/MJ175pQIFPvn3L9BnYG9MXzBZuv+38DidnKSwzwI/78Pd6/fiQVYunnhpmYAsO9bukp+7y1hOlmLwus83yNgRzJgyNwUFDwux6r/WSDHtqVefRGBwAHas2y3F5r6D+mLGwqnynG8//E7WRebUr731stytBCp4ztMXTpXnb/x6i8TPvgN7Y9bSGQIOfPfpegHFeDxPvrRM6gQbv96Moocl+k0vsXzM5FGYMH2sFOn5d453UEgQVry8XPYD//W7jzFi4nBMmD4O9zMfCMODe+CBwwZg+sJpKMorwud/+RIvvfEjMdPevWE3bl29JUwFFpl3b94jZtgcs6dff0o65+nFERQcIIyKnDs5WPPRGjkWAhWzl88WkOWrv3yFeU/OQ/9h/XFi3wkc3nUYySOSOyWatq3eJudB1sWAYQNw8sBJHN59WMVPzc+DMXz5i8vRpXs89m3Zh6vnrsr4/eiXP0JkbAS2r92BK6lXkTxsgIAilH7a+NVGWcdef/t1ASfIrqCUFReFGYtnYsTEUThz6DR2rd8p/gtkVGxdtQ1Xz1+VsZu2UDEqCFTs3bIHb/z+DQQGB2Hr6i24dOay5CrP/uw5xHeLx/Y123Dp1GWtqMsahhNS5qZg/IwJuHT6EjZ9tUGuW4/ePbDspeWor6nDyQOn5JxLCkvwyR8/luYsBqQX33wRCYndhClCQOPV37wmwNGGrzbIsfFzFz27CANHJGP/1v04vJNj1SEF/UXPLkZeTh7++u7fVE2lvR3vClABvP3qOxg6ZjCWvrAMGdcy8Ml/fCw1mZj4GDz/xvPCEPjmb6uEsfH6O68jNDwUqz9aLYBPj3498fTrTwsb5a2X3u6sI6lmXYcAP8tfWirMrA/e/asoBbB28tZffiOADRkVvAZLn1+C3Kxc/OXtv8renOP8uw9/K/Hs3dd/i5Q5KZi1eAauX7qBD3//scg4kd3x8z/8VCTV1nyyVmLSky8tF8DjL2//Tdb3IWMGY9KsCbh5KR27N+6V9xVAgjUrJ1XjYf1MeY2owrhaNBUzUzUgsy9QyURRnkn5MSipTN7bnIs8Jz4e1QIVRVg+SWM28NtOXx5NsUXV11RtjDnLpseAisVPNKuanNYEzWsprHtNdp35DmuUnBvCTOB/Uitko7BSSZEalxbxqKohEm+aoouoqGgAAp+iaouq7saH1Ca1vbQOiOj+KdI7TYknTUJfnshaGFURqPiggxWaNL1ukq3XVnUfG31sVC1WMVX1Ohv3nzx/5Sermsd1NowYhItfiekHRkXnivbDN//XjMCMWB+FAmoabjo6ypuBiDg3Rgxw/Lvo0xpUEJDA9pj8kAQAhVZoXWaqqK1MYog0EthQX1Xh3qYKkaRZiQeDMkPSqVQMWHwomp+iULE4pv5OKScRyVShjhRCIoyaVq5O59KPU2d36L4Tohen+WBIVyqDop3yT2rTxO5CtXlSjAbF1FBggd6ZwY/mJo4/s/NDdPhUNq+Zc3ETzY2hi2gL6rrKOjr+dwFPkF4VEEXaiouDFtB0lFbvnu0EazQzNzHzbqHOs2KgCNODAVpL9HjsYuJEBoSgyEoXUI2NGnsW3oVOp2nq8Xqzs11fiJTxmBpuATKYSBPo0aS4dBN0shR4Hixc0FibXbiUo6GhMAEKyj4RUOg7Ybxs2G22FpHg8WJXoBM3oNRbZpGD5kLcPHfA3aJ0itvbqGHJom6FdHhTPzskJEQKOCwqskhhdrOI1JGMo2aAye66C+fPwVpaDB2ooKY1C/rxBCpcnOHu6dPJkJGNPDv5CarYbGhoapJOf54zCxjcnNfV1cPF2SQFIY4igQpeF9K5vX14P7Wj2dak+D8Oh5wPOxbYCUqwob6+ES5mVzHU0yWCKAvF51qrK1FZWYHqaquMja+PrxQG3TWgotFWizqrFelXr0tHfNeuCVLAiI6PhbdfgFwovhcXLX6ueHd4eKCutgZ1taq4wvuYRVQWlFhcZIcXWUQEjshq4VcyKlqFtmmEB4vFdjuC/PxRml+I+upqYQg42lpQkH8PJoMBriyQi5+NUUww/b294enhjaKSEtja7aiuIxvFLt00rbYWeHuapVjn6+0Nb08fuJoVyMMxYoWI89nF3U3GvqKyEgVFhXIN4mOjkditq8iDUPOdzAELixX01aivRX1VNQxGC+xOboCHNzpcXdHkZEBDq02Oi/cD73VXi7vS4NeYSwXlxTChHfU1FWiyVsLW1CAd1SxKX7t0A/Hx3ZEyfRbCYuIkgWLXv9niLPe9o12TwIABtzMyxIgtOiJS5mNDc7OcJ9rtKMzLw/ZtW0X6qXvPBJg9XdFka0VJaQVoROtmdkFuTjZcXUzwDw5A/oNsHNy5DfnZmTCQHUWD9xY72hztUjAilkcfB/FJ0VhhetFGNNyhzNzFm4Pama3NUrhivsX5QVkpV5MJnmYTIiJCERoZgdiuPTB99gIYLV5obLbD0zdAgBAmdQQqeP8PGthf7jEfL0+ZIzSoJTNE+YiUYfKkSfDz9ZE44OTiAmttLYKDA3D71h1EhgSKR4Wz2Di2w+5kQZoGVCQIUMF7xgl2gwk5uXnw8faEr5eH3J9kWLAYyzntTg1XvoPDIUBFdGyMgI65+UXiq1JXVYP4mHDA0IGbdzIRGhWBtJvZ+N1P30RtbQXa7TbY7TbpdhF2GVmBZjPmzZuH5UuXoaS0FH16Eaiol3WI7EEFVFg0oMJJup4ZRhVQoeI+E192ggYHKOknAdYfM039Z6CiDbXVzcjKfIjevbvCy0vp7IoO2f/nRycvEhAWjUDPsFrrcOfeXVRYC5H/4B4Su3VB8oBkePmHwVrfBpu9A84G4MGDXKSlXUV6+i0UF1MyrEliRVsr6eRKF1j3OeK1ELNxR5OsEW5mCwYOHIA+fXohLMQffn7eKM7LQ3hoEApKChAZ1RXh4T0RHBaJ4tJCFJeWCthK8PTi+bMoeJgFV5c2DBmciMTEPqisssPs5oeg0BjpgDp18igy0tPgaG9Fva0DgUF+6NO7B4qK8mCtVgw0P58AhMVQMsGIthZKZah42NTUgDu3b6Ci+DrGjumHmKhuuHEtH+l3LyJ5WBd4ugehvc0hfg4OhxmFxbWotjYjMjpWYnp25lUU5Wdg3KQJaLVzrXKBu6sntm5ZC3tbFebMmojwiC5osjmjtd2CpjYntNiBnJwcrP74fZQUF8p8arY1Sh6lMyuVbjWbDUwC0pFdKps4ATJUTDVp3e1UaaacG7vm2WzxyBjZAJPZFa5uHsJsrKyuQFl5KZyNLsJOc3VxhsUIJA8agD5J/RHcfQBaOowor6wD+xmYDjE+Bgb4wcXFCdaaamkS0JsT6KnE/Ky5VVHRGV/4YCzVzbQFqIBD/WxrFQBeARWKyZN28QLOHt2DEC8josO8YSEjhGCkmxvcjAZYXM1yX4uptoebgOTSyWYn86AdtpY21De1oKq+Efml5Siz1sicVo0W1Og1SmGcICllp4IDwyQfYDxoaW1HS4cTcovKkZH1QIAKAmwtrQ3o0jUWKZOnoqGJgIYz3C0ewg7kQ2elEaigCaubh4dIX3F91uUqdeBR8lUNqNBBjMeBCnoHEIBgzsLNtepiVHlvqwZUeD8GVLBpgWtiQ3M9WuhRoQEVvOaUoCNQbjKZYXFxR3FxiQAVXu6ecsz0oRFwQrzQuFHnJhdyzAQquKluFUYEGRVkQitWhZbCsqulU6pUMSpa4e3lKb5LTgQ/Cf78w8Zdib+rAgZBa84FFrwJKBCoYI5PnXO9a1AfGyV34CTzl1rZlAN1M7uKRwWBCs4xBVSwQ1PJ63EM6ElG4Ej2DwCai20ikaaui7OwVpkH60xrXX9dD6vKsFntWXTzZrnvlBWtAiqemomAQF/s3XYcDx8UyrMTesSKhBIN4jd9u1eeQ6Di8N4zuH0985+idu+kbpikySVtXLUHI8cPwtBR/XH7RiYO7Dwuz4+Oi8CM+RPFJ4WAwnOvL5O9z54th1HwUJl4JyZ1F9DhXnoWDuw8hqlzJiAxqQcunLmCcwQq4iIwfQG9FazY9M0uObde/bshZeYYFBcQqNiJqXPGi3xT6ukrAlSMTRmOwcOTRPbs9o17uJuRg4qyamXZpqE6OlChHwMBlbvpWdi/7ZiKY04GzF8+A9HxkTgsIIRDAAV24h/Ypjr4+Ya65Ky+Lxs1aRiGjRkkLID9247g+Z+tlP3Sro37kZ9bKJ9PEGLslJHIuHEXqacuY9HKufDy9kBOZi7u3MjE3VtZnYwAekvMXDxFupk//8u3SvPfAaTMHIeBw5JknHhNR4wdLKyUvVsPyaHFdonG7CVTBVxa+8UmxHaJweyl/LkK677cIvdoX00KqaigBN99thFPCkMhFAe3H0bqqYty3BNnTsDgUcmgVNTJQ6cVUNGvB/bvPIz0S+kwOZwwMmU4hk8cjltXbmPvpv2yp+w3pK+AD2Q4rP5s4yOgQnwugCGjkjF++hjc5Gu2HMSLbzwj7PFta3YiIbErho0dgqsXrmOfnI9qIBg5fgjGThmF9KsZMp4rX16KiOgw7NuqgIrpCxRQ8e0n6zrBu9d++SP520f//jn6JfcRoOL2tTvYuWGPaq5wOLD0+UWIS4jFvi0HpEj69GsrBMDY9t1OPMjM/eeMxeFAv8F9hQlBEEKK/g7gqdcIVARi25odyL6XgwFDkjBz8XSRdVr14Rq5JxmPfvbb1+Wc3n/7b6CkF59zIy1dgBF2qFNSa9FTC6TD+q+/pWSTevzknVekcLtl9XZkZ+R0+g9w7zNn+Qz0H9wPx/efwvH9JzWfSiftsxz481t/w4IVczFgaBJO7D+Fo3uPCnOAEkArX14ha/V//Nuf8dIvfoTImAjs3LBLOvoXPDlPCtR/eeevnc2UBDaGjRmKU4dOyxiOnTpGWCWbv9ki49m9Tw8semaBsEo+//MXWPT0QgwY1h/H9x4XP5FBIwdhznLlJbF51RY5t4VPLcTA4QNwbN9xHNxxUH6nDLRVXv/4esR8gj+/+MsXhJ2xdc12pJ2/jOThyViwYr5cw41fb0TXHl3xxIvLpebz/m/e7/TvnDJvMsZMGSfsjW1rtuLlX78iQMXmb7Yi7cxlua+nLZginfqUfiKw9eTLT8r7/OnNP8mxcZ2bv2IBRk0aKbJZMu+l3kJPo3Y8//Pn0CupF7as2oLLZy/L+Ep+qfm7kJ0xYcYEnD9+Hhu/3qQpOzgwfvoEzFg0XRhN6z5fh9fffk0YP99+tFrAIK5ZK15egeThAwW8uHL+iqxzQ0YPBs3lyU754F0ap7tIzHjvk3dlrr31ylsYPn4Yljy3BGnn0vDdp2tlz8w1lIbrZC0Q3Ek9eQE//e1PBKhY9eG3wvLp2bcHnn7tKQVUvPKO8oUQlRHm9QbMWDJNgLzzJ1Kx+uM1su9gM8Yv//gmgsOC8OUHX8HHzxcrXnpCju+9N/6oJMna2vDHz34v4/lvL7+Dp19biSGjBmH72p3CjOB6x476p15dgTEpo7Bv20Fhp7z2m1cEuL155RYun0nDlfPXOgEHaczVjKGV94TyP+BD99bgPo9yS9KURCNxqhdIvahd7gmCQSJ9zeZabc2U+pJm6i0NCdJURwananl9HKiQfFfbU6jGF84LpfTBZsDHgYolK9okTyC7U56jrdOc+yz4M+8hMCD7et1fRvNt4WeIB4gGPvB6Sr4jjVxK/krFnEeG4mrvpnIB5Z+iPHR13xnFmFASntIkTYlnTVFG9vyaBJTKr1gHpY+mYqvoAJGwNjS5J3qyircHj1FUBB7lJ6pBWQeUyDbWFFA0QEf3vRB29Q/ST/+8Dv3wm//ZIzAj1u8RDU/rDuMmRm5CkUZSaKpQuFgslhubqKcytZOgReNtu9poi16aRvESx3oxTVWIpir8q005iz4EA9jxrorxioognSQawEEJKSngS3FRZxBoFCrNQEnLgeUcGBzEXIjditw0acV8vkLMiyQYcXOtAh6DtDARuJnjxoymWuwaJDLLDQ51+ERKx0kKVXyunJuYQKmgo2vYSdVQUFhNx08oZSqwMEhJ8ZibOw0QUcGPclAqwaCUjLRYCrJNvV6aQTLoqkVDtKhNJikasROex0EpEi6yPF9q+XLBYPLGn1lQ0xFw/iyFTQnCGlAh0l4CaUigJSuCxWF9cyLH5syAqGiautEPwRB3dw/pUmQxngiuLLYs3ra2qoJeu12ACermN7e2oLFFmWI3t7WJ9FPvcWNF85lxN8A/UKTCKMfE86qrV8bYAlRw3Cyu8hmyCFAnvq1VvBwIWAQFBck/gh78HI5ZeER457FSyojX6NL586h+DKhwcqL5MhDftascu4cXgQrFqJCNvEXJk3H8CK5wAWHBnEV2bp65AWa3OOeL2ezaucATTGBhgdedxWoughwTFvlYtNURehbXvTx9OoEhSizxM/n3yooykYNiQSM0NBSuFjdZvHWgoslG42crrqddhYuTCQkJCWIGzkKtDzuTHwMqdPkrFpA4brW1VmFu8Dw5jzgvxEyOxRWhctKrxg1VldXCuKDBtLXeKibCLkYjwkNCUFZQJKAFVSebG+pwI+2sFME83T3EK5AxwMVkEgPXYP9AAaucnE2oqKwWyZ7qqmphgpAuKwyYgED4+AZIJxi71zkf6BnBRI9zJiAoCHZHO65fu4aGhnr06JGAxB7d4eftDXeLu8hTUSbG5OKC6uoqVJaWwz0wGAYvX7SZLOhgDDEY5Bo6mwlwsru8RYAiFj7FrNXZGfmlRXDqsKOptgI1FaWoKC/VEgrg9o076JaQiPFTqaEar+a6BlQouRYVexg9qBVeV1Mj8lmUA7A1N6mEqL0d+bm52LljG37z639DbHwMDBZnlFdQTqkDAex6RgfampuQdfsW4uIisHvHVty8lApHW7N0+LLLmmalTGF4P1tr6mSesFtYzNHc3FQ3CRywaOa7cq6UwiBdtqVJpLY4BjT5ZgHd02KBm3TomhAVEwW/gCD06ZeMISPHwmTxgLPFCw1NlEhygL4ljOdil6SqAAAgAElEQVTJA/pLx5u3l4cksXmlSvqpsKAQVRWKUcHuW8rFGF3MqLRaERYWhPSbGYgKDfp+oMLNFV3CA+DhrHT47TAiIzNLvDo8zGaZK04sPsmaIpwoYUUxDmVl30dMPL1nTCgsLoGPjy/qqq2Ij42UBeVaegYioyNx9VYOfvfGr2GtKkdHezNa22zCkiKQw/nDAt68BfOxdNFilJaVoXfPXtIpLmCjmGk/AipI4WYBlmMpXcZOqquNQAVjNoEKxibVHfnINPXxTSTXgDbH/2GgQts8wGGSuXLi1BHkPryF2KhIDB08DMEhEWg3uKKorAa37mQi7cJZkS+rrKxCU1OzSGiw+KjYeqqTTRVXlb+LyEbybw61PrIwzhjq4+WBsNAA9OnbE3FRkfB0d0Fzqw3Jg0fB2ysCHVASNtkP7iIr6x4e3M9BTVUlErrEIbl/Is6cOY5BQ/ohIjocRpMPaqwduHMnGzdvpKGmpkiK2GGR3YSN16tnN1RUlArYwTlocDghtkscwkIjYTKxsKo6vVzMJhQVPkTqmV0YNTIRCV37IO9hPc5dOI4hw3vBaPDFrfR09Ersgm7deqK+vhU1NU1wdqVMnBPu3rqB0qIHmDB5DNpAPy/KOnrKvXdw/w54ubVhwqRx8A8IREMTgXoW6duw+tv1uHrxOJqbbLDWWZXkE9dhRdgEIUVpKNCYoswlWHRnemUyMJcBXC1mkZPzpewg7wdq3spGSMupHE5wdfcSlt/D/AI8LMxHExluzmYE+gXAw9UFdlsjevXqij5J/RDXbyAMLh4orWpAs53gpREWs4eMp5sLDcWrZT2WbjIHDbJtcs0Zz/UNk3SiaUA81zgC4vxZgK1/ACrKyyuRcesGju/fAW8XO6JCvRVbSmfUihScAxaTUdYTgg1k8LHLr1mkhijL1yiMoPziUhRVVqLZTgNxV8l96GHCYjj9F8wuziJZQy+B8PAIPPX0U3Dz9EZNQytKq+pxv6AYZZVWVBPMIXgWEYLZc+bC1ioK8HB1VRKNzOV0FqzVapV8jetNfXMjqq0KqFBM1kcSbf8dUMHchdeR119kdXgRuSYRqKirgw5UEAQlo5NyTw3NDWhubf4noIIFDBZeXEyuKCsrR3FRoTRTsHjg7uqmGn94v7JrkuMrXieUBVSsOwJAzKuZe9N4XHVGaoWDDiWxwI03gQrmQvSEYOcm49njQEWnIaTk3ErSSjEqHOJ7QkCB10bAkZZWYSzx2IQhrEnXsfHFZLZIPKfsJtcvD3e+TnmtfR9QQVkpSkzKGNLovaBJckmJQ7r0kwZUsDGlk1GhGZw+pkOhCum6YbLmE8eVdPHKmcIy2rPtiJhpE4SJY0F8/kRhT3z1X+ux5KnZCI0MFskmAhV9+ncXBgEBDr0bk/Mp934BNn6zE6MmDMHQ0QOEwbB/+3HZS8R2icDUueNRxS7+Vbvx3I+XyrX48m/rFMHOABDwSJk1FvduZQvAQdCBjAoW4M8cvYDouEjMXJgiYMemVTvlPu2d1ENeU1xQig3f7MC0uRPkdxfOXMXJQ6kC/IybMkJAEMoy8ZpVlFUJmyLzzn0FWGg9Ydw7kB0yacZYZNy8h4Pbj3WarE6bPwk9+3XDif1n5RqnzB6HOzczsU86+NWuYtiYZJFyolSTgEfa49qldNy4dAtzlk8TWZrve+RkPcT6r7chJj4S46aMREhYkOwL2AR2+8ZdHNl9QiSPZiycLIW9fxRN5J199eJNNNY3iQdG+pUM7NmkivYxXaMwd9lUMc/+5qP16NItFnOXTUdleRXWfLpJnkMppGnzJoqvw5pPNyqGQlSoFAlPHjol8oDjp48XoCL15BWcPXoR0xdORK9+3XBw11GRj7GYXDB03BCMShmJ9LRbOLzzmLAcKRdFVgSBg9Ufb1Cnr7bdEoOCQ4KEIcFxJUNi1mIW/Yuw/qvNmL1kuoAKZ4+dx+F9J9V+0skgPhsz5k+Wsdmxfg+efmW5rKV7t6rC9gxNZunbj9eqvXN7O17/DdkLwId//Ay9+ydizpLpwkrZvm6P5sFoxNxlM9F7QC/xuqA3x7M/Xim5PKVksu/el/0lC/wET+hVoasGcBLn3Hsg2vhMh1a+9oT8nWAL/TcIZsxeOkOAiq/+tlpreDTiJ2+/IuvPX3/3CXoP7Il5UrRPx7bVO2Xv1qV7HOavmCN7rPff+pvMV8aUH7/zqjSBbf9uJ7LuZHd22jE2LVg5V+R2dm3cgxuXbqrmxI4O/Py9H0s+95e3/oblLy4RVsn3PSjR890X6zF51iRExUZi27qdsl9Z8vQiuYe+78Gidn1tAybMGIcr56+KZBcvcEKvriLtVVZUhk/+9AUWP70Ag0YOxNG9x3F0z3EkDe4noAmlzjav2ir35+JnFspzju07iQPbD2nSNyy8co9sR2BQAGYtmYFefXuIP5D+oIcB3+PKuWtSrJ+3YrZ636+3Iq57rHTf0y/hoz9+qor3zTbMWjIdo1NG4dShU9j87Wa8/KuX0TupNzZ+uRkXTl+WuTNj8TRhqBzefUSYIQQ8CCB/34OSWRu/2KIUIzSm3xu//ymi46OF3ZJ68mJnA4d09Tscwo4ZNnYoDu8+it2b9mpd9EYBa5a/sFSAijWfrsPPf/cTBIcG4au/rsK9W1kyvs+8/iQGDO2PTV9vwfljqfLeA0cMwJMvLxfGwp9+9X6nh+l7n74rt91br/0Og0cNwhM/WoJLZ69g1YerO33Blj2/CMPHDsX6rzbhzJFzeOO9n4pk2Gd//hI5dx6ge+8EPP/Tp0W6+Tcv/7ZTBURvnp29bAZSZk3AgR2Hhd2ivAac8Iv3foqQiBB89cEqkRdb+cpykaX7w5t/VsVwRwf+/dPfyX3xq5fewS9+/xN06RaH1Z+ux6lDZzQmgxPmPTELU+emyPvvXLcbXXt2wbLnFiMqPlLWRTKPyPgik0q89tiooHmAKbNyNqMoVhbXejbW8vjEA4NKF+3t0sxIxQXWY/jgfcj5zxqCnCfrde00YzfKOkyAg/kzPUvZOKAaCJTiCD9fPDTJ8CRjQ1RDHq0Nm9c8atha8ESr7LHYFMdalXikUgKeygFsyBOwQDcYV3kqpeal7iL1LpXLdvpUcP/V2iYG1Hr9j3Uffc1WNUXVFChSmZphOz+D56mDH/q1ZY7EmCNsh8dyQubR1VVVIqVKMEn5e7AeqaQpdTko5mi6qbtibPD4HjVg8/PZKCKelqxFdpq9qyZx3Xj9B6Die0PPD7/8nzwCk8I8O70HhFWh6azpFCjeUDqlSAr/TJ605+kd9TqaqN+c8h4aIsgCKbvPpZguX5VslG5yp3f2axCFLC5MdsT8WjTdFBNDPB9aWjUqnRbIhJ5vlM5CFg51HT0GAG54FAtBdXmxOMCOXDGWFvkoJoFkUzBJU/IfLL4p8x9uqtRCqgAPpS2nqGOPPdiNrUlIMXgxyOhMACn8mxWwocblkbcG35u60MLCkK40gxRRqcbMY2LA0rNVOT5uNDXwgcmqGDPJJpoghTIUkuOX4gZlIFRhjBtPBWAQqaWkiAZOSIDTTIWEAaIAGo6xMhqn+RDls0yika0MwBVYwddx4eRioTaaijon8gr8SokUAhUs9FPDuo3m2jYxeeYCSEPtgVOmSCFMuim9vIUBQkSbsioEKnSpJC4eFppGan4b9Chg9wEDP4EO/uOmn0V+AhUM4gQqdAkwAhV8XE5NFaCChtO6R4UOVDiZTPDy9u3UWGbxgcV6mp0KE0JjdnDBoBQDC3csjnChrK2vkzlBpJ3HyC5HAhWc4/TZ4LESPOJmimOqd2eSKUHJI5HhaWsTE2ueOxde6kyXlBTLWEZGRMrcYNc6CxC8jgQqaq1W3Ei7AhejCd26dYe7lwei42Lh4x8oixfHR+ahXjRqZvc4zbs9BPwgG4WLKRMFq5XjWNGZrLiI2bxDFlwWm5hY1DVQbqoGnm6uaKipFT1/SjM01lqRfukMzGRduKlihJNQjTpEmzo2PFwAOpH0qqtHY32DFH6li4Od6C4WeHh5IigoRBgVnIeU7bG1tKK4rEyklyqrKQ9mFPN0yn6Fh4cgOjIMMZFR8PH2lQ5KAiHs3OdnNDU2wTM8HM2u7mhzMcNoMsOp3YE2XgNSaAG5tkaji9rUMQlzMSO/tBjGjjY01FSisaYK7fZm6QqiHMedW9no1r0Pxk+eivCYOGELtdlbxBCV96ColBGoMDiJDFlZSSkCAwLENJzdt5JFtLcj6+5dHNi3V6SfSBFvZaGR88bNXRVXWLx0tOHW1TRUFD7AySOH0NxYC4dG8+S8ojY//Wc474pLypTxlsitkXXjpmS8tM0az4/zltRTxt6WFpskXXwPmnyLtJ/JCE9XM1yMgIenK2JiYuDrF4DBw0ahd9IgWDz9UdPYjGaHk4AwOlDBOe/tya7dDuQWFcscLyjIR1UFzbQnwtfXRwBFZ4sryquqEB4eLEBFZGgQwoMCYSQASkaF0YIrt7Pg5u6GruEBcDcJvwF2gxH3su8jMNAPfl7eEt9tzZoRu7MJzhr7jMlv9v0HiI6JQXObHWUVleJ5Qo392JhI2XjcvH0XYZHhyLiTi7VffIPqynJYrRWoqakSAM9IOTAY4OrhglmzZ2LR/AUoKy9HYo+e/wRU8N5S0k+KUUGQiiAKM3wuDwSEGCRDAgOUbNs/ABV/v3w8BlRkPUTvXl3g5W3+38Co+OeMhPc7AYjUCyfg6mZHQnx39OjeF2aLLwpKq7Hv0EmcOHUS1WUFIk8k1G2ZtlxDCeKSkWPTwFbNQFfTkhXPInqfGE0yluzmdjEZ0VBvhZOTAwOS+mD0qKGIiglH7z4D4WoJEOm7mtpq3ExPw82baSKb1i2hG6KjItEh3d8G3LqThr4D42BweCD1bLpIQXV0tMFgakH/gX0RFdkb169dl/uZevUx0dECdj58kCPGhJERUSIbxGvEzRWBlqzsO0i7dBTDh3ZHv76DUVxsw5lzJ0Qz3sMSiZvpN2GtKcLI4UMRFxuHvPxiGIwuMLm44U76LVSXFWJcyig0UtawzQNOJn/AyQJrdSkunz8CVzcHRo4eIsy6hjoHLp7PwJefrUGTrVo8Z+ob67XCKlmJqoBnptcTm0GEmeYsQC9jKeOqr5cZ3l7uInVHhgPnn3h4kXFmYuc4Nz0QCTkXi7sUnzMzs3DvwX00MmcwWxASEARPdzOa6msQGR6APkm9Ed6lC9x9AtHQZkCrw4y2DgJMXvD3C4Sbs0MBFSxKa6wzWyOlDJ3Q3N7Saf6nN0JwvSZQSdkwznd+b2tqQRTNtJ0Vo4IyYg/vZ+Hg7s3wMLQgPMQHzY114q1T32QTbzLKDbkYneDt4Y4QetaEhQnbj+0xTDzrautRUWWV+9zBuOlJKSRnWQfdhInhKoCOF5mKzi64fu0K6usb8NLLL8MvMAROLh6wtRtRWduIh0XFuHfvNm5fuwJPiwmLFy+BvcMIo8UDLq6e4nWhd8HxbiJQwTWVUky1jfSaqFEx+/8BqBD2oi79ZDQK44fHowM6IhdoUmhVS5MNdTW1ilXI51qtEsM4j+tt9Wixt8hGlzkGwSnmPOwsb2lmvsZ1p0rMtD0IVFC+0mxR/maazxhzC7JO+N4ED/i1pY1AhfIro2/E40AF2Xtcz8TIWgMqxBibc8LRLmuHxDZNKkGYYowH7ITscCAvP18DKign5y7XQwcquFbwoQMVilFhhIlM1jb6plTCbHIRdgzzLK6fRcVFcl6KUaF81wSo8PLoLDw0FdrUfSGyW5pHhd55qck6qE6oR2wBPVKqwrbWPylABX9uFxAiIMgXe7ceRf5DlZcldI8VUIEd+Bu+2YklT2tAxZ7Tkn+woM08PS31BjJuZIlfxYwFk8S4/h+BikO7TsnxR8eGYcYCxajY8I1iVJAxs3PDIfGX4CMxKUFAB7IZ9m4/iunzJqJPUg+knk7D2eOXEBkThlmLJqOq3Ip132yXces7gEDFeAVUfL1djo1AReqpKzh+8KzGPlbXguy0pMGJ6DuwF5qabNix8YBIRon4m3SXQv5GhkLGTcWWkIINgGXPzZeO/UO7FEOEkk0EKvayg99B6ad+GDd1lIAgV85TU/02+gzsKQV6Pm/Xhv145VfPyv1w9thFmSt86P+vrWtAbk7+o4XN4RBwZcjIgQiLCEFa6nXxfJi1eApqrfW4knqtcw+lUwbIkOjaMx4jxg/GTQIVGw/L+8clKKCCUk8EIWITojF36XRUlFVitQZU9EtOxPT5BBMUULHypcWalNJBnDl6RvLcSbNSMHTMIKSeSMPxA6mYtWQS+gzogQM7jkg3t7OTUaR/Rk4cLpryezbul89PGtQHU3WGw0eaZ4RBNaIJoO1Ew/Y54kNx73YWevbpjpOHz+Ls8VRMnD4Ww8cOkYLqwd3HlDSLAxiXMgJjJo3A9bRb2LFhD5559QlERodjz5aDch1nLJwiYMfX//Wt5D7cx/2YQIUDeP/dDzFoOGWOpojnAw279T3sipeXisTYns37hdnw9CtKwmnz6m3IupMjHeULnpwjDAcWna+m3kB0XBTmr5gt8lSrP1ore8Vnf7JSfE0o4UQmBovOs5ZMEybNlx98K/sOxqY3fvuaHNMHv/tYzMcJZty4nI7N326XtY9AxaKn5omR8Ptv/1VTdQDeeO/HMLtaBBC4e+teJ4DD91r41DwkDeqLQ7uO4sSBU53yLm/+4Wcy4z5450PMe3KOgCdkAFRX1yg9eolZCmC+dT0DL/70WQ2o2IWa6hosf24JrNVW8evorFOK8oID1RXV6J7YTYCKy2evYsPXm7Xjj8fyFxaJ5Nvn//m1gC6DHwMhyK7g+aUR3Fi9Q8Zi0VNzMXT0YBzafQx7txzoNNXlvUhmD1kvlMS6dukmTh48jYf387DixeXoP6QvNq/aLteFQNKip+cJULH2s43o1bc7lr+4VHwSfvPKbwWQZ91h7rIZGDN5pDBCtq/bhhd++jx69++NzV9vx8XTVwQIn7l4skiXHd13HDkZOVj56gpUVVThzOFzcg/qqg/8nvJqeffz5f6WOpLRCc/8eAX6JffGd59vlCK6WpNY7G6T67Zw5TxMmD4GJw6expY1O1SjrJMRMxdOE9ZP6slLWPXRd3LNwyJC8e1H63HzKn19jFj50hIBD9d+ugGnj5yV9ZqyTk++vFSk1v70y79IMy6XyT9+/q4Ue3/x/FsYnTICT/5oiYAxX3ywqlM2/GfvvoqEnl2w+pP1SD19Cb/8vQIqPvnTl+LZ071PAl5641nxz3nzhbeVB6rsd9Uxk81DkJAgx6qPv+ts+nj7P38pnhKfv/+NgLUrX1mGnHu5+MOb70uDFI/7/a9+L/H2p8/8Gi+/+ZzEvo3fbMOBXUeVTxkMeOqVpRibMgq7Nu2TucE9PlUKyC4aNGKAgCTxCTE4uPMo1ny2SdWRtAZerm30wGHOIfUjO5sX6FGkGOesZbBJRpcrYlzifpOfK4wDMyXGVaOD3rzMXIC1Nn4GZcAVM0U1uFCthd9zjypNs2wY06STFNsB2Lb2kUfF/Cd0P1oFEgjrQhRbVH1RyTwp2XXGQNZWOD/ZiKbyEzJBFCgpgu9s0jSaxLeL8UqaJwxk+Sp/CWnA0pqJdRCGdRS9GVlfjPTaoJ4P6XLSekahszDE7028elsll5GGamlsUwx11TjK8WLLjmJM8Jwo4dVBVrHIV3EsWWdUTWLMd/gavTlc1E5+YFT88wb4h9/8zx6BGbEBnWghF2B2o0gnlWbQIgVPOKR7hXcuNz68yZWHgUIZ9QKsBC5uvrRAIYCFvA917ZS0EG9SBi3Vwc0OABWE5eajqanGjBBDbI2GpRDLv5fC0LvTZcOj0dJo4Eq0kcFQ9D21ri2RbdJMhsX/4R86XHUvCwYE/omBisUPKWJq/hJm6vqSziUOBwqw4CIkiKyY9CptPkF0hVamWAw0+zY5GyWR4gZVKGH6poiBk7QwKUA6JDHggiBGYp3m26ooxLFQnf4KxdblNxjkuQiJXIT4VSipF41nLdR5oriMcE5OtBBSuqeyKZNAz0WUwZsSGarjnMGaxWQTGRUCnygQRIEZTlqhVxV5VVelCqpt7cpkmGg6teRb29vR3NaCppYW0Uu2tTYLy2LYrJkSZFlkFmBGqIXcfNN8mObUzSpoE3WW31uY7aGtjcVVhVrrchMEIwTptpjh5uEuUg/cNHChYYciH5dSz4uZdkRUJKJj42QzrUs/sZPP28dfdUVr81qAj+ZmdRzi78CFwYE2dvprxqGCuhscIlXFOUs5DqUT6SrFzbr6ell0H++oE/pka6uY0RI0+3ugwiLnTKCiiJ2R7u4IDQmV4gGpjm4EKlqa0WirQU11NW5evQYXJ2f06NFDzluXfuK9qWuFS+JBrw2CDB5u8PLyFJCC//hZAsS0tqCqulIKRTYxqCJg5CZjx85H3u/s6OT8pWF2RWkpaq3VIvuDtlY8uHMDRnQIUEFdcTtpoNp4hAcHSWenJ0EMownN1GdvaFAyc2DXp7uANJwH4vHh6goCJR0GJwEDyEKhhAQBIQJedTQhN5KF44Oe3XvAn6CGrQVunh5oN2oGWy5meEVEoI4rusVNioxO1AJvaRU2GAsQqlCiy9cY4OXpjYKyMhjsLaizlsNWWw13V2cptOfm5iHzzgP07JWECVOmITgiGh0Gh4BGBCIJclBqhR2mBDXJGCkqLESgf4BslNiRIo/2dly/chVnTp3AL95QGq6+QTQD9xB2DuXmTDS7b2lEbuZdbPjmM9RXV8HgsEsMFekzAnrONEM1yzjW1NIXwB2NkmQ5iTcJ30cSMI2pxXjG42JS2NLaJEUuOJnVvIUTWuhF4ustbA6z2QlhocGICAuFn38IJk2djcj4niiva0RzhxPyCwoFqBgyOFnuCQIVNKvNzsuXOVpYWCBAxeRJExHg7yf3gNnNDaUVFQIwUfopPDgQUaHBMNipsdmOdpOSfqIeORkV7lK8NcHupAEVAf7w5VwjK68dqLLWSgIaFhIo8nM878pqqyTXdY2NqLJyrnvK3A4PDZGNQGbWA7TZO3Ar/TZupKXBZmtCRVkJKitLVScN2LFkgNnViKHDBmPhgoXy+vjYOLnfed+yo5nxX7p/aAYrQEWdYlQQqDAy/iud138EKh73qHg8W2BcbXW0oraqBdlZuejVKx7e3pb/30DFo0YbXfalHaWlRTh+4ig6Omzo2jUabq4+CA/vgvyCCuw7eBTnL10W0LK50apkApV1kypU80qx+7pdAa5q/VH6r3pzgpI9NMDZaJbiOMFce1szGhrqxGOkb98emD4zBSNHjoXZxRs5OfdRUJADq7UU3l5uiImJgpkd1a1taGxi/Hfgzr3r8A10xqABQ1GYV45aa4OAQ15+nggODUFoWAJIjaNJ+/37OcLwiYwMQ0gQPY9cpUs8NzcfhYWFwsxhgZa+Og9zbmHgwDgkJw9GtbUDZ86dxPARg2EyhKGouBIPHmbA4uzAtCkTpKEgK+chzO4+KC0uQk1FIcZNGIm793LQ0eGN0MjugNEMZxcjykuLkJp6HL6+Lhg9cjhs9XZ88clapJ67gjZDm3gi6L5PXL+lYYOx0uQEb083hAT6IzTQH94eHlJ4Zwe7p4eLeOtwjSeAIRspo0mARyPZIiayTg2ob7ShobEZ1rp65D7Mw817mbDamuHm6iHvGxLgC2tVKTzcTSL/FBAaBFcfX7SbzHCY3NBhIAjiBx/vAGFrcM3ga3lNOzoMAlrLfdDRoswEjUZZHzkf9LWS9wbXYv7c1NgsoCfzOkolsuO/pqoCu7d8B7OjCR5mAwoL8sTsvFVwCK4JBpG344wj0OXt5aXMA53aYW9tl1yGa6Kntw/aOhxobGkR/wbqPDs67PC0uIkPR1BAAAJ8/NDS0iB5GAEno7MbzO6+aHG4IL+kEg+KC1BdVYGW2iqE+nohqW9f1De2ICAsCmbvAHQ4K7BfMiWDAZWVlWqd9/RAVV2tMCy/T/qJ4VVJEymjQ35VXgwm6djmuqoDFdL0IYbg7QKk19bUCtjD15ExymYHyj01cv21t0jxiDGerBG+r3+AL1pb2sWHhXJJlRXl4lHB/EUYNyajdEEKU1iT72RuyfuA50IpLRYEhDHc0qY1EamYQfSb6zg32WWVJXJfEqhgoYJVHcUMfnT/y/fCjlCdgAQquJl2c7dIbsT1QoCKZjJMFVDBNUovAAjjiUAb5T3LK+DsZJJ8wI25bYcCKnheXL+YV/E8yNTgWFLukFGpqbBJAA6CY8wnpEAheSvnl1rv9QKiQIS6HwevsSZbq8dn7hEod/jEs3PFSPnwntMCEPBajZs8AoNHJIlUEhkRS56ZLX4Fh3efhI+fN4aPSZa/7dl6VNbebr3iMXn2WJTTR+DrHRg9cSiGjaY3wz0c2HlCrkF0bDhmL5ksc2TdlzuwaOVMxHSJxMnDqbiami45OD0qxqYM0977MGYuSEGf/j1x/nQaTh+9IKbfBCooMbbuK3ordKBv/x6dvg78HYvtfM25E5dx5cINLH12nsyFnRsOyvHx++XPz0V4ZKiADunX7nR6BvI69B3QC1PmTpDu+J3rKF3ULp4Ai5+eIzKquzccgKe3pzyHrIs9m5W80sxFk+W1505cwqlD5+RzBo8cgHFTRyLj+j3s3nwQS56dJ14Sx/efETCDD5oad+0Zh7u3szFi3BAMGp6EKxdv4PiBMzIvBEAQY+gSbPp6O556bZkYM+/edEB8K/hgx39giL9IRbHoOnLCEAFKxGNDgIpo8dggMPHdZ5tBCSn6ZZBRseqj9XKs8jkamLD6k41YuHI2uvXqgmN7j2P/zgPCREuZOxkDh/0v9t47Sq7qzhrdlbqrqlN1zlFZSEggCRBJBIkgDJjkhMHGYQbnsY3H4zTB34zns409Hoexx8ZgYwPGGDAZTAYRJIFCK7ZytzrnXJ6W1ksAACAASURBVF1VXV1v7f07t1vYnnl+6733xzeLYrHUalW4de+55/zO3r+996l45dkteM4RFctPXSxLJlrsUDB/zkVn47xL1mH75p14iERFJqOQ6ne86xK0H+vE7d+/29ZUNf+ayp/30ZozT8VFV1ygej6dSuMXP75bpM8ppy3HFe+6VED37T/8tWpJ3lc3ffx6AZJPP/YCNj3zGj70qfejtqFa54WgHAFojrUffetn+rzyylJ84OPXa19w69//AKvWrsRV73sH9u8+qPBw3t9llSW48eZ3S7lOwPhwy1F85DM3oqyyTDkWLbsPCAjlOX7z9R1SS/AeW7FmuQiGrvZu3PbdOzTe//qWDyv75bd3PCC7oCUnL8Z1H7xKx/TDb/5MdRuP6SOfulF113f+4ftYdcZKR1TsxL13PKC1Yd7iJrz3I9dpP/itr/27qe/TadzyT58Wyf3rn96Llj0HNKdqWptJ44JL1+GSd27Anh178cv/uFvNgiS7PvLZm9So+K2vfg8XbjwXG664EDu3NOPXP/utOUkgg5Wrlinc/cihVnziCx9FfWMt7v3lA9i9bQ8+/eWPI68gVyTE3uYWzZEcz8WlxSJ1rnjXO7D+svOwedMb+M3tzCKB1Dsf/MT7Zf30na9/Hzd9/P1Yc9aqWRLi7AvW4roPXKXzeddP79W1eu+Hr5XtD3NYzJbL5kRhBsEA/v7WLwrHuf0Hv0LL7oMaY7QLY8D43bf9Dq89v1mEGlU6b762QyoeYi9/f+vfobAkhl//5F79nt+YpMj5F5+Dpx5+Bvf/6ne4/q/eh3UbzsXvfvkQXnjyFe313/fRa3HuhjPx5ENPSyX0xX/5HPJj+bjzx3dj88tbVYtVVlco9HzrK9vfAmZzjF/9/iuw8eqL8NIzr8p6jXNzXVMNbv78h5SX+OJTrygTpr2tE9/5px+ovuAYuuUfPi2C5d5fPoinH3kef/u/PqPr+J//9kts39qsxo4Pfuw9OP3cVbjzP+7By8++pn38qjNW4CN/8wGd87//9D9rrSBJ8Pl/+qT227d89Ks4d8NZuOkT78O2Lc348a0MZJ9BVXUFPv8Pn1Bj0o9vvV2f8fff/lsRgD/61m2ysFu6YhE+9Xd/pTHymZu+ZOubw2bYyLr6zJX46Gc/oNB4jjO6B/D6/NN3vyQLte9/4yc6Xzff8iF0d/TgHz//Le3R+Rlf+sZntc/i+77rxitx9fsux9ZXt+HWr/9Iax3VM/946xdRVlGCn3z3DjQtqMf6jSSQnsedP7tXdeP5F58t0pLqp69/4dtaq9kMYOSQNbyxNiX+w7qF842nelRThZw8bO2nFbfXvCuSIEMHCbqVmNWw1+xruRV+4VuWUWFKDtn5+gPCHvjg8XGdszwPcxF58C6zGOXjqvcxvNtUrp7tpGe/NNsk7bJZBfC751nDCZutrOFYGJccUSxzlg++j/caHpPcSVzOmDK1XMMJ63cenCkeZtx8Y/ZR/J3IB15z5xBjjcOm+qDSmDUymwB0jmUvb+dDGKrD0dwpmiWH1cjB2oWuCFNx7ZP0O7mj+NUY7JEgaod+m6g4cZv99s//E87AxdUxTTy6qWnflGUhyuYVbyoA3mwsnAiKc6LhxCP5klhPew6LKRYJYv00IWTEVCpsh5Od29R4neViFd0E6REE9OEVu0hgnCyirKEI4FKebp5t9AmWGoBgOp/pfHLpJ19UWKSChZt62vRICaCu/6CzYSLkYmyl8he4WSKYzN+RihXQZJ5zCssNZskWx+Rh7Fw0Jtjz9dPkpVwLIxssO8PeRwqLrJBlJ1AOlrA8Bi8Eh4sjJ3Jvw8SiwHIfzPPVPKvNN1BvKAbZqUCcxM6zthIJpM5uy7ng8crv2imI+SeBpkDIh4xfLR6zXqZmtWVBQCxABSITKE4Ze0uPc3XKyirLVCUsdFn48bX0KSTjTvCC321yalI/UznBbAoqHWgDlfTIi1QSKy/aoHNC2yQFSrpwWk7Asv2JUwFAgNYCis1ugItJQh3Q/Gw+h+efm9fWtlYRIQWFMTQ2Ns6GVhMU4PV6fdMmDPWQqKhDfWMjfP4gMn4fmubNl+wvr6BQBIMIDyo43Pvz+0y7rkGNSxeULq9lkS9xAZjceHMcEQxWh5kWkaAyK2SZ5kgBdkbwfQoLiwV00lqM34dgvRfaefx4q7z+q6urUBgr0sLP/2kBZUTFCIYG+rFr+w6EfAEsWbJ0lqgoLCnXUPFCu3mOPLKCnabsQCQQQhUKF1+PaOT3oCc5gVe+tqSkTIDgxHhcGwZ2s5Okoa3N0aOHMc4QYY755BR6Wg8qqJWbMIJrhAV4zXguYlS7BLNQVhCTD3mauR+TE1psA352PIYQzs1BKCssNUxhUbHukSgVBsEsfRd2rpKwGBoZxvH2doyODWkDU1dVrcV/mgGyRTGwzKJip7CsHP6cPIxNzyCR8aszlkAprZ9IvLFA4ZjjvUrSkmO7sLAInb19SMYnMDrYg+G+LuTlhJGIJ3Dg0CG07D2KZctX4YKLL0VFXaPuM9rYsJs3mGVZLtzgsFhgFyyJChbJefl5Aoo0HjIZbH71Nbz+6iv42le+IquiaH6M7R8KaGeneNBHD+9xPHjv3djxykuygWK2xYxUShlk1BkT1TlmlglDbzlPTsTjUnYQMJctR3qumAuQbHX3STJJuzIOvSxMJuiPbvMnfeG50cnK9iOWG0VTXQ0i0TysXL0W52y4HEMTKUxMz6CtvV3A31oRFVkoyKNkN40Dx1r1/eeIiotQUlyIsfEJBMPZUsVUVJQ5oqIM9VVl8KfZsf/fEBW+AFoOHxHhUZSfp7kolfZhdHwcBw8ewsrlSzVfah4lzeIDRscnZTclm4FDR9SdS8C0vb0Tx2mHc/Qo+nu6FFbPvAWOYcqQkeEaEdL8yC6/M047HStWrMCaU1dp3PCepvUT5+K3EhUjpj4KU+FCIMy6ebh+naio+O+IClo/DQ1M4eCBI1i2dD4KYv/viQoL0bYOJXaKMQD76aefQE9vBxYumo/6hnkYGUni6OEuPPf8y9i3fx/6B3sULj41xfNHIoKFPJsFTDZt3q7WSGCgpxEVBrjzBeo3VHhxKBRGXjQHyExjaHhA1yASCWL1acvxnne/B1PxFPbt34OqqkLMb6rVcycmx9DT14PevgEMjTDkPCDyuKSkAAvm1aOmqlxKpT17W3DxxncqiyQvvxiFBUUYGR7HoYMHcfhwCwKBDBYvnIfqmgapO0h6DPT348DB/ZiYHEF+Xg462w6hqakAZ5+9VlkTm157EatWnYIg6tDeFUc8MYrB3qOIZqdxySUXo29oAoeOdaKj8wj8MyO49GJ21vZi/94uKY7YpRsIk3guQMfxI9jy+ksKjU9MTOHXd9yNgYEhTGbSsq6TrZOf6Rl2X1aUFmFhbTHqqktRXVWJEmb7sGte55jdUZAileuDaq6UEaKyJPKH4cuKyBItkUqLxDvW2oFjbW3YsbcFrb0DyM3JQ21lBWqqSjE82I1UYhRnnnkafAS6K0oQKSxAhrUDiePcYpQWVcMXKsTwMDv/83Vv8FrwGvLCU1HBGoLrhLdOe4oK3ht88O9joxNaizmPc11hvs1gbw+efvR+JMf7EMwkBPZHc/MQKyzUueD6SLKcBLGsF6dTUrUFAxlkpjNYvnQpzj33HAXI0lqI2TejyUmti+lkAiUFhciPRpCTHUZtTTXKi/OV7VFRUYXs7DyEooWYSPmxfe8BvPLmZoWcn7VyOVbMaxTJfvR4B3JiJahcuByZaEwklUdWkDjgZjKSE8XAyJBIWAPOzTLSe4QCRuLwuZap4IVpBwV8siZhXcCHak82BZGETk3L6olrBmvenp4eERXKqKCiIv1WooL1HclZEgPJqRnZRZKoyM/NU73EeZ/NG1x/uI5a047ZopA8UMCkFFNm28r8KK6Ljoe029mpgbt7O8xaMJKled8na1aOQwMkPIW1ERUEAzOzYdq0mfKICnUT/sVEBa3IwohkW03V3dN9AlFhGRUK02ZGhctLGW9ldpgRFV7zE9d77Sh4L6kg9tp0xF64hh5mAZgX9Rx5YV2hN3z0GjTOq8Pw0Ah2vrlX13TF6qU6picefA4tew7jfR++SkTFkw8/r7nykivPV93Frn3OYUuWL1AWGBUBv/7Z/Vh30VqRGSQqHr3/GV0LdvVTdUHrp7t+/qCUCwzg5rV5c/MurTG0XSJRxS75h+87gah4YSuefeIl1NRV4bobLte4YgYFA1sLivKx8Z3rwWyFX/30Plx+7cVYsWopNj2/Bc8/8Qqu+8AVWLJsPtqOduj7lVeVyDaInvv3/uJBqTNmHxmGSi9R8DRPXMuugzje2iFbJAJ9e5v343d3PqJj33j1BtkOPfybJ3Rez12/Vl3KtBPdsXWXgoU5b7JOZOf3o/f9QTkQF115vu45EhW0ymGQNomiF55+VYqHK991ie63LZu2YWJsQp3YFTXlePX5LQq2vvCydTh7w1qMjVBVsV3XgYoFkifsIi4uKcI5G87Eji278ODdj2s4NC1swLU3XC6i5pc/ukdg53s+co1qopeffhVdHT0oKMyXrZRyHX5wF87dsBbnbzwXI0Oj8oKvqK7AkpVLNB+8+OSrePaxTbj6ho0gUcFciW2vb1d7GzMK1l1yDnZsbsaDdz2ivRo7nS9/z0YcP9ohosJuWN5HVCna3pR2Pjd87L0Kym1+czfuvu0+29/5fLjxY+8VacIO8W1bdmLRSQtw0smL0cbw6u//SvcuCQWGKT90z6PYs2M//vrzHxLxsH1zs5QO7LavqC5XCPa/ff3HuoZXv/9yfcauN/dqfBBkrWmoksri1z8loOzHBz91vT5v66ZtCtPm/UZrKu5/Ca5zvqBVFMkjEkf/+e2fa76gJc+i5Quw5aU3FVi9i0D/Vz6O8upSqTAISjO/hN3qBJS/9dV/l6XUNTdcIUXFfb/4vWqPeYsbjaiYjONfv/wdEePc37O7nuqzu2/7rc4LzzMBUe4xi0oLBdbSJoi5H21H23D6OWs0hgkO/+vffQdFpTF89G9uUm4Aj23Xjn1YuGSelAoH9x/GT7/7C3ziix9Rvsk9t98v73/mjNAWjWPiledf075t7brTFI784N2PoLi0CBddfoHUL7Ts4V562YoluOHm96C7swf/9r9+hA9+7HqNhz888rxew4yW93/0XRgdHsezT7wogHnDZecpt+TJh55V/gj3H57XPfGXz331Ywpxp/qG4fXMseEYJxlN0mnzy29i9doVuP6v+b5jIgJ4r645+1Tdt1R/8HfFZcU4Y91q3aOPPfCk8hDOunAtbvrEB5Tf8vzjr6BhQY3GDtejx+5/Ssfzzvdehkuv2qA586WnXtGaznufSoG7brsPrz63xXAUNgL4fSLQPnbLTQLYX372dSl9SHzUN9bgkd89id/d+bBICBKszKR55cUtUoWtWXsKDh84hm985buYmkriq//6ORGsP/r27VJ8cT/2V39zI84gUfGT32LTc68Lo2ATzddu/YKey98xv4fkJUkl3t8kAgjof+TTN2j8b3llO3bv3If1l67DgiVNeO2lrfjB/75Ndc5XvvE5zUEkTklkszb55Bc/jInxSXzqg18ydw6nDuC9SkD8H7/zRR3/zm17NEdRKXTKmuUYGhrRsbfsOYh//t6XUVNXKQK6o70b511k5+N4ayf+5sNfUfbTP3zrC2iYV4fNm97UmnDuhWtF3Lz64hZ8959/ouyhmz93k9Zoqq0G+4dwwSXniphl9tGdP71vFm+SU4erVcwxIz7bUEwcjntKrzmFTRcC/Gl3K/tzw9kEsCsPy5pxOSa4T/BIAM4NrEeMNDTlrUcGCKNyeKJUGJzbAn48fPccUXHFe801xVunlZPhGoO5n2e9yOsrC3OXO6s9GZthkik1NKiJ19l66neso0mKuCxaObF4JEOAjcpZSNLiymGOBIGMyEnL5pyf61nLm7KETiq0bZ82IkPB1ylhoTpPIp7nbOiJKbLxbraBWi4xtrdifaU8TM/+yVlqsVmE+Km5zCRUi8+pKt5WVPxPwOXf/g5/dAYuqMjTjeZZGHm2Odw8cULgzaJsBnbrMzNBVkqW+aCue09poZvWCAFvcvL8fanHMq86MpMkQOgZH9fvuB/ysi64sBAsp0WJSbOo5JiTfnFT5uU+8CbVxOgkwiyMCMLKYsoB7l5wjiaSGZO5m++hd9yuM5TfSZZLTB01L1sjW4yIYeHPiZsTkGeNZRsaStCsi1aTDyct2rmIGYYmRgJdHlitYz4hjEfWLAoKp2STgGfKvPQ0S7ssiRkqKSIu0yONcHZE70fvewFD6qRIIYuAKW1MgkHJ98w738xlvZBLZg2kZtjJPNcJZ36Ac4sJF1W73gS6LDzbjoe4olkH8O/ssCe4rByGlIUFKZuB6o0AQeOEkRRSUtAmw0gLAn51q1apwCYgze/jgWK0XBK4yDBubt7JTrNTPGJEBb8fJ3UugHwOr3NZaRnaO9oFaHOhampqQkkpVUJps2aZmcFrIiq65VNf19gkuzB22DU0zdNGMi9WKLsnW2QsjJGLKK9NUnI71x3gBbyzY48SxnRSxS/DtKnk4fkmOM8uPxJ1JCKUx0L/RZIVScsLyMtnjoXvLYoK7945dvSIQJ15TU267iaNTGsxIsAvoqK/D7t3NEttMktUNDWiqKxC9yyfywWMgA+Phe89PDyoMMyioiIpKnhM/L4Enjnu+voZUj4si5Ti4lKdO4JNBILVPcDnppI4duQIwtn0pGT3IrBr6yvKzKDdE8kQZln4JKkMCFSPhrJRkpePIpIx8tqcBoNZkzMZTE6ZryQzJNjJQVCmpLQctaWVKMyPaVPOLgwu1ASG2rs6QdCkoqocuQRj5McbQF4sJtuIkfgkKhubkJjOYGIqhbGpFPzZWboPueCTWCCIwevE680gUv5M+WRHd6+IgdHBXvS0H5UChQRry4ED2L/nKE5esQbnrb8YVQ2NUpnwWmaHgwixCzzNsNeUiCyqRggy8T7i9+GY5Bjk+dn62uvYtnUzvvi3X0TT/HnIyi1QPgav0/T0FIL07N+/C3f854+Rppf9dArTDDB2VnF+qimiOUjHJ2XNkpcf0+dSLSBgjHk/tGqTSi0oiTqt3ziHKrMmGTfLO18QU8m0uk2DvgCSibjusWBWAOGAD401FSgrr0Q0rxhXvecDyETyMJFMo7XdKSpOWyNrGikqptM4cPSY7MmYEWCKivXymJeqKDuM4dFRlJYVY1ezKSoaqivgn3FERSAbW/e0yC5ofnUpcjSt0/rJjwNHjqK4sAjFsXyR5rRQ5xyyv+UgVq9cJnUWN728BryfJ6cS2LV7N1566UXs3LkLo6PjpkiSL3pCAekEJzkH05LIxnQamRlOdH6Eso1sZNjt/PnzcfH6DTj1lFM0f8YTU39CVNDShvenCCIqQdhprtwfqKvfs37674iKaUxjsH8SB1uoqJiP2P8HRAVBOYGMDJNOpvHCC09j/4HdmLegAfX18xAI5uHNN/biod8/iaNHj2FychhT8SEkUuOmuJPNH1VkJn02uTTf0Jv/Xde1U/ZpHfQxnN2CfVncE3gdHxuV3ZEvE1LwfHFpBCcvP0lBx7W1ZZg/vwrxiTF0tXVhcGRQXeNsPksmM1iw8CSsWX0WYvlFOHp4F3JzMsjLDWNsPImKykU43tkny7emxnkKf6Xt2+jIEPbs3YHhwT40zluCeU0LRAKzG37r1s26XyPhLLQd3IfyqiysO/d05OWX4vWtL2PBgkUiKjp6gGQ6iaI8P/Y0v4qGxjqcvPJ0dPSNoHnXq8ike3D5JZchMeZHb08czbv3Irc4gIaF85GVUy/rncMHW/D6yy9h97Y3sbd5h9bnUYZOT06Bw5v/F0YjaKqtwaJ5TairzEZJLE+WR7nZIdmxUaUmooIKSy8g2DUycN5jrTETDAOhKILK8gLGJ6ewd98BHDx8GLv2H8auQ62aI+c11GF+Yy1SU7RgasdZZ52hDePQxAiihXkorazQmslrl5WVh1BOE/z+bOREed9xI5Yl0pojKp6Zkh0kLRu5BisLglZP8bjuE9YG3MCPjoxrLeY44lqye9duvPLi8+hqPYCivCC9jjAxNaE5jGsS2yroezw8OoLB4VHVadRyToyNIpaTjeJYDLUV1VizZg36enrRevw4BoYHkQyw3DBlWFlhESrLymQbVV5UjOxAGpPjo6iprkcoOwfRgnLZXO1uOYznXnsR0WgAF56+GjGGUwcDOHSsDeOpaSxZez6ySuqkVPHsrXp7e1XvsAmmb3hQc7YIgaDZCniPEzMq3mL9FAyir3dA54IqQ76GtQYLG55D+nfR7olEBd+3q6tLVoeyEJscRSKdnFVUUMnHmpl+6FkhKpcy6O7ukRozV7lNOVqLWNuw285sWCU+0zpBooKbZv6W4AA30sxJ8vIqpI5IG1DP+rCrZ46oEJihvpk0QgFThVr2mVNUcM7IZNRUwHqQ9qGyflJopHlCS1EhW4O3Kiqy36KoCKhWstw0oLevZ5ao4Nom66fcqGwvzXIKmGgdM5LCWaIF/UHzxCZh65vLCfIAXo+U4N9JzMx6PIvAMMvVGz56tcBhkky19VW63uOjE3j5uS3Y9lqzLvv1H73aiIrfP4c9Ow8og2LV2pMVDs991OGDbaiqKdd1vu0H9+DMdatEVJAYePCeJ3TuaGFz5bs3oL93CHf97AHNu2eceyrOOv80KUe4jhEsrmuoUgj3w799UnkUUik8vxkvPf26rtelV16AU04/Wfch7aCGB0cUui2i4j9/i8uvo7Jhqayfnntik+qEjdeux9LlC1RPs1bp7ekXULl/9yEb1h57BQgs3Hgtsxq6BSzm5LFunsGRA8cUTk3gk4QDLaZ2b98v4JIHwwwZ2kEtO3WpxgLnC1qbLFw6D51t3bj9h065sHoZzr34TBSVFOoeIeC3fcsugbK8XlQ2nH/J2bP/zqYpfs7TDz6nvQbH2JkXnoazLzwDefmWNUPA9LUXtijk+vxLzhUISrCbRAUfDIe+7sbLBdjf4TIiSEowT4Nj74WnXsHwwDAuf7energLgaAP1954paxe5P0+GZe9FkHXV57biqd+/yKuuXGjSK0H73kUzVubVVucvu40XLBxHba/vhO/v/tRNYWdvGY5rnjvRrQf7cBtzCRxVsGeOtZroHvPh65WV/zjD/4Brz632a6Nzm0Y73zfZQIp2e3NvQavx8P3PiGVCM+jiIqGGvz+nkex7bUdApcZ0M2xLcVSW6fsN/nab3zx39Rxz0DxtiPHRWBQKcAxSXutB379MEaHRnX7EGTdeO1FIoLYvf+ft/4cl1y9AWdfeKbAVN7vtMSpbazWnvF7//Qfskc7fd0a2fbwffnvt333F1JxrL/ifCl07Ji6EMlh3UpFxQ8FCF/7gSvN+ul2U2vMX9qE6//KwrS/8XffQSpFVYEfX/3mLVIV/PLH9wist4Bm23PxMX9xoxQj7FTng+A4j5ff/zt//yOpbitrynHN+6/E/CVNaggi0H9g32FZYXUc78Znv3azMlPuuf0BETXcSzD4nWQFiS0+qBBhrsiLT23ChisvwGVXXYTXXzKigvtuZph88OPvk73bN//he/jwJ2/EmevW4InfPyMykvPvzZ//IJafuhSJqSTu/vnvRAytPXc1Hv/9s3jygWedqt81b2aM9HzPTVehaX69cJ3ern6RbSetWITHHngGD95lSp7PfPWvsXLNSXrfO350D958bSdu+KvrsPa81Vo7mPF0sOUIFi2djz88/Cx+84v7pBj/2je/jDVnnqKxxvuTRBDnr8ceeAoP3PWY1kyqfC67+iIUFhfoPJBk5D38+APPWPODspO4PmRp78x57P0fuU7nk8dMJcVLz7yuXBr1jQf9+NjnPiiyjPcR50OqVu76+QOykqJDwVf/9W9QWV2GH936CzRv24/k1BQ+9cUP46zz1+C2H9yN55/aZE2ryOCcC07Dte+/XCoJ7iGOHmpFbl6OxtpnP/I1nHfRWfjwJ9+LA/uOoK6hBrEicyHgnP0f3/kFhgaIN0xj/SXn4Ma/fhcKiwqwgyqte5/Cp//uQ6qXPnHjl0SWKENJwdXW6FnbWImPf/4mEV+8vp0dPRq/VON9++s/RvP2fbjkHefj2us3orKqXOfpyKE2kd38zI9/8Mual/hdb/7MjVi+YpGaYqfiCby2aRt+cOvPNR9x/Tz3gtPx3g++U5k+XGdIQL/03Gbc8eN79TMxCu1PHelpQL2pA1g7E29hXWZq56RlrbrmYNk+0S3lhBB33reyu3KgPP+dWISnaFLjrWuA8KybPJU297mW2WHOLLxOT/5uLvNl47vMbly4BRtZZdduRAHPMT9HykyuY8yAlVOHTZNmDWU5VEpmDbow7hm6IyQNi3Qycu53FC5OvJCNQVJxWmO2rLB8UGMr8w1VO7g6ZtZhhs3easCd1rngmCO+4TmteBjErL2hckKtQdpToQh79XKA6cTBxsIMXQ8sa9YyLoKap1iXCnd1TdhvKypmy/G3f/ifcgbWVxfK8scACQvJZGGvyYJhNc7rnt/XUwx4YYqaKARcE+g2RpY3s5EdnBhYFNgmiTc+FzD+G/9kwc+OeZOOGeDv/WkhOaYOsAnPuqJkBeV+FsvrfP8ErDiPXE6C5i/nZV3MWVVoQyn5mWd/ZJsTTlmSVrlZzZO0ewSHmNuZaQFSUlVQLZJFBtfZE7GTzCkhuNkTeUDCgeCVrBMc+C9lg5edEZwlOAQpOabVDtEIIp5nZUDwNTxGx/qa/IwEj4WX8/MIjPK7GMlin6lJlPkXXMSYKcE2zQCJFNf55oLCFdbknk8lisBjl+MRpH8jj8OdX06+8hZ0uR6UjFLkwkVLm26SCZm0rJ8I0jJAW6oDgv6ppLre12y8DL19/QLeUwSrAwEBgPw7iwAAIABJREFUHxXl5QqX5XO4eTYbMXbWGWOsTbVb9Bg+KfuD4hL09fYiRZuRsRGNCfrVs4uPnRw8d6++/LK6OamoqGuYBz+BtMwMqmuqkBXJRmlFpUBe2bjI45jWOEZUsDtQOQAiG+x+oHJIXdYJC0qOxQowOTFmIEQ0rA5RLkyK0eVYTs+I6KJapKgwpnwELSvqkKWlQq7GExe6lv0tOi9NjY0ur8Rez+MjuTc61ofRoRE0b9shz9uTli5DTn6+MiqKyspECLGYIOjBccDwbG5k2o63IhQKyBqLigqpQlJJ3VOTE+Oyf2J4Lsm+8rJKWX8w6I9AOgOcCe5OTUygq6MdeTlRJKfiAmObt76MPbuaNc7oz0/yROeHxAXDMIMBZPt86oovK44hwnsonUJ8Oi1vcsogBwYGBV5Q2VBbV4/G6jqUxoxQIcnA68DvxY7+zt5OZOeGkR/NA7EHdgzHSkoQzI6gZ3AI1U3zkAlnEZGRP726kAl4KeeB94rJRll4zdly+TA0MiFSYKC/E90dx1BSGJPtz969+7B/TytOWrYSF2/ciMqaGqlxxicndF+FcwjWsyPWigyOT3au0P4rjxkOmLa6fGYG2159HTu3vIHPf+EWNCxcgKxIvqyjJsbHkEpMIjswgzt//mPs3LoZM/FJEQ4aPyJZLciVmRYkP7lhIBBOtYlCnrPDrtgxezoSCSR41PVLQiJE8NgsfUhQ8P7lvcUOE5Jt7D5n9gXtn2K5WVg6fwFnDpy9fgMal56M8XQYR9rbaNaEtatXIRIIygs+lclg36HDSMykZVk22NOPjesvQnFJAQbHxlXQEXwsKyvCju27ZftUX12BAOcLksPBLGzb34JIdg7mVZcjyrmMNnj+gCx3SguLUBKLkQ5F2ufD+FRK6oM1K5ZoXKaQQf/QiObCRx95DI8/8ii6OlrVjcz501NCcS6gsoDnhkQe51mRnkEjr/g/lyLOrQZOBlBfV4/1F67H5ZdfLgCRRC/Pp5dRQWJPRS1D2p2/qWe5VVFWhPLy0tn178/VC5I5+6ZNUdFyBEsXN6GwKPoXWT+ZVYk9SNJIuu28WGVxxrk/7ce2zVuxfeeLKCzPwxlrz0fAH8NrrzTjoYcewZ49exSwnkwRcJ5Q7opIDpdZxPc2AtoIb6qCzIKRm4UM0jMkxvn0NIKZNAqVGRNWd7Zxcxl58tPGjXMBC34Cl8uXLsLpa5YhlRrF0FA/An6qp0gURVFRUYOTTlqJeHwaixefjL6+QTTv3IxUchhnnbkG1ZVVyMkrRl/vEHYfOCJrnEOHjzBeHrG8QkyMD6O76yg6u7pQUlos+6/hoUFE8/JRUV2HsckpdLYeQXfnblxy0Wo01NehuXk/yioaMJPJR28/O5gyykbhnM4NcUVFHWcO7Nv9KlJTR3DBheswlaAyIob+/lEcPboHU6kJLFm+BrFYuQKZn3nqGfzqjjvQ13lcypLRKWdb6AeqS/KxtKkWjZXVKMrPRW6eTyRFfjiijAp2ixNU1novVadZzKkBQiRS0IID/dkIZOWaGk+WS5Noaz2O3Xv3oHnvIby+6yDG45NoaqzBqUsXA4k4Bkb6sGLVCqxafSb2tnbhtW3b4csksXReBeY3lAk4SKbDyIrEUFrWgOxoGRAowPjEjBRdk9P9al4oKa7A+GgCqSladY3ps8O5tO2jRWIKwyMjIpF4nAQdDh44iBeefQb+6ThS4/3ICfnQ09uJUJhNEX4RvPHkhJoeEokMEvEUKsoLMTbYh8vOXoOGhkYMDIwimBWRXdTRtmNS2fkDac11uZEwKsrLUByjqiKqeY12f8xeqK6pRV6sGKFoPqZ9IRxpbcezL7+AqspSnHvqSsyMDsFP28X+fnT092H5OesRqZoHX5D3OusOU/axViVw1tvfr827p6hQdpdrhqEyhGuMzSuhWXsDXsvBkREMDg6qxggFA4iyrlHAdMJ8zAcGpJKgGo9ZR0ODg1qrx0hUzMwRFZ71ExWCzLpiPdHd3YfO9k5EQ2HZblCFR6Cc9Y8ajPw+Ox6pPQysYY2utYWkBBUWxqeriUL6Ardx7+s16yc2KLDWdN6hAkKk6lXGhHUAsh4iydTe0WGBnNFsAYC8RnwhCW3WVrK9koWT1aKcp7Oyo8q6YUaFlIDKasnSvw0O9Gucs4bRuhX0K5eGndpkGfj9xo+Oq+nA1JJBU5DoT7JZat6dPXZLh2Gxbbalxu26Tk5nDWpNQ6xszDJGWXCacK3O9hLrvKYq7gesNqZa2+p1ebFT1vZnH2ZHpe5iNTCZtaqEHTooL6TBFNB2hEYkez7bGnday9lpasfmPdtAJF5QwVBvOQKeH34n2XB4gaTKa5rFyWdt/vS2bi2leoJEBe2aHr7nceczb+fFs4DVp9lWS+9xopLFA6U4Bq1Rxmp8d+jeiuYWtlmBi52IE8kkF9DtfSlv38MnUXVPy1oRWK5zm/s7z07YzsUJyhq+e9rmW+9cel3BvD5/+mDzGp+b0r6QAOLI0DDCEVr7csxxb2g5iD4fvcXjCLPuZSYYa3Pl8zEjzRShXEtNpuhUPnY2BKxxD2TbUttL2Ll1fiH2N3eu3T7XhdOb+tHAuNnXzQ2oue/vMojs+daExjnhtHOYGXGpLLLuv/Mx2x/KP92y75SD6AYaD4/3HOcTjjmuRbIigRG9nCe8pkHWot6D487e98Th6TMrNwbJOpWy1wRnWYauc9t1qSvLQmOTtcq0CFeSYoYbBK3z2B2TXAb4cT77XDtOu7/ND97Old9nOY+8Ph7+wN00975yeqBdqBwizDnCfPLNFkcW05xoOKG4oSPAUjgH83WsLufzrSOa+1hrcOSe1ObFICYmxrWGaO85i6XMNY5w7yFgkjUwm0TlGmG5D7LdYW6Yy9vUWBKhbGPEc5Pgz4bRZExtohxLsyMkMMpjvub6y6QQ+8Mjz+E3d9yP9uMdqK9vxNRUSopLfjZBX9aRxEdow2h74pj2kDwWfTabXVwAsXdP8VitsdUwBs7vwoZcroMwIGdPrQZUqact24skuVwVuNcU9mF2Pt5ax3HPccfvJetD2pbTKYSgscOfmGXEfZWuu7v+3BPwYpy3YS1u/swNUp794Nu3ay5RTcEMTzdczbqZOQNmK8TzzX083R14LnmsU1K7hzQGtU9j8yEnCaoRaIfEcTidxr9+70uora/Ed//lZ9j+5h43pgw81xyqLn5rmuR3JJHkjUOzDLL3M1cOe0/hQm5tJf7jqW6IaXg5DFwvFUTN3FN3T81auVNB616n+9q5e3hzOM8bGyE49vidOF75Ha0JwYKrbUwb8E8S0Rw/mEnBgG7Lq5hdK0RUGNbHMcqx8dTv5sLgL7nWmvY8RYewGL6vu5+4wHvWUZ41rWdj69lKaS4RpsN5k/esjUGOJzbJsmHPax62ddbwwlmck3ZXmu+syViqdafs8MgNfTd3Tji9cY7XntKt7byW3jn0lniOLe9ceTZSdmzW8MwBqjnaXX++J0+0rOkZAG4yd7Oletv66b+ot97+9f+xZ+C88vxZn1hOdLzR1QVMS4sIu5mMqVQx6xQQtCnijcXCfK74s9BNj4H07IQI4vAmlYVT2p7PRZCbKE64mrg0uTkVg1M+SIrFBYa/V3HCbiyzpuKkYRsidtyzq9r8ZnnMfI2CTWkH4iZwPkfSby6I0zPqmOTEZQuYqTJMKaAqTQuR/l2TM1UWtpPhlEW5F31wbaNHuyuzyuKiwcWJwD0LHRZQnHh4TFpE5OscFAjN11iQr8m8eH75BQj0cpHgxGOFT0byfSokuDDpOzMgSOQEN2AmI5P6woXwcCCym1Ud+m7jZfZUNKun3N8suvQ87kxnN0O2WfQ63ax6tLBxvtY2XQwY57V30j8BWWajw3PB9+bfaeGl7iZ2SSbjAnKVUZFKaDE477p3q8hQIHZfvzofeA2i0TAKimMWysSAW+eRbufVrhMXToLMBGv5KC0qlp8zO3ODQTvX7Hasq6sTYM8CZ9OLL2Cwtxc1dfWoq58Pdqaz2GE3TTozjcLiEuTmm40CC4msUFjHxwWcXZVmz2CqCA+4Y15CMjGljSntCQqLiuTdTEsekjZZ2RGEo9YNIKA9kVAXPnMVQOspjlAuTskU8gjIS56YxI4dO9SZWlNdPft5CqrKCqmojU8NY6C3D81v7kA4mI2TTlqG3PwC1DU1Ir+oSN3+5uGZFshBRQULwP4BBggPqlOcBACvKY+Lz+XvWRiz8OQx0GaK50KZELy2pCEyM5gYHUFfbw8Kc3MwNjqC2qpK9HYcxvPPPmPFIjf2mQzycqz7inVAfg5BIyAaCqKksADlJcXyWk/4MohPJdUJ3d1D25k0SkvK0DRvHqqKypDHUNBI2LAEZBSS3N7VoXuXNishfwi50VwEfVkoq6pC//Awjh3vxIJlJyOnogShSETnRxkt6RmMJwnG2yaA15Egk0Bst6GaSqSRSsTR1d2GjrYjykAYGhjAzh3NOLC/HcuWrcSll7HDpQqpTFph8ry+tDaaSqQErEg9k0iJRCAgVVRcqE1zypeGfyaD3Vu24Y1XX8fnbvks6hctQna0QEoodg0jncBgdzv+43vfwmBvFzJJ2pwZIekVqySR+BgaHtX5LSsrk5UIryPBd5tLk5ojOZ48AsOAM1r7mYpABfY0i+os2wiJaKG3JYPFfFI7rDnpJBTk5SNWUYFzLnkHMtmlONDeirQvjbWnnIoIlSx5RlTsP3wU8XQKx463YbinH5dfdIn804cmxjX2RkbHUF5ehO3bSFSUOaIirU1jOhjC9pZ9CIeYUVGJMItrfwbpAHDgYBvKC4tQGivENBJI+4GxqWkcaDmK01YskcHRtN+HPfta8Lvf3o/nnn0Oo4NDyExbeLypZUz9ROJzeNgIJPmX85zMAnf2dy+k1ebphDqUSCKuX78e11xzNSqrKmwzlSTZ7NNGjEW/iArlDbB7NyTwq6KsGBUVJSCbdiKpcGKhcCJRcajlCBYvbkLRX0hUWAewPZi5w3nX3P2pmLGt1KF9h/HaS08jGJrA6rPWICevBhPjPvzkR7dj8+YtmJgcNaIiOSl1GB9GUDtwjnO6y3by1gaSg7KLkTIxhVBWBtFwENUlxWioq0dJaZk0A8EQibMsHGttw94D+zHEvCCeGx9QHItixckLUFkeU2AsibOc3BjOO38DqirrMTA4hrGxKXX0cw3Yu2c7xscHUFNdhlNXrEBlZSX8/jD2HW7D8PiwrOOSiQC62vvQ3dGKquoi5BVF8dzTfxACtWjhAsxfuATTCGJsMiHwe8urj+GSi04VOdTW2o9QmGRnATq7SU74UV5RKbsjBg7n5xUJWNrf/DJ8qXacc/6ZOHD0ONLTUZEpgwPd2L93u5Rpy1ecDl8gFw/c/wge/f1D6O/qQHbIj4GxMeXAlBREsPqkJixurENxTh4obM+OBpCbE0FeOIJoNv31HbAqayDaLgYREABLVsjsgvzctAeogmLGT0gZOQw7J2C2Z+8ebN2+B6/s2I+e4UHUVZfjrFNWsHUfI6ODqF+8AJduvAb+gmo0H2hF87YtaG15E/lR4OSVS3VdaEkXzM5FXqwCubFqZHyc00OYIjiXZk5QBeKTVCrRbo3jaAKR3ByniOG9ZkQF77+RYZvj+3u6seuN13GgeQtqyoswNNSLvoE+3UO5OVFkfFT3sQ6KYmoyibxIACX5WXjfZRtQU12D7p5htPf0I+3zy2Kyf6gfifio5vXsrCByI1H9z057Zt5MTXJDH0VZZRVixaVAVgS+ULbWkuc3bZLl3YLKCsRCfuSQUJkYw7GuDsxbdQZyahfBH4ogPc2GEZ+If9aV4Wi2iArWB96ceyJRwWBvb25hnUfQR9eLAdmjw+gfGLCw65AFXrNeFlGBDAYGBxDLL5CigiQFLcu4Vsv66QSigoHSWr/8tJ2LIBSKoKe7H53tXYiEwiiIETBl3hzzJNhQkdAxnKjwMGCPjRjsziPpSADLABvlb8v7yR79JCqYXxemlZXZ7LG+5jrjAcECpBxoRPCFRAU31jwGZltIUcHQcBIVk5bbZISDAWwiKrIMxOnr61cTBtcsgk2swwf6+04gKkxJTKUGiQqCDrw2o0fG9XzLp2B9b/Z3XJvZLMD34/vLps91uApwJC0ja7s5ssBAds8aynByr5FJtbbLZ5u1vmMjFUFOBxTz+3mNUR4o8aebRKfc8MBo1yhlvtYGPnkgvxTFsnS0zA3VVw4MEgjompQsj8Rqdlvr+XdTTPNcm1UXa3+C3l4zl2EcnNelsM4Y8Cowl+/hHVcgYNZP15GoaMEDv3pE7I/ZWZg1Ld+TwA/fyxT1No68c6tahvstB6LNHaOFQKvac0PP64a182fHqvdSOK19nnFptlfxyAcqvtQkJvske6514jqAmddeTXZm28aaV1leslkyC1zekwInXdONnQvbB/EwqO7mHq8glqcmPXrS8x7KpLnPI0jpE5mRyZD45lyRrXuouKIcY4NDGKMiKxLVUet9BY5bzpM6f2Wlm9Be0SMAjNQyYk3gWijLXSOzbPNCWA08s2spMNM1u/H13M8JwHZOBQQKqaQYHRm1QHtXH9N+6Job34GdW/fgvjsedk4EBMItAFbNgALeA7ovmZ1oZIeNAbseBlZqjLC5QfmWnN8dSUZKn2t3MjFLaJB04MtMkU5r0ozlYfK+dQAoryWvGfEKfpTZUVv2HO8dku2yvHOECm2ReZ2piuX8oD1siEAjm8AMqLbxxMYms6eRkwQtcOJxcw5whKJAZmGvNuYEpAskNqCar9F978+IJOGx8NqS2OZx81hoT2qd4DJq1e/oNMC1wiMgNZ/6LSNAyINrLPL2bbm5ecrn0950etr2ulxLUpynw9pn873oWuB9nvnz273AZhuOT84pxGa4Z+XvrMYwlR9/vu6Gy7DxnRfgyYefwwN3PYLDh4+gqXE+ksRigtlI0KWBezKnKM5Mu3uE+BAts6U4tLrUVLnW0MYfeaw8VcqcnJrSmj0+YdajutZBI4p4jBwDyhRwYDm/A7+LSAIRyeaYIbscl59ENSePbfY8TIw7dwtTQXtEmtfwKpBXZHEA6y44DR//3I14+fmt+N43b9Nw1pzo5jbNk1oe7PmmnLcgZM6XcstgTa7GxiyNB1mrs4GMhHCIJIdZD3Fv8u3vf1lExTe//hPs3LbfrYdGuBFz0jnR7ZTRdfbskzje+O9aw1w4OY+Dc4ZHTPAo1UBMa3aRiUZ28D4mUUFlBesaficSfZbdYIoFzhdq1nR7ZctVsKxa/k5rksuTlSKPDgiu3rD5jHO9YWl8rhoT2BTh5b26OVgkyImEJesQZPDM/XNExcXXuZw03sdUFDscTHMBj5N7Eq7nTjmh/Fc1+/IzzVpd4L9rKvbWIo4fUz2QqDDMyJo4jAgQoc6mi+yI8D2+zpqHGQgesSZv5zDjzc+em4zhICQDbe0ib8P34DFxLuJn2hrLDA9rgtb8wZ5iR5Lzs2VRrEY6s6YyPNHeg7iSMDr3ureJij+ttN7+zf/hZ+DMInaX2k1kLL9Jq7jAcuHXZkMSd7LsBJ85ybjAbBeqqQmXN6MkSgl1f88G0rhuffNbs9dJdRBwvnEC3K0jQ8WTik8r0r2Him4uRFpcraPKs6PQwuDVqm5z4BWwLNBYjHIiI7NOcoXfS+/lZGseiK/v7opGLuBSQvA4POVGkMUjpALh9/M6QazwN9WIxyjz36yJybp4JNVyBaFCCBleSMKB55mbKgJmLEyV22FFlhe248kcPXneHDlhkyt/L8LIeQRqwye7HismeVwiXLjAZqa1UAmgdOyuLb5aFWYf1gtjmz8+ja/XhlR2AcYum4SSBQ2DgbgBZCfytAgh+eqxM5lBzBPjsn7i59K2hVkV6665zt4vPYNO5g6MjCAajshKYjI+LoA7GslDJErAgQGSDOk0SwF245H1ZgHpm5mRomKwfwDxyTF191ZWVogA6ejokHqAYO6Lzz2Hwd5u1NTWo7ZhAfz0MfVnMH/hPPnST6VmZD9BqyKqNxjuTABfGxh1GdGqbMrslCbGrSBmCHdBvry11dmhwCgWun51XzIUMiZLKZMT8zl8xAqLNC5IgGiz64gKXrOe7m7s3rMHdXW1KC0pnbWMUudAyIiKVGoMvV3d2PHGdkSywli27GSRLMzeiJWVoq+/X58jOw12JCoLJEvfpbXtKGpqqlFZWaVj4u8ou+VGiyBuLFaksdHT3acChuOHoISC2AGMDPRjcmxY4a493V1YMK8RQX8ajz3yCHo6uzDD7hKfXyGomk9CPuSwo98PZPl9yItGpMKQ9RRl0Q60YVYJbWpolURVRWFOgQgGjk2OpcGhIfT092N0fAyTUxNSwfA4s0Nh5OYUwBfKwpHWNnXKrn/HFSisrUYgnIWsQBYiwWyB6RyDYA6Em49IBnlkH0c7vfG5+eztPY7OtiOor6sWUNS8cxda9h3DSUtXYOM7LkNldRXS3JSok4jAvnWQ88HODpI19Atnd2xpSTH6B/uRmEkJ9D+8ax9e3/QqbvnbL6BmwQJEcvORnRXBxOgo0skJvPbCM3j8gfuQmhwT0KTx50AJHis3I5yPunp6wI2K17XE+doLaE2mSJ5RCmrzJ6+/7Do0D3E+MwCF15/XQQQjQQt5iwOhSAAzyTgWVtdg2eKliGfSOP/SyxGrXIj97a2YzsxgzYqViPh4vYyo2NNyEITa2jrbMdIzgMvWX4TCwgKMJae0mR6hoqK8GDu370ZtBYmKSqeoIFERxI6W/cgORTG/uuqPiIpWlBcWozRWgGmkTiAqjuG0lUs1H3f09eH73/8h/vCHZ5CYTMjqBTPJWds+gTMq6Kyw5bxHYlObGucl782p9F3nzzx/3IRR5cV7nZvws88+Ex/68E2or6+XVJ6boFmiIiukDaefqhSSkDNpVJYVo7KqjHT2/+9EBVcfdrAzi4NqruKyEvT19eK5p5/A+FAXzjnvNDQtWI5jbZN4+KFn8PijDwqwTiY5p3GeizsFI4t9O0feuNOmz1kmsBtaG2l28PkIOKSRn5eN5UsX4qxTV6G2uhqlZeUCHKM5uZpnOzq7sXVnM17d8gZ272tBXKR7ECtXLsbyZfNRWBxDY9N81Nc1IRzJk3KhuroBscIStLa2Y8uWNxCNhHD22tXoaD+KxOQkFi1YiKKSUgwMx7H3wD4sWroMw0NTGBmKo6+7A/7AFIrK83HvPfdgOkU7kBk0zl+A2oZ5RurEJ/Dys/djw/qVWHnyYowOJ5FMRxErqcbBIx2YjKdRXFwmq7FkYhq5eZwXQ9iz4yVgugcXbjgfQ+MpHDnch5HhOFavPhnp6THs27sdk5PsJqzAXb+6D7t37Mb4yJC6UMemaJXnx/y6MqxetgC1ZaWIRXOQzdyZvBAiWQzNzpJ9njVpGADo1WT+kOUdSDVDxSvrphD9+Xmefdr08nqS9Kd14KYtO/D4C6+js68PdbXlWHvyMvhTKUxMjaG0uhIXb7wWBdUnob3fNjl9nUfwxuZN2LNvFxqqw5i3oBoV1YXIzYsgGAgjHC5CcXEDRlJRTGeyUFRUonNDG4/x+KgUFbl5+VrXuE4ODY3K+onqRIZpd3Z2SeEw3NOO5s0vITgTR+uxQ1ori4oKkcuMKN7jzBqaSCOIINLJcaxZOR8XrV2N0uIy5Wi8uXO38ogC7p7jui87TTZVsMGE9U8wqPl2YHAENfV1yI7mIppXgKzcfJEPI+OTeHnz6yjKy4UvPoG2PbtRXVaKgpIiTPuB/Pr5yK9fAn+IhD3Vpn6tVUSjqAjqH6ICkBlFRg579wvP4/8dUdHT26vNMAkVqgW4ZrA2ZH1EooJh2KwZWBP19vRoLR1nmPYJRAUtwURa+wgKkRgJo693UD7nJOcLaVORSsjqkHWcbeTZvc35ydaCPyEq0swAsvgyj6gQkS+iolt1PYOtBRarJiBIaSSDB36Z37MpX2n9xL2DZVREVdfyhVTW/jmigsAuaw7ON6oLglmaswlI8MH8jTlFhREVfF+CrBwLPKaxIyNvyafQfeTU4eyw5/F5XbVeXW6hnwagabNPb2jX6epExn+ywzOiwrrdzUrGFBZGF/zp48/9zlAL19Hs80iUtABCIxoIoFrgJx9eQ4GBY0ZUqJv4BDJDgImzuBGAR1DaXXs1VTkbT67z9rw5FblXL4hkoJWs91wRItbgxceppy/HO959sYgKKioE4HJPqE5VktyeWsFUOhp3AnusRvL2jm/dbbhmUAe2ecSVt4/TfsrZiXrKem2vPED8jwgO7lFmYOu7QCURPFSJG8Bj3dVW83iECcetAcUGThlYbR3PBIKsQ5sWhkYuss6PT01gMj4hpTOvD9csP0je2d7W/MwJyE6ayj6ZQmlpqfY55s9uAc8WYGvHqmvi1l8SmdYZb9l2dm6ta99rZtO34d7DZcWwlvdsf0kIeMG3UkO4fb5IDGU8cg9mzX38TiJOZmak0j3r/NNx9Q2XYdvmZvzmZ793JEhGqmN186tr2MBYfleeD2OO3JV1XAW/jwekKpPHA99mzBJXWANzb5yaiOdDgCNr1whz4qzpyptnvWw9XiPOk1Sxy4bFNeypWUc5hoZByDKUC7nGCkFLlzVJ0lT5Y3DZgnZPeNecDgJ8T8uz417Xp+vGmpn1kBeMO2v34hoWLYuTZC7Bywwmxsc1r7B253fk53PvQaWp1znuAdbcQ3Mc0IOepA5zF6RKk/Wx5XOSViV2YOo1UwdLEe2wAH6G51zBvR3xAz5sDfAcGMySOqRMO9qrjetn79iJQ3D/xXNz7fWX4vJr1+PxB57Gb+98CAcPHBJRQfKeKm2BpyKv3HzoOrvnSE6/5ilZ+bgOce+29RogeT55fLKc1nbT2fiIvDaswlNfCTw/IU/A3CUM5+H4YkaJ5k9hN2ysNEJT1ssJNh7lmKUzm2edKsEaU41U1dGqAAAgAElEQVTg0DyQlSWi4pOfu1E2ST/4zp2qr7RfdwA9MRsSbMK1REYQvwoKn+CxmmrbhSuT/CKe4NwOeB44p/B7mH028L+/+7eorq3Arf/yM7y5dY/GomP9dD50fG588vnCbE6wNOd54prhKQC0pjnHE76PN4fYfMw5isSa1QVS/NDhRMSCy9lzxJy6/6WGMVW/jWFTVXrrpVRhtI5kE4sIcVuPtd8Urkg1iGFJ1uBk5IVHGrAfQHOf8bQ2BtzPz95v54eP86+ccGolW9c4n7OBVw2SqkuoWjEi1cgrXnvOwYbheCo5I9Mte1WuHSIlQyL0zL43oDnO5kkjp7jf53N43Ty1igK5mRtBkoquMRy/DBt3Y8QjMTk+vOYDKTMcufiW2snN3/yepogy1ZfqETqnyFnBNWJzTXPEhJSwUlzZuqaGhbcVFXPlxds//c84A2uLbAHlw2Nk+bMYPikguADwhjYGUeA0pWIqAmyz4k2C3hlhUcZJz/IEnHzNTXZe8W0dQbzRrYYwhZjJm1TYqlA3gbWe6xUyJzbQuOOUDFXd/27T6CZR66DxQkWt4PaYTm3UXAgQP0usvzqqbBOkhUIMtfvZb11AnBh0rjQZWTeDNgBi1m2C1MMtLvzRY/u5+Etu7SyZvO58A09N6mabP5vgef64GRaxwgl4VhY3bUxqIjErRZXknMWAY5C94l4SRDeZ8ZisqLAAIW12XOHoSdzdMjH7B0N+Jd1114ATNjfYXoeUCnplD1gHFzu61WXBwoAhzCyqCbrS9illf1JRoU09F/uphAB6SiSLi4oE0BJkGx+bdItiSF3N/D8UyZalFDfp8fEJne/SkhIMEEAfH0Mw5BM5IV/Onl60tbXp73uamzE80Iea2gbUN8wngi5p+KIlC7WIJrkIpzNSO+TnxxTybYoKqlfsPLETmwWhAN68fPOXlrSZHt0TAvIJMtEXlWBaT3+f1DDsbuHixoI3JxqV5zQVuJ4kk50NLJ5yozmyYjl+vB2LFi1CQUFMi7HIAhfyTVBxfGIAxw4fwf5de1GYF3uLoiIky6dBVNfUCGz1CiYL6p5GZ1e7ztmyZct0D0sxMjMjn8Ourk6Ul7NjPKxO4q6ubgsDldWDbQmH+roRHxuGn12PPd1YveoU+Sc/98yzOLBvP0YGh/TFSC7R6iE7al0w4VBQAafZoYDUJ1yoGVDFLmUW/pRgCkzODuvaRoNhbTRkE5eexsjYmIoEddEO9CMuADwbBYXFyApHpcx48eVNyCssxkVXXI1CWnpFIwj5g4gEwmb9NBUHZhICsThWPbstr4Omr39Qqpy+/k4pKhocUbGLRMX+Viw7aQUukfVTtQpT3kvyjBTBFtdmlaBdrCAfR48cVqg2iyEeb3F5mUDv/dua8eZrb+DzX/oiKhoMQGM3E8dLYmwUD/7mTuzf8SbGBvtVOHIzpPvYFWQe0NDV3SsiitfHC4zneeNzkymGa4WtQ41kDs+3N3eqW8NAaI5jKm543r3PkcVYThghP5Dj9+OCtWcj7Z/BguUnY9Gqddh/vB3JTAarl69ENgkpEhW+NFoOtWJyZhptHccx3N2Hy9ZfLKukOOXAoaCIivLyEuzcsQs15eWorypHIMNNgQ/TgSB2trQgOxSZJSrYfTTtz0hRUVZERUUMaVo/+X1SVLQcaMXqFYvR1dWDO35xB5548in5uRMQleIswfNm8zS/H8+BByZmO0sWKl7UneI28CKFAkbs2OY5jJyozTs8rwycv/DCC3DzzTcjP69AxCmJCv4ZyvbUa1zPOLdOo7KsRESFa7/7s8WCp6gYdtZPS/4fWD/9saKC8zJDizmO29qP48jhfUhMDeLUU5agpKwUo6PsFMzDt7/17zh2rFk5UCywE0kCAewesk4dX2bOc9/bbOrgSdaSnPNlwNkzNxLEvLoqnLZqOebX16KMOTSxAhQVlyEnN1/5LwRgSOKNJlI42tGF+x54BH944UVMZ1JoaKzChz90PdatOxd5eYUYn4yjvKIaZSVVmKECMkNCqR8vvPAiqirLseqUk0Ebwu1vbFH3fVNjE5JpH1oOt2D5ilPR2zuOgb5x9PV1YXCwA0fbDiG/IA8nn7wcra2t2LN7L3LyclFbU4vC3Aief/p3OOvMeTjztFOQTIYwmchCfmEl9h86grbjncgrKEY4uwDBULYIZ957e5s3Ics3grPWrUP/MIkBesf7ceToPjTUFqEgNyQf+V3NLXjqiWcVCMr1eHxiFGnfDArzo1izbD7m11aiJD8Xsdw8y4YJB5EVpCVPQPMkASALzGaHq9lC+mRnQwKDACQl/kEEw7TGy9H2hONe6pipKa1TW7ftw90PPYHWrg4pKk5bdhJ8yQQm4mPIKczF5Vdeh6KGU9AxzI1VAD7Nx34FXL/0zIPo7W5BWUUQTU2VqCwvQyTI/IkczOQWIZCdh8JYORJJbnL9mBhPIj6ZQE4sqnXViAoqKuZLZcr7squ7T4HVh3Ztw5G92xFMj6G/pxNpqnKoXmVdOR2X9VM0HENuJBf93W248PzTsGZJEwrzC0XMUG2zY/ce5BUUSF1HclnzMIMbuQGmdYbfJ6vF/IIilFdXIb+wGDP+IHxZYYQiOUilMzjSehwBbuQTcRxq3on+brMUbFi8ELk185BXuwiBYATwEUwMiNxkRx47cQdHhjRnnqioEHBNMFj5IabWknJW5IApKvg6KktIKudHc62DkYAmu0unLSeKRAVBLa4fbAbgujExNY7kTErjl3M7N/y0m+RUbjVuFvr7h9HT1SulBsm/TJpqJ+ZFWb3O47OuVBfELkWwy6kSmEuigh3TBCAM1PPmzMG+btUiDCFV7StMwAALrw4UoeZsnFgHMkOEVhVUVJBQIPjGGXkq6YgKBxJ7ZAdrKVoP8rUD/QN6PutlWcVkMrL3ZMMF1xMjmANS4EaZ06GO4AxGjw0gm9eYzT8BUxV6YIKs+QS4m0Wp1kFH2lu5Ppd/p74dBxrbF35LVWxN4rLicEpjB/DMFf9/2d5Q2xYPzFKHrrNZJTAnkImAhamWZ7vknXWOfucIFV4L7R0EwtpeyPs3DgAjJLg3MrDGGl3nfm9Ha1/SCCzbI3iKcu1HZjvOrX5SN7NAYbO0UDPs7ObHqRmclYjZ2hpJYD1Rc9TN7Evch3tdruqTcv7nPM+eDQx/5405jVLu2f7odJv2nc1wTjlOooIgklRDZqWqa+4Iu7m9qu1reHja67r8Qc/WTMA694QC+Ln/MzUlSUs205SWlGuuIHCq8kOAHDe302q+IujORgLumZjXwKo6KD9zAyXtmjgbOQdUznWH21iw+5cd+mafJksr7Uutc5ggmTcXcY/unSuv2Wyuo34ug9K+rSns+V2lYHDgvvf5XoOPMiLdmKKVqABOz77pxOvgiAred6YYMfWyWZdxfTe7JtYHngWcLFc8VY5UXtZ5zO/IeUBZPqA/fFjqFH6u8viY5ebIDdbT3GNKieCcDDj2rYnQwE3uSfkduIfQ+XTjU5Y0dhdYl7jDBQSuuk5725fbeyt30wHsUp7y2LLDyo/U93R2ewJJqXbgdU8k1ZDF6+/NmWYXZR36HrFmwCjJXSP7lN3p8i75Or4PL5r3ey+zU6QTu+FnZjSH8rx4ewGzOfKUGpYX6jk9eESAZwEkYN6RcxlwrhG8i8NHjqCutlENCbJLIvnERokZs6nlemNWVmZZzWvv3e0iyHlvqJHTuvSlBHbKBKlGpCI1VQJVFprrlW9qa5jmXfMjmH1fzWdyfQgom0EWVGoCtY51j4Sdtc7mZ7r7U//mmjv5Grn0urnNI1/NytzOHe9dnlceizfG2DHv4WXenkPziwBpz65tzrJNWZVZXIvt3rE62zAeD0vS/sXlneqakLhyThsecePtXWZf52oQTwVGIoXkoylNSJ5ak6qHvXmEt+ZapwDRnOWtMVLlzeVXGIhv592zI+fvPBKH35kAv3L/XE6eTetGdnACVlaDm2M863QvH/ePFRV83XMPzBEV511Jm1rmZORo78LvZfOSjTBTq5iTh4hdrXuO2Od9T9USlfPOEs5QDXuukRBmyabfK5OXfzdFrNeMwAZnWeM7YoHHYRZtbi2UVZldc2/u4uGRxDG1FxX5xMfs73actqZ56hQdk5eLquxbW8fkPCOLbVotOhySuJsjl3gjEXN4m6j4y+qvt5/1f9AZWFuU6ySqFj5jFkdOescNspOPWmFhi4zXYckbX4vCtE22XES8HAvzCjQfOgK+JtO04s8yHMzHVWQAW65NTz5rNyT21iMqnD8s/1WTkifDntP+2kSirnZb8Pm++gxHphhwb4ujt1ER+0v/t9mNiifQOuFP162iicV1T3kbFYH9UliY1yGLV6kN5DdnC5vXuauNnbogbJEkkKsOKHozMriHQdru+ExKbQuXMeW2afSKGBW46hC2c8gJlu/nbQZ4XNY9bD6NKlwkQfNLYmqqFEomTQVgi4g3bVuhZifZNi1il7XwZ2shkDzY+W6a36MRS/JDnknJZ1ie2ezWlZJiynInSGKkklJUqOBk5/d0WiQFrQ4Y0EyvaZMWpzEyOioAhEUd3y87J6zCiISGrlkGqKqoQm9vD8bGR7Uxr66p1kLE4yK4QLKivfUYpqfiqK1vRF3DfPj8IV2fxSct1DnKzskRGM5u6PLySoED9LQnWTE2NqHz5zHqvB6eZQ7PN4E+Wk0RXCKARoCW52psbATjk+MqQKjOyMsl6Gld/LTVME9MAypoocNN1NatWzWOaJlBAN9TPfBPghcTk+Po7DiK462t6DzWLpuIxYuXIDevALUN9fCxKyYYlIrEK2JIPFi2yrTzMG/FipUr9R1kR5VIoL+/T9ZPNTV1boMaEGHC75+bl2v3TWYaw33dGBnsw/hQP5LxSZxx2mkoqahQUOobW7ZgsH8QE7I48cm3NyvMbk8/ouGwQsZz2GUykxF4z8KyrLxMpBDvIRWA4QgKC4vVxUCigmA8N6iyRmNIazIpwEJ+qjm5yI0VytojnkzhN7/5LZrmL8LFV16NotoqBEgS0R4qK4rE9DTGE5MIzNqe+QT4GNlkj+HRMYyPDWN4uBeth1vQ2FArn/Dmnc1o2XsMy5evxPqLNqBx/jyRFFRoWNeODyPDI8ik04hGskH+tu3YUQWbcn4pjBUiEA2LiN35+pto2b0PN3/y0yioKMVMICAiK5uhWMNDuPeXP8dQZxsmhgYwE6LsfEqFIj/HA8V4rFR/8Nxw/vA2IbyXzKKPWTqm+OJ8xaKa1ZrmLvIrTk7OsUfAjK9j9y43QZwLQ1GSa9mYHh3HhrPORnFxPqLFxVh9/jtwoLMHqZkMTj35VEQCIURysjATAg4cOi5rreNdnRjs7MYVF1+qc5RW4Gmurjf945ubd0lRwZwKZhpQRcPt+p7DBxD0h7GgpgaREG06Mkj5Mjh4qA2lBUUoLSrEjKyfMhhLkMBoRV1NKe6957d45KGHRbJxDuF5YiE7I0LRCO8/7vplxzNJnfGxcYGyHlmszajfLPVYTJJE40aRc4GF07MjKoGrrroK73n3e0VoMluFcznHuWfb4AO7MqdRU1WOcoZCmnHa7Djzumhspcsok4cd/QzTXrq0CbFYxFlZ2Lr0Xz3e8p4izE3mzHtj06aXsGf3VixeWovSshL4fXk4dnQMjz/xMrZtewPxqT5133Nu5xrOm0udadyk0HJPKkKzVrTVwGXtzKQQ8mdQUVKAVScvwcqTFot0KszLQ242FSj5mosCQd5XXIe5oAcQT01jIpHC5jd34Yc/vwNHjh9VUOXnbvkUrrj8CoyOToiYqKtrQDCLjRMBTEzGsbN5Fzo721GkkORSNNbXw5dJY9NLz6OhvlZjd2/LHiw7ZTWmpoLo7R1D+/FjaN61BXWNDVi0ZImOnxtKdqcfbNkvQrGuqhwH9r6KxYsKcf66tcjOKsTohB/DYwm21qFvYBDH23oRCESRm1eI8ooK5ORk4ciB7YiE4jj9zLMxOAJMTkUQiRZibLwPA32tiAQziOUW4Oknn8NDDz6E7u5efX48QS9loKm2AqtPWoj8rAD8M7bJ0vgL2HzEvxcVFKC00HIW8nNof8d6Qp51VgNwi84aQ0RwDL4gu/p9Wkfi8XGFMnKs7m45hrseeAyH2o5hflMdTlm4AOmJCeVAICuDq991LSoWnIHWQUJ6YfjYIJIVRElpBabHJrB1y/M4cmgrhgePoygWxbzaeSgm4J+XRjBMe6EK+JAPHwoQnyDZOYNIQRbSPiPXCTbPn79INoojI8Po6u5HbjiKTU8/ho5Du1GSG0IiPoxp5qLws5kyEg4gO0LiJYzpeBLDA11Yt24VFtVVobSoDFnhPExNpdHd24+9LS0K9WY9wJJOaWjptLKTphMJ1FRVoaq+DtH8fGRHc5DxhzDtDyIrmot0xofJeEISgom+HvS0HkVH21EkM9OoW7gAkco65NUsgi/Aa8LOyCD6+wcEkFBRMUALuUnLqPA6fQ0szkhR4YErsxkVvF7BoJoXunu6pYQjIcG1UABXBlr/qL4rLIhZl2YqhY72dikqxuJjSGFaFpEEONhcwTqDBADXCGKKgwMjIipysiKIFeeLrOFaQEUCP8O6yjm3sXPWfJW5qZX1gMgJEla8z42oIHEpK5yZGQwO9MpOlNlUmreEqc/NaZwrBLCoRjUQ41hbm7qPcnIjIhRY43KOjCfMBlNAt6xm5vLs2KHL9+K8GslimHvEGqIAdHV2qmZhPoeRFZYXwvPgY26Oj9ZPA7MNDiIqZhUVXnjrrBjEiApnoaNamQrX2bBNCwgVAHviw8VGyL/eCxF3VhZevfXfTtp/9I/qijzBpkd7LfeZHjnhjSuzzrD52HtYF769h5qOWE/KbsSaqgQtyo/fzrWU3eo+NSWF/pttUnOAkqx/TdHNJibPw96zW5LNlrNh5T6F8w33bx7oqfHhOqeNGDGLEIV/OhCSYNXs4wSWwQNsPMBKx+ZIA++82O/m9isCzt3jxB2MNa95hJJZsni5DXau7J40f3EC0XMZFXwdz5/ZY1mHt51b20+KEKUCfiquupqfRQvTktJyTKe4P7ZcIe7PlNHoY6uMqUKoGGZ+luwjOW8JdLJuPY884meq+3eWEDS7UvvqpoyQMkUKBY5bHqvtw9jYw9rAwEnrBvZyGLwsA85ZVEhxD8nXC8BjFowj3wiIct9oRJQB8ARj2RFu84qRVNzXS12hRkOHG7hrYVcI4Bngz55nu7r9OSfJMtgUXiRpBfS6Pb+XQ8l9JIluBdPSGz5jSkNdVwLVzLFw4B1VFVQQ8MOosvLGupQ8DvDlfkbuBWpWMjWUVNAzmA0h5/cSiaBOZvv+Al9nHR486xgDJmWnk0yZxZPUDmYbZYqoOVWGgdvmvqDsG86VbBzynuOu36yCStfY6llrWCB5RJUOO7cNiPdQCtkvexkVTlnCOVigKK+Zc7vQve+AUbMTc8fjCCq9Z4YZHxHLMEwkTN0xzbFic03rsTbU1jZoTUy6wGNya2mRGc5CS5SGYTBqRvVyCVztwt8bEUyiwuy/PTJAxIZTTXjNkapPebzCPagSMqzFWz94rPwd9z3ci3OfzbFqGRTW4T82RmtoO48iO0+4np5tnbdn8EKv9RUI1rMJVgC2EZ06Vt4XzlJN8zDvoySVPAStzX3EO9dz87XLbVCnvud0ZHiUbIZcrqCNHzs/3pzI2sxT2J/YJMB7aI6UM7zJCB2zq/b2hbTVYuYk11DuEfj16ZTCe92b74QvOcs4/k62ee46ydHDva9HIMv2VrZsNtZJJHIWUCPsCQ/eC5Z/YaSb50Ki6+safJUb600aOvE2vF98cC5M+4JrEiKvPODehtictZ+tZdYwYufAxiwfGm8uk0X3nLN2UrOxI/35PDnJxK0+8Ygte1tPLXbCORIBaeNLGa3KmjVlnEhkp/LgPUVShvehl6mhdcUpf2bXTK3TZiWnPbtyam19UjaYq0k8ssj7TjZGbF7SmvG2ouIt4+/tv/wPOANrYpT2m5eoVwyqEHESVI9VtsBty0gwIIebU5v4NJk54MXdY3ajuiAovh8XdAtUUhuR6/CyjbrdgC40iBMMm1Ld3916Z906sssxptTk6x4jqnd4y8ZilkV3RbmYa48IcL6qUoZIVuVe6zGTlJ1K+jhjJIv5H7k2eDu2WSWJs1cR4ODk1DYxUkpr/nVeN4vH/qqIPKEzyGxJzOeODx2TK2iUueEmKBXYrttSnUxuUvSUHB5zbROyyZa9DgF1+cm70ybh2XOujZExynrMNTvZROrC0HkuWCBZZ4PBZCpAWGQ6QoaTMb8HC0wWzFRUkJggwMxCkwUp1RbnO0UFQVraSXFRZ7HH3IPR0WFkM6Q4HHW2BSxSZzA+PoHxyTFZRXAssYAqihVKMTE5TtBxVL6P1dXV+jdtiuNxkRU73ngD8fHROaKCiorMDBYtXSAsjZ343DzTNzY/l13BpSp6CeBOTtHyIGrqAicP9TblXBcIMBDkZ0dsNBoRMMuTGJ+c0OJFMJSdziQjCFpzoWLRa9fGujII8I2NjGDrG2+irLQMZaXlyC+IacOvLpxkQiqFru4utLUekCrgaMthgRCLFy9FTm6eLIkKy8skWyUA7XVCeUQFzz+LQp4PFi/M8OAYonSaQC8XVQKFNoZ8Ot98rgeM0OplpL8H/Z3HMTU2CF86hVNOPRXldY0Y6BvA66++JhuvidFxywEIBpAVCZgElioLBkETxKG/OD1aA34jIuR3n9H5pvUUMyBCAZP7knDJjoZF9NC7tKu7WwocPrJz8+CnT7dyBrJw16/vwfyFi3Dx5VegsLpCiopoIBs5wYgyUiY57gm0OksDHhevqfcY5RgaHcLQUA9ajxzAvMY6DHDs7NiJ3bsOYsXyU3DRpZegvqEe/qwQ+HzeCyR3GSAeK8hT9zMDeA8fbBGplMPgtGQK0wppBNoOHsPmV17Hpz9/CxqXLIaf9lrJBMaHhrF/53a8+MSjGO/vQnpqEpPq/DIiUx0fLk9BQM7gsMB2bdRSJLrsZ7Mqo++vyVb5Gu878v5XoR8w4Ir/znFHVUVvb68saqgMCOdbmOv08ChWL12CJYuakJWfj8Wnr0PfZBLjiRmsWrka0WAI0dxsJP0pHDzUjvFUAm0dHRjo7MZVl27Uxpf5ESSs6MteVl6CXc27UUPrp8qKP0NUZDmighkVQMqfQUvLMZTFiqSqSPumBCKPxqexZ/9RHD60D7++81doPXQYaZITVJPMMBx+GjPqtnPgjDe3u/kqBPqyWm4FNzWe/YC8Z2kHqK5p/ntIWS1UVLCDhyQoNz2cg99//Q145zuv1vyiYl0bWfqmcG1ifk/qLyIqeK3YKf1WooKFOSdhk0b/V48/JirMKiCB3bv3YOuWTYjFApi3sBaTU2kUxRagubkV3/v3f8fEBC2fxjVWPHLdCGnbNPjcRtEjVLyaQFj5dBz1NWVYe/opWL5oPipKClFRXIpwKFv2C9zgBrPonW+B2wrnFNBI1VYK7f3D+NX9D+K+Rx5CJD+Cmz5yI6656hqUFVegtKxStkwc6wxqPHT4KDq7u9DYVCeLu6GBYXXk19VUYyo+hu1vbkZDfQUGRwcQzo0hK1yKPbuPYO/eXSgrK8Apq87E6PgkMj4r9plyOjbcj727mxGfGMXQ4GE01IVxyUXnoTBWjfHJIPYfasWML4XGxiZk0tk41tqDtuPdyA6HkJsXxv/F3nsHSXre54FP59zTk8POzOYckUGBCSREEiRIgkqm5KurunNZdpVKJR9PlqwLf7skH03Ld5YsS1USrQiJMimBFAiKJEgABJF3sQmbd2cn5+mcu6+e5/e+PQNI8p3/NAvDQnHD7HT3973fG564tnQdE6NJPPz+D2MzH0alnkYkkkG9lUcs2sbW8grya2v49je/iReefx5bWxvyu1fqVfSl47j/5GHs6u8DKmVksyn0Dw7o+pRqNc3DVNsTCNo1MoqDe/ZicnQEmWxU4Hg4ZqB4p2sACXUddDbEElTgJ9xaUhVhx7n08rUZfOUb38a1Ozexf880jkxPoVutoNaqotqu4nM/85PYc/JDmMsH0EZUBBBB4KHRMdblIL+5gW6rgpvXLuLWlYsobq0jk4pieCIoIDzJiKLkEOLxIbSadH3GEMmk0KJqrtnC+toG9u07oDHBWLKlpQ2kYkm8+r1ncfPCa5gayaDbLCMSsUgVRjZFYgH1T+Q3qrh59Qb2TI3g1Mn92LdrHCNDY8ikB1Eqs2ejJGHBndkZzMze0TyczaSRzWSQy2aQk7sni2QmhWgyhTCzhRmDEgjLUcGRXik30G00MXftCtbmZzE0kEO+WgQSUQwfOIb4yF6VooeCcQRDUXVUMD6T88BmIS+iwju1tP9ye1ESFd61IGW/i54jOLa2uY75hQUJLdivxP0i1YeKvqCjYnVVexoBkc0mFuZJVOREVDS6psQlSE83AfcTdAwxHqTZ7GBjI4/F+SUkIgl1VEQjHPdN65Vz8TcG7BiRoigH7gnYr6b8eK43LvqJREXXlI8EKNbXluVEyKToqjHwWwpwPzm5rGj9mfKx27g7O6vX8ESFBDfcL9H5UyVQ8neJChbGc76hkyoZi2vtoACE8xJJG09UCHCKhEXU0GXiS2sLNze1R/WOChF6LoqFcxznO9/PZi5Rc0XYvpfK/G2FpVe475yBPaYucsDFgAhoNnluDzh895y9DYq9829MgGSgJr+0Z1ec1HaBswdfTEVrRIW9nqmL1SvhuhX833m3rhzpThyl/kDvlHAgloEv7uTmHBYKTfIEtURe7PhwGez+WjlhF6+XwG9FXhhQ7c8W/vPwM/YIWbee6ZruJCj+DpFvojivl/LRUvqZdhB0l5ukwbucHO4SW4egEUp6OafwlsPGXWc5jah6l1CM5y8D+fgZdFbrOWbsrWxHh3TlnKJriVVHOpUAACAASURBVCIgCrHyWwUMDA6pn6LdZD+BxeFIKB+kEIeSDEbTjouI43vjHkXkiW96d1FgBLF9n4MHCklI8rXsEjogzAnarAPAiQscQC2gzRHYigVyuer2HFrZrp3pTc1vufGuo6D3XBOYJUBs8T1e/ML1x5wI5qLimqP7/m5riy68fRbv5DUlvZEM2nc4lb8/7zIKR70Een9RfQ/nWt8pKTFcvSHSls8yY6pULhyzUuDtyDQDbb2CfOc+msIB7q2ZQuBjp3TOqtUlHOLP5JrEOGICo4lUEsVy0caRsAuqt6NaZ71jlw44zjvqW5ATui13F8kkuVOIa7gzv6nnLR7I1PRtRNjz0TCBDV/bnFHbpcSeXNT+1qvcXUyNB5jtnluqhNT/FC512shksgLqKW7w6QreicNbxvk4nclo3iGJZkQRkwUDKoGv18rqFOX+9+7dOUxMTKLdMRGrKDiCtEE7p/g+GP8ceR6R19mAbPtM+j4SRU0WAVuvgAkmHQnpzjwcOxJDuudY4991yesaiTTznSeQ04T3wAtE+Z4VyeMwJk/cMDKIz5R1aNjA9eNaY7pW0+cjliDlv6KqTXwqR0GbgrB4Lx7cx7VxXy7RpiOFvBrfMDLraRCAzflS3ZMUEfIzmpvCjzE/d8ktxfFCQtSNFX6Px928K5yv4/EmjadIROPQg/r8ewLwPq2EY5M/TwkZTPrQ+cfisnZY43o4mwm6jBgwAspccvzyIgjfcaPOLU+QemeACHXbM/j3rP4Hdz6z6/R3v174Wqr3hx94koIm21/4Ofqdv7ZS7J1kjf5ecUou/knPjwf+jbBSf4cwOFvXORfwunvM0q/P/Lz++vFNKVrOO2dc+beRMK443gm+SGrH4hSG2vnU5iQjgTwpZ3O03QNFUsnFZTFQilT30Ydu36V/6yKvFGXuXEr6nO8RFX/vWHrvD/87vgIkKixLzS2MPsfSManKPXMbTG/dtYmQD5Nlw+nBF3tt+gnbTBq7SCDXb2h8kavU+dGoFga/EfMLiSkKTCnnM9V5KJGy2IF220w1Fzi+EidXKxnr7bHcJOAnEk2ELvdNiw6JANojlRFoiwivg1+sesKdnrzHfrJXs3CT58tuCfJ7x8n2m+DPjkmprBxb934EOrpsWWNdLeNO75MHDlljbdK2xdvui194Za93tli/8SGw6B0fZPo52Vlckx1sFH/FrD1wA205/fqS8spioPzhxzzL23wFVYu+fEh/LrLHO2uMqDDrcdtsx+gq4klZft2OYnq42SVh4YmLDzz5E5qEGYXEyZbXiJs5XsNKpaisZm4+CBAqszOe1KLAfgLGIRBgzG9uSpEy0N8voIbvIZFKYHJyUmOL14v/ccPx8osvIr+xhqnd+zC9Z7+ABwKLh44eUOlebnBId7le5aHfSpRorebPicdTypGU+mOHMlG/h1lBa9Wy7mkyHkOa5Y7KMC1biR07FjbW5czgQWNoaAhJZmM7lUm5UFQXx8L8PNbW1lQaysMOo5+oNFWpb53F4V1cu3ZNmfAcSxdcmfaRo8eQyfZhfGoSwxPjaLq+AsYucBz5jgpeW26E+TU3N4eDBw9q7BGkLhTyGhMkeXRjuiQTKrrOpVIRsWgQYXRUDLu1uoB2tYRooIOTp89g1/6j2ujeuHYdr77yCiqFksYz7fAIWicN7x0tqFZUbrncoQDL0xN2vduWI5vr68fYxASGB4cs6ise07Wn6oNRPQuLi2hU2IkSQqq/HwXGbnG8t7v49rPfxmERFU8gOzqEWDKJeCCKvgQdIUCZCvKOzTv83HzudxIVJKkKJCo2ljBz+zoO7t+DtZVVnDt7TlEuJ0+exsc+8XGMjo9x92BxVJEIctmcFXsx7qxZx+bGKlZWFpBJp3jK07NDzTrJhdXZFbz4/R/gl37lV7D/6BEEfOl1pYKn//wpnHvpBTTz62iz9JZKL/ec+flOh7FmExsbWyIZOPY4l253TfDQaRZYPo+eXOO/F0nkbNR6Npot5SWPjo1ifm4eK0sLQKCNZD9jbuKI1BvYNzyMD37gQcQyaew6fg9q4SQK1Q4euPdhxFmAnImijiauXJtRzBOJitX5BXzuk08glkgocZ5OIBIVo6PDPaJi21ERRB1BXL5xTTn4Byd3IUHlFh0VQeDKlVsYyQ1iZHAA3WATnVAAhUoD3/jm9/GXf/kUrly6hHqphLYKB9uoU53N/zVs7HMONyLCiiV5XeJSCoZs7nFkJqPPeC1JsErlqMOLRbewC4Rjl645gRL1mkDGf/pP/xkefPAh/XweegTuCDRhTCKJihHFXb3bUeHnUJvgu6i3G8hvNcAy7ePHDiDX74kKrhn/8MZiZ0E3VfYEa2/fmcH3n38eoUAV95zZj2x/FrU6VXU5/Nsv/RZee/0F1Bt5tOp0iLV0wPdfcuOpM8fmCP/SWn8I3AS72DeUxoff/wBOHj+MidFB9Gey6M8OIByMokt1Z5hkLsskmVHruhSCbBvg67WxvFnCD89fxL/5f/5v5GsFfPrJJ/AvfukLOLjviHUvCHAJ4PqNW5idm8ehQ5yruxjIDUqaeef2DLkqHNi/F3MzN3Drxls4eGQ/Gh3g7twWXnv9bbmBpndPYGrqGDYLFVOJ8wDQqKlkvV7OY31jBbdvn0UosIZPPf4RTEzsR7OVxM2ZRVy+ch7ve/ghZFJDKBY7KBVrKNfKyBdWMHvnPA7uG8b9D38IG/kw6s0cwtEMynWC+BEEGwHM3rqBP/z938Nb515HqbIl4otr4P7pMbzvzEkkO230xekW60c8mUCXlvtuUP1N8wuzuDtzBzEEcWBqGvun6IjJIpNNIEFiNhhCsVTG0vIqNvJbaHbCchnkclkMEfxO25jm/Hr15iy+9s3v4crNa9i7exIHdu0SUcGopWK9jE985kkcfejjWCoF0WRLfZuRBmEMjo+Au4at9QKS0TShemytL+Hq22dx68YF5NduIJuNYXRiBJm+LFLZPiSTfYgn+hBJjqEFggQsht7Enj37NefnGf20aI6KK2dfwQ++9VeYGkojHuYeyRwR3Es1OzVUag2srxaBZhdHD+/G2FhO0WKjwxMYHBhHo0HXkI3bzfwWrs1cw/LKMqKRMAZyOeQyGYHb7EbK5LKIJhIal22E0GEUE0kLEJCpoVWtY3XmNvKrS5gcH8Pc2iKSAwPYdew0GrEBNDsEaRlVGBGRxP0MlaWFclFroycqdopmFGPlXLy+TFviEhEVG+rOIgFPEKylEl/be3Iftby6gqH+Qd1DXo/FhXntA1imXWvXFRupKMV4VCB+rr9Pax/PtGtrm5idmUMiHEemL6Xi60azJiVzDwSSSs+inxS70mLeMpXd3Kd00Wjx4EygxWYAEhUEDdfXlkRUZNNpE6/Y9r73ZcIdO7Qr2qfTwczdu3ruRCakbK3VHqvJvq6avkfuY+eoMLVhXEDO6sqqIiI5RzOqj6+5k6jQnoJFxn0ZRT/JWktHxQ12VEQEIhqwuU1U8NfqFnDnCn8+oVDGK0R91JHOGXJXBF0siTnMd3xi/Z1U4Z6ocLE2f9+M7QGdd/+dqfotxkWRrW5f7h0IXk1rQBAJkZ1nAgNMvdrSC738nobrkmUFeXDMssgt2nA71kvHAInCDJ+iYp3j3L+2zg5ufHqSx2KB7MtiKLbLsntxTe6sxveus5LLqDduxEgiWwPfcVl7sbf6495Z1IBdc4a6s9FOQZX/EXI72G9E5joyTOcXV6DNz8CxoFhX1/Mh9S2LhTtWhmyCD3utaqWmxAGpZp1aWT+j20WtUkJfrk+fgSCslZTztaUPtgglqtF53FJcUgBjY2NyBVMtr9sj8ZMDQB3/4mN8eDbhOcTHUfq0Ap/3r7OoUwPL7eHOi1YYbUSFB3lFMvh+CCd4c8d0EQ18Tc5tiuN05a66BT6lwF1jXjc7A5sjwsaPEUs7TFbbc4OAWwdSyunvCtt7zhsHdsohYiQv9wpyY5DAcyXGIundnMHxy1gbnu3oeOX3eAW6opBcRC/vo3dNC2D2Smfu75yrxA8/f74m1lCvskjdRJF8Nnn/iUd4ARBfl2p0uVKcc8neW1j7MH++J1Fg542QeiC4FnrC0FyqRizIvapiIOuq4V6I90RYiltPBL46YkKRzyKc7TPt/GyesJKoke/N9e/wHMp4YzmFHODuH0ABpO7PPOgsEJYF80HqKkqKeeXrzs0vYHJyCs0WO12iqrakAI59hCqP5muIDDQynGPVg6/e5aO5xYlGOR7k+ODaUK+bG9yRAhxQwogoBlL5teEg/jrw59vPMZep37Ta+LU+ED7jPI/afNMVucDPaM+4bXR5/fyZSe4N9gE4pb7vrdHa5hTrPlKcf+ZFCj231Q4Bqif2PG7Fe8bPKHxMxLiJpvzc759VXjuSZv5z8DnwnQmeVPEPmEB4ET6MEtqZxGHg9bbrxrtpLGbdOnsMW+KYoJhv53nDHDcBIyidANf3y4rw5vPEz+rGlAfKjQhyeJhcSVZkbXMJ44sMn/IOFU/I/X0cJ//ND/4605tL3vfpQq+71ZxoNu/4lBJbjzhP23zK8ePnbEuGMYJje7kgWmXnA+FlPgJepIqLSBbJaH2wvt9K484lHYhAc/O4YYAW4+S/tP45B6jcjrSvug/rCXw7N26T/PrXevv2HvR6WsPsa/vZ2S5/tzQcJ7R4j6joXf/3fvEjcgXuyxGEdQ+EJwLcok4QWROZU+7zOeD3EixjT4EUEc4e5i+HcjGdukOldO7h9YSEsh8dg6mHzqmJ/IPvH0yzAroH3zOPjs3ugeXeyaHFzjJY/b+xn7Ntefa/94eQUMQmdb9h1gTGycApRbwivXebXWO3n8AUKeIYbjkifLRUyJQBRoJYHh0ne76OirSdWkG/7k3k3JBwgbTFwTa4PoPWVNVepScnhT8IMzKmVrW+ClniLIO4FwHlOzw8E8+FJ0JSwWVhsuyQbDqzid19kArW29I4cWtoGCHEQx2BFx2kqARkHqbiq5hJaBMqJ3NuWHjwpntCeaH6Mzoq7NdHf+wRjR12PegA5myOXAjpNiiXK4qC4iRPJwH/4zXh9abFmp8/v7WlPgZmUnLjyIghbqb27t0r5wIXBapIWGx88/p1AdxTe9hRsU/gEMfovgP7tUgPjY7qelcY86T33pJleXh4RAVkIpMcgWEbdJcvyc2ViIqKwBECCJlsWvea5aK+H4WdG3xOSqWKniWCDH39WW1c61X2G9QUtUR7JsF6btQ9+Gy9FCWByfx5o+PDWF9ew/k33pRC9dixYyrTnt69G9nREeW10tVh97OrDHQrZ2MESU2gKg9KfL8sAyc5wnvK98yODh1UW+zkYOFfGY1aCdXiqsDzrfU1NCtloNVQNMnY+CSO3vcwylQut1t4681zeOvcOdliqcjsNisaBxqPVKgzl5tgEQ8KXapOWtrwC7hotdGX7cOuiV0YHB7C8PCQNpV0o1Cdxvu8vLwsAivbP4Ts0DA6sRg2yyVsbGzi6f/yNRw+eBAfe+KT6BtkMXoCzVpTQIflbzLahxErLEuPOOLEykH56JfKRayvr2BjYxVzM7dx6OABdaWcfeNNnHv9HO659z51VAwNDwsgY7Ywu0A4n3FTSUJna3Md6WQcm5vraNQriCraKcYgV1SqDdy5fhdff/oZfOFf/iompqfRiXDOAqr5DXz9qT/FrYsX0aiWBCBVq3Xrx3GHQM5r7Eygimu9UEQmkzLnSojK0nSvy8THuimyTf0MBvTwHjN+gyWlfH75HI2MDOPY0aNy1BBYWtlYR7Ivo7iWeCCMgVgMT3z8Q+jLJTG4/xA6qX4UWxE8cN8jiAUY6xRDO9TG5Wt3UGu01I2wOD+PJz/9GZGMfP7Z2bK+sYHx8RG8de68VOIs02b0E8dnKxDBxeu3NVcf3TuFVIRAWBCtYBCX376GoVw/RocHddAnwHhnfgm/8cXfVPxPtVzWuKSDgcScSs0YL+hIOsYwSBWprN0gsmkCeEk5kgayOfT3pTXWS6W8YubyxRK2SkXUCOLLvUeyNC1VM7Pmg5EIMumkDqijIyP4Zz//8zhy6JBOc1LRaB6zDfHY2AjGxoYt2vAfYBw8cLdVLOP6tZs4ceQgBvpsY85DwH+VqdAMxW+hEieA1bU1PPvsMygUN3HixEGcOnkUiXQf5haLOH/+Fr74xX+LtY151KsFNOvMd7WoPgGV3Cjr8xJoMYJM1cR87x0eFBsYH8ziI/cexcP334O9uyekXGcRPEFqBAkEd7UGMPeZ8VEdgrxSl3M94XzQxVapitsLS/iNf/+buHDjKh57/GP4lX/1azh25JjA7VA4iuXlNbzyymt44MH7kckkUS4XMTY8KgCKirDbt2e0RrCc/aUXv4vJiRz2TI/hwvm3sZFnjFIOzU4EBw4dwcbmlhMhdEUktpoVtBldGA1hZZXl0d/ET3/2ozi8/xBayGJmpYaXXn4Re3aP4vjREygX6CwLIpKIoxMs48LZb2E0F8K9D7CjIoROoB+BUBLl6hbSqQSC7TCun38Lf/B7v4WrNy6quFqZys0GHjlzCGeOH0WC+bwqIe1iq1jCRr6oaCwqGgnO1islRLsdJKMhjA7lMDzch4mJEQwPjaDd6mLm7jyu3rwtZX4nEEA/ycaRUQwNsFODMW5FHX7L9Ta+/q3v4cr1a5iensDuXROo5QvqCarUy/jgxz6KUx98HCvVCOr1CLrNFpLRCIbGBxGMRbC2vI5kLKN7ydrVSjWP1eV5LN25hSuX38JmfgmpDKMWSXYOGGicYJF6P9rdCNbzNeyaPiDn2+ZWEcvLq8gk41ifv4nv/PVTSHbrSNKloxiZJhrtughKnrdIRqRTWUQidKqlcfzQAYEjyURGBFaxVBHRQ0fB3NIsFpeXsLbMqK4gxkZG0J/NKDaLRB3FCwR7lD4djCIUS6EbCCO/WUKtUEZxbQXl/Kb6pJrBACYPHERibArlACMDCe4x0iiEra2C9ggkKwsVIyo86W3ADEEjU8MZIRwWSaD4Of0Zo5825Iokgcli6gZLUJnX3jYAhhGWdFtwLiSgsaSOiqwEGiRhs32MfmLvkMXT9ff3qbAe6tBYx+1btxCLxOS2SKdT6nQydW1vlyuAgWsS5yn+Pfcl3POxG4TX3QSTFLYQADIAcG11UUQFY6gUS8qDM593B9x4sEdOAOUxd3B3ZkaCI15/65Fgsw1B3LaLNLSYVHMZG4hKooJgwdrKmimaGX1GlWkwILcmnbYRxXdYLjr3Wol0Sn/G79m6vqHrztg+f80NEDHRlJWBmirfx1NIJe/ALgF7AskMTPDiLQ/iCwZwOIeEKi4GV+phnnl6dnIvet+hfHfRFwYgO5e0j4Bx5xiJvlyEgxUnm7pYZLiAOgciE+JygL1I+LDt3wgiq8/GvTfr6LB+QV5jvrYX8Rg4YsCGV3ZKLx6yIlvtt92HFWjsVLp2ZutoPhbA45TS/jOZIMyU+B5ANXDIFbVSRes6LnYeoTVOebZkDrvOSxazwvvG79/5ZWcBO7N4t4rOLA50tDOpsWYSublznj+jWf+hkVgcBxTVcH/kgUVTPRvIprOXK1/V9VJ3SEAu2nKpiOHREWW/5/NFA0E7PINa3JbEeLSnaeQbCD04NKR9Jc8sfA8EYHmeNpLMIoEEegtMZ2pBuTfP6B66pAEvvLNx55T+0uI54Np9nz6TG298xqRmduXBik1SPr05JryAxYQxJuyja5//b8kHFhNFhb7iWJ2oznoHtAPQ2YikjURBbgyZk8ecRwSIGeuqManzuZGm9pktQtMnFnjxmsWV0h3QMRW767H0Cm/u83q8l+sOoHhP0ZokrDSOLKWAX3xvPhJUc1cgqDMWI4N8h4kvbBYQ2m3r3MovxkrxLGLktBFingDpRbK4a+4jxnQWEzlnz6bWEYpbGtsgqGKcw0GJR3xpMp9dYRiuG8EEnuYW8POm78gwwaPFVKnLwj1DHsjntdC19xFfrqCewKnibliu3esTtXWMzxTfD9fn/j7e8xruzs6p67FMN0I05p4bqsSN4DOXkHN89XpJDOeRM4f4gYhC6/ngnp2dI9ynC9tw/RS8oeaY4J7S1lQTEboIIte5wzHgRUI+dsg/AyJJXCyWsAWHg+xMRvB4Cu8lPzPxmjY9ps5tLwU/STTXQ6Hx42IU/TwpB4Xr4PHzKYWh/vmwz7kdI0fsTF16bm7xAjpiJYoh45y6o1xcOJs7L3E86sypcnQ/Vxg433uW3VgQ5uRcEiJjNQ+Y8Nh/Bv/eJPh1cYienPRkp6n/vfPQuA85AHh+czFLvH/C9ojFBTkWLPrKrwHCs9R36UhFAe7WX2IOK/s1x5yIWhfd/so3sr2p/32fLrr5zZQS3uGiOVHCCj7jftm0uFrFILp5XLFdIgK3SQtzwtjP4hpgjiD7+VrXXeS93XcjWShA8Wu+3LAivdiDY2ICCRgcWcd5juPAE/YiM52Tz3pNjIzVPN0Te5CdtevgCSO/ntncZVHsFjfshHUwx4hw1veIih8RdP69j9G7AqcyVnwkpQpjWFw+oGxFrmBak43baDo8Xw8iJxofw2TAqOW89hT6TtEjBwMfMMauuIdS7gEuak7VQvTcs6BizdmnUOOG2Suj3KZRFmhfCuWthjyM2GQgFtjlsXJxoHKai4I/TDp0B+2ALRxeZWXv0VQRfgLxuYm8NuGIWcL45ZUT3j0iYqFp5T7cgPQWK6fa8CovLZrMHyaz6yY8qQe4cdZCaJmVxgRbubbPqvPKAyrsee0U4+IAdG0IXZarV+P4CVATsTtcyQS3o6TOu3WNBfY2U6dkcQcS+9lm3bVDrS0EUkfwgMTDRcuuC1+T/5kioW0HYSr5Gf9Eu23HskaPvf/9iksSWOY2sVReM8KGYBXfMzcBlWJJmy4e1rPpjBZxAqy2SbMDLxf19fV1bG2uoVzasgN8LqdNlzJLASwvLqJWJlGxG9N7rQiM42tweERuBoJEJDUYUTQ0OIhQLIqtQh6haAS5vgEtylJMtb09mjmUNv45JkSUSOloIAEvED+vPQgshV0RQErAnRt9OksY30ACgUSCFph2R6RTrVKX1ZhKSqlMpZS+rbG5a9eElA8rC0s4/+ZZZOJGVKTSaezeuxeZ8TG9BokQoh8cY3QtkAwgUM+DLC28HD03rl8VmOEVlhyH/f39ys5UyW61go3NdVQL6yjnF9Gs1dDk4YR9NK0W0okkwtEE7nv/o70osGatjh/+8CVcvnhJPzfarhmgwdHKaDFuYBxZx8MeB626bGhljUQFpI8MD0spOrmLXSMRzM7PI5PK6CDI9z84OIJ9h48hlE5js1pHvdPBytIifv/3fg/79+7FRx//hMgI3lfauDmu+Bp0ZdSdRZx/5t0G/kBK9alcGwuz+nm8riTD3njtNbz56us4ffoMPvLYR+VCiNLl0agrNomExfLykj4vs7hJTtChwgio1eVF7J7epR4OFs6eP3cJX//6N/GFL/wKRsbGEEjGEI0FsXT3Jp556k+xdOu2DgOVTpMnIM1DUiIqN7wr9dhmPo/NUlGb+1qlqpgms6ia8j3qNv3MaafDh5+PHQpkRKhQZcE4YwvYvzEyNowH7n9Axa23Z2Zx7tJlRJMsr88gGogiEwrjk489jF3jfchN7kE7PYhGNIt77yFREVGcTTfUwaUbd1GrN9QHQ2fQZz/7WXWbcK6KJeJySBFsPUeiYmQEeyYnEGaZNo8EwTguXp/RfHJi/xQSxN1o5Q6EcP7SZQHikxPjyiRmP8aX//gv8Lu/+7tYX11U5BNdLHQw2EaO14obdkaqMKYQSEQiyKYSyKXjGB7sV7dJNpHGULYPg/1ZpBJU8bawvr6KlbVN3F1Ywt2VFazk82i0yUFEkMsN6t91SXTF4/o3zUYNJ48fwy/+wi8oksXi3KjkssMDVdMkZ3QQfhfQsr39YNdJB1vlPK5du46Th49gKNMnwL/jnYJ/716F87iVkaPLAtourl67hqef/hoOHt6NBx+8D8MjY0AwgUKphn/7m7+Drz/9V6iUC4pN4ryiDTTjXryqWyoErqFUWHNPEBbhGO7WMZSL4+F7T+CBw3tw9MA+TAwPIZ1MIRSJIZLIoBuKimSX8isck3uv3eaBiiCEkdxcXxmjt7i+jt/5gz/As89/Hw994P345V/9l3jwoYfQ6QRRLtfx3Hefx5Ejh3HgwD6VsNMtOdCX09zMeaRWb+HW3XnMzi9g9+QoVuavYXQgonuyttnC7fkGSo04Dh7Zp3tK5Sv3/9zeNJs1A4d5mK8X8K1n/gRPfvxBnDl2GJ3wIG4ud3D7Lp//G3jkkfsRCqRRLEQRDKeASB0Xzz2DsVwX9z3wKNY2g2gHGDsTU+wgwZtOA3j1e8/hz//493Fn/iZqrYq6E0KNJh5//0kc2LdbcxwdAfwM127NosES4HJFZOPE8DD6Ugn0p2JIxzmfhDG5axSHDu7H1K7dcgHcun0XN+7OYXltjfg0JqensHt6GqPDo0jFU3LIXb1yHYVyDW+ev4S3r13B+MQo9u3Zg7XlZSQjzPnv4v4P3I8TH3gMG600GvUkunUgGYtgaCSHSDShGCKuG+bgZM8SY87a6NY72Fxfx52Zy7j69hso5BcwNtaHifEhjA0Pyt0XiqTRaMcxMLYf8cwQtgo1LC+uI51IIdSu4Jtf/RM0N5eQ6jaRDAWQTMYQjNkcVanWsLqxqciuxaUVracP3nMKe/fs0bNF14FUe+GIytsj0YCu39zCAhYXFpGIRTG1axRjQ4PI9GdF6JoanTvECKKJLLqhONbX8thaXcfcnTtIxqKIp9KIZfswPL0Xof5hNMMJqf8JrnDTVCyUtdZzP1kkUcG4x2i0dxjvgZoC0sM6zDIGSk6BYFjA0eLKFpZWFjEyOoBkIipHhUi9Fvd7TaysLCkOkV/lSlmCAu6JKrWSxB8kKrjHYPwUX4OfS+LYjwAAIABJREFUjY5POpgYJ3Prxg3te7gfYDRKpVpxyjw6KeSN1v/zWeGzVK1b9xevTbPB/QGzvx0Y64Hybhcrjqhgt4ZcFgJMTSnrwW4pSzlWuG9stXF35i4CLDlPxRTBFXZEBfe1vnsp4t0dAhoYwWPRT+wD4efj/sRf47m5u3p2IiFzJJOoSGfTSKZ5f+0+bF5ftQJuOrskMAlZfJWLa/HOYMXaepDAual9JI13XffUibwZTsqoiBLnpJDvuweaWaQFAWdFtOjauZgip7D04FmvMNaRCXJa+5fwNm53hhHwqBJgy/XnftNn0wsU9RGiTv0tIkbv1/cdcCHxJx5THqv8VIpTB1y5n2GKWDsDcK9EksiAcR+fZACkAY5GzHiHxk4CR4Zcgc1WEOu7HkSWEbhyAJdXM3t9q1ei6gym/gMCcSS7qbA3gRffmwe4vZLZAHS71rz26pJwzn6LfzThloHhFgPC9cmD43a5LMbG4oZ55jLSxEYl3RI1kcgcz4qqCQZQLhZ0NuGYJTmRL5QxOjqhNS6RMuEIHQp8v3yW+cWzBR0Y7Ozx5xNGgug6u3QCjQUP5lGc4f7cyB8HsLvYHNvz2VnMx8ZYprn1SkgU59zy6pX0HQKaC8yN0RK5al0kFkflejgU7+uILLupLtKE79WdV103it+iWJyPXUdeQ4tI41s0EJrPr+YMR76J0KXDWkXTvK5UtjPeysaOroMbS3wI6WiwOCObd7S3ZXyqA7C9yE9dFI6Y6I0Tuogd2UJRmxXX8j2aeInRfuocUtG3YQk+woWfLxK3iGs6zY3I8YJCjzk4XELPnoGaPNMogsyVZetZdsSGf18883GNYNypdVOaSppffA75jHlXhn1mc0Ro3FJwJ+LJnjd+JooVSM4x9odudF4rXg/OmSQ7ef189I7AeJeq4AFRi5VyRfIkd3k+77YRi5gwc219ExOT01jbKiAS4zoiWaqwC3PommPP5ibbD/PLx3/7z+2vgyexhOmQuA6Fe/1PRkTZvCVRk55rK5MnMWDYkXPyeeeISz3gPOfjwnoioiCTDio6B/WEpY6Q5DXi9eJ5m5GJdHb4ecz6IygGrWv95TlUynhXHs35WW4mJ4z1a4s+K58dHzPokjBEnDuMh8SwEf3EE7j+2lzF+Y/nVBHpvB9Bw6dsXrQuWP6az4kckg7c316PQ45gtffpSQ2bT6yTyu6FWx/cM2dEhhHQum90S7IXxAln+V74vPFjtfQsG7xk5L+LV/J4m0soUcRci11oHeEufp3ivbO4L/8e7DN6EoB/98o3th0VD30qr3XdnO2uW8MJc60PiO/d3DqaG51bhGOfr6nP4OYnv9T24pwcKe7dLfz3Hk/0z/vO9ce/ZxHp7t/6924EpRFyO50u9vz6iDM/tm0e8VFfdOwT85QUxEdHeTGv1m6b63nv7XxlcxHdUr118D2iojem3vvFj8gVOJWxCWl740e1jG2eZclzmyKvYGHOoQHzFq3jFzX/73sbULfxNQbVFAUiN9ymzCssODF4C5RFRtnER2WAKYRsgyq2nkpDKqW1MTGrqBZWv2HnazhVgI6XTjkllY77OZpsyIxycXVZrQLznQLFvxcBuHRKiE0PKoeUawE/u0VEma3UlEzmZuACygXPv65Nim4hccxrT8njFkgP7usQ6fISCQpQbS8VEydZZ1XkRspPoFwCTShjkVVaTFRw7VXYps7ym3VTzYR0eI3KYm/2PSrcuCh5O6nfVOzsLeFk21MYuIOdJkdmU7rNBLcrPsOdWe/8Oyr4+WsSFVSkkNAgUfGhz31Oh1WOn62tTRQKplbkGLGoIh42wwLDuMljWTE3F3RgkDDwzAv/jfodikUUC1uK3eGvbQG3ci1arefu3kUpX3RExR4VknJhHxwZsc2oG/9jw8MYGhkRkMUujHypiEwqizgz+9kX0DILutQmyiK0wnNeO+43uIBa/AZtrBUt5pVSVXEx8Rhtv+xTCCFf3BKRwc1Ng7FXVCtmsnITlApF5EsluSs41qiUptJy/759eq+Mb1omUfHGWZEFx+moyGREVKTHxlFvtXWtTBrJ5yUupwcLEnWwjIZVbH317csolQoYGx1Dh/FdCCCX60Or2VAp6/raKgr5AtqNMjqtslTqJFMIjpPQJAjT6gZw4NR92L1nrxV3xQieV/Dd73wX165cQSZsG34eTmO0PSsH0srfC6VNjWWRBiz5DFMtGcbQ4BBy/VQSD4tYoMWzWm6omHxocFhqnqHxKcT7cphb28Dq1qbA8T/68u9j3969+NgTn9KY4BfvCwFAEgoCUMT7cZNnSldPRHJ8t9oNLC4uYub2LdTrVRw+fEjj7vxb53D21ddx6tRpfPKJT8lFQTJyq1AQQVWpVfUZBgcH7OAapAq7qOs3O3sHo8NDskgvzC/j5o07OPvmBfzar/3vmJicQpcRFpEOzr7yIp77679CdXVV80yFBXOuMNB6BHjQayOdzqLAzpNyyaLxmHMbT9gcw5gLOigIorMgudWWQpqHQ26GQ9Gwxpg/uAoEy2bkQCIBEo0l8L0XX8R6fk2dJ4FmEAOpFD700FEcOjCJ/pFdaKYHEB2YxLHj9yMWjCGbIVHRxdu3ZlGt1THDkveFBXz2s58R6UVnFNVaa/9VoiKGC9fv6Bk4vm8SyRhVNxG0AkGcPX8emXQG+/fuVo7z9Zu38au/9n/iwoXzcvowI7otgpgHItuYdrstjecwQsgmUyJGJkeGMdhHF1MGERa2ZzIYyGaRS6flsuBzXCgWsLpRxNzyKi7duIUL165haXML9UZH/QC5wRGbBxp1HWzpnCFR+5knPo0nn3zSyGVF7Zn1951EhZf5vHvTEECl3ka+UsCVq1dx+shRDGVy/81EBdfJl156WeTF4SP7MDQ0oEJrKtsXVzbxhf/1X+HK25dUFl+rlgSK6rl0IIechJ6o0JrOAwfHVwN9qSgeuvcY7jt1DPuHc5gaY3k2CZ6kxnU0kUQgEgd1aCryDFKJR0WUKUJNRWhZrCSzVrby+MrTT+OPv/IXOHTiOH7xf/kX+MQnPyEQ/tlnv4NIOI6PfOQjiMVCWF5ZwcT4qLopTMHLE10YzW4Xf/4Xf42hwTSW566iXV3HY49+SKXQZy/No1gL49DRo1hfW9MayYNSLMxDQ0MupIDm76aIih+7Zxrvu/c0wskxXFtqI19q48rl17BrIo17770XC/MlhML9RBHw9oW/xcRgB6fv/SCW19roBDJod8IoVUsqSC5tlfGtr/4XPPP0X2J5Yx5NNFWYHG938JOP3Y8xRoF1OnKJ3bgzh5WNPPqHRnDr7qz2GI996MPo0Lm2soCBvoQKvI8fPYLTJ09hbHQCS6vruHbzDi5ev4Xbs7Mo1Kpynx3afxBnTp3C5Pg44uEIbl6/gZdfewNnz1/ElWvXMDk9oag/zm3RQBATYwM4ce9RHHr4QygFB9FokqgIIhGNYGA4g3gshZXVFQE3fp/GuU7KtTbQlDMviI21ebx9+RwuXXgDlUoeE2Ncb7PKsM72k9AdQDo1jk4nhcVllk/3YyCZwrd5fWYuI44CMnFG/nGtS4uIXNvYxNLauojKO7Nz2lMdPbBbjgqud3SjSNHGGm/GYUWtGLtUr2F+YRGLi/MiAY4eOYCJ0WHksowcZLwnx48VkCOSwNpGCRtrW1iYncXW5ibGJqcwMjmNvtEJBNNZIlNyNvKAzWFXrdSlpCVBzM4IiiB89FNPHKPTv60vFHhwTeN/BMa5Z1hY2cLyyiLGxofkbOFzqKiCJkEXc1SQqOCzQscGBQ6cm8vVElody2WnCIH7UHNWkFTOKjaPQNutmzf12nQTkuDgOtti7r5cwkHtUfiYk5jhfq3ZspJHupm4vnD6MiMmo94cBNHt6j1zHzbQn3MgkQGa/mDeOz/0iIoWZmbuasGNJaOKuozGI3IA/X1Ehckg30lUcNxls5nevnN27i7i7yIq6KhIZjMOeA5g4/qKHCW81lR1ct/BdZHAka+Y6zkRuI+T28TABAMoKBbabv+h4MaDrwJ4HDjJ/aX/XsGwXnVLgMHQNY03DywqJ53AlwMTPVCo2AjnaBDg4Ha2AswdwKnzjHNVemGYVJMeYXIRRSordY4OkQ4+R7y3X90upvZKb0+oeEeFV2RyTBC0M2GW3RuOKznW5UqxgSRlN+85xUk6qxiZ0ovecHG2UkdL2GQgMH++xcVug2hGQFgEBz8HX5tiE4lZHNDrI7F80bgHfXwUhpEw5kQ34sHF5rooGF5rnittb9iQ6MCXnJJk0jXTjTNysufIUJxJUMQi3ZtcT65dvaLr0Kg3kc0N4Oy5C3IMx+JJ5AYGdHbkPpFnAooBBBR2u9pj0/nE57y/P6f9Ec9CBEBJvhlQbCOBZycDPy1iSZ/NZa0LYNN52kA5U4mbQ8LAXeve4J7dXJNuTLqyWRES7kzIe9kjoQIWR8PxJEDSjWM/5kh0Klo4GtNZyzthDCx1Bduc/6JR7anYX0DC0TtILMbE9kG+CJzncwmHGEFDtbED+40sMmKDoJ93Ckip7tTi9RoBZit/5vtSP4HiPrcL23tRQe4a8pzBaGKeVziPq1ScUTLu+SQYarfAnjMjIYk/2D6GXUg8P2tfrg4EIzE0D7geGP7eEyu+P0MxbRxHznHhUyTseeLWxkBcAv6cp4gB8EvXREXUVIJ3HNjqkRIKMKxonffbn48FZLozjicc+XvDbGyMbEfPWJGzjwIVEeBicgiaRkkghTjW65idncfoxCSrsyUsUJQ0neEuT5+RZh5INRCdpAJdPYZL8Brz33BNTiRiijbzcyZJBJ7xSUIYHmGuXO8CkDu1be/bn7s5r+rZcu/XXFi23sot4O4T8RGei9mryrnVuyE8LsT4Yo17PnNsp+K1JGnBrhkXj63Ir4TFUPveUcOlTIRrc66RgBbF4+Ki3PjlZ9ea6dT6fm61GPXt9dQLcSXI1Lhuq+OAqRRcyzifkEgmcaK53CV29J5VSsCcU1qOAP/6vqvKO/rYuUUBYQD6WRxfvHe8Rga023iz62g4ER8LjxUptk6Avs25mgNIsFGgxnJ59WI4p47cV/Yca2w5QlaCXNdbI2yut+baNX7pr7fLtB/4xGbvALUdVWhkh2KVKEWJGMFk0X32d1zffUqJ7QOti8LSFLY7ifyz4edTOQk94eHm753RhtsdRjYXeyeenyv5vXSXGllu19F/eexB48FhaMLYnLOEDhrfF6LrJiKeghITQ/D+ekzOi030XPMs9x5R8e6D9nu//+/9CpxMW2m0qY+sa8CUJbR3eSuUqSM4u8ja5YrZlMGrzYXFEe2cRbj4iLU0KqOnePFOAZ/Pyo2UkQem2ufkwYWMk4wtIk6hQKWIUxf0Nl29zfp2WY4sZG7z5kFJHSxc4aHy/xq0F/vFzF7fLF+2ubWiMU60ZqeWpTBsilNtHNX34FQwXUg5o/fkGHUpN1yebG+ScSonfwjhZsgUHQ4o3yFLsg2ps986dYNtLOzQZWyxu6bafFl5ktmtQ1rIWKpMFbJy97joOAOyWfi2Ld9ExXpZo77DwxX6eEWRWc8ZEUUV3bYNktdRG2iXZ6hFhgeLDuOTGtrEWQwUiQr/XxMf+emf1mfgZoWLPzdXBPN5OOdmhQpvXgOpQ5wqgRMzI6B4uLB8TjtgEtCmon15eVFl3IyEYNcCCaPr16+LBKEboNvq9IgKAnFURw+Pjml8cqFnhijBBSr5B0dHRawQFGap9ED/oEA3qihsE2FMNtVI3CBpI0n1YMyyo3kNqNDnokOlY5TKY21mA1IAMtOzUilJacV7RUfIYP+AQGO6ElQ4Wa+iUChieWkFA4OD2DW+S5uoaqOKpbkFnH3tdaRjSZw4cVzA/J59+5AamVBsTTqZFNlIxTqvFwvR2i0WyNUVnzDYn1Pm8+rqMjLJJGrFIpq1imUhMgqnkJeynxtt/oxOl5+vq2JoEhVU5PMeNFpt9I/vxfFTJ7XwG3gSQ6PWwF889RS2lmYtAsNlz9IhQUKP961O+bHrt0nwPhNkj8bUOUJCg/eaxxHZdVsd5PpymJrarbLeaLoP6f4hxDJ9uHz1Km7dvoU//M9/gD379uJjjz+OoeEhXRPeF44pjqXBQcZaWTQanxUSGMoHdZsHjhOCc3OzMyqSZWk2jyjlYglfeerPMT01hSd/4nPYw3vUamFpZVk/O9ffr8eJtvFkPK4or3x+Uy6emZnbUnLzkEGV58rKJn7w4g9FVOzZux/tYAeNVhXPP/t1vPadb6NTKsmpUaWjwllWGSPQbFiu98DAkIr+Nop5OWRI8HAu5rWjO0cdDMmoIpH6WQLtVDEkPjN9GZF2BN+Yt87omGQijb0H9uPgoUM4cvgIXnrpJTz34nPaXLXrXUwOD+O+E9M4eWQ3BgfH0e4bRmbiAPYfOI1omH0sCREVV27Pq3Twzp07Ins+85nPYHh4QL0s3MD/Q0QF+xs6wagjKtpGVEQpf4+AVM1rZ9+SUp1KdCpDv/il38Qf/ec/Rr1WQa1WFrjHUy8BPxKjQUVxANEAMJjN4ejePTi6bzd2DQ2pQ4AZ/NFUXHFg6XhKRAXHXLNNl1MTjU5YDoQrd2bw6vkLePncW5hfXUObnSaJDPoHhu25b9Y17/CAMTw0jF/4hV/Anj27e4fA/xaiolxr9YiKM0ePvYOo4LPXy/J+x0aDiwvXGC6wVOO0sbzMeaIPPNfpQAcWfAfx7N++iC/+X1/C1uYqNjeWRaB6R5/Af65VjqhQ9BMPaqp86ug6Hty7Cx/+wMM4enAP9gz1oy+VFvgqZbf+P6kiyBaz1uls8RRbiCpnAnE8XJpln8TjRrGE5154Ef/uP/5HjE9P4n/8J/8T/tHnP49r125hdXUT9937AHK5fhFOa+trmJ7apfdixXHM0gXqrRau3ZrByy8/h1Skg+EcHQhRHDh4FFdvzmFxtYD9h08rt5+RBIyLkJqx0dR6QAV6IhnA3z7zpzi0O4VHH3kQ0fQEri22sVUMoFkv4K1z38Xnf/bTyG9V0W5n0OokcPXi85ga7eDkmfdjaZVERRqNJsuyywKe1hZW8JU//DJ+8L1voVDdRCvQQqfZRC4SwecevR8T48PIpJLCZUvlqlwPDcaESFkeQTIaQ6WQx/rSPNLJMHK5NM6cvgf3nrkH0VgKM/NzuHrrLl4+ew7XSQqu0UEYx57JSRzavxdnThzHmWPHVUx94dLb+OrT38DZC+cxMTkul8rN61dFTh3ZP42Dx/aKqKhGhlGpJ4BmCIlIGLlBlsdneo4KD2aaktXAbe5zUoxAq5WlLF5dXcS5s6/j6sWXEApVsHvvMKYnx5FJZ5FM9COXnZDDIhzrRzaew/ee+TZuXz6PcHcTfekG+nMZhINp1JttzC8toVCtiqhc38qjXK1iOJdQnGM2lUZ/KqM1YmRgWOMqGk+q66dcb2JuZRG3b9/A6soCjh87jNOHD2F4MCMiWaBwMIZovA8IJ7BZbqBSa2lNe/GlV/DRTzxu5ESIhdsJRKMJE4jUDdgpl6qmxkynUSgXFMmys0zbOypIAHiighEP/I9EBQ/oC8tb2qeMT44gTJeR4vkYD2pOsJ3RT5yj19ZW5ayko6LeqmkuJOne6TblNOFzzjk8FCZRsSWigmAV3xeJCjkjWxY9KvDG7cZJSBGE53pYYzdPk2WeFGLwWbWJhqSGcvU7wPLKgg7GgwP9/99EhQPtSVpzbo4mokgxTjBOQMTU/AQvFP/KtVgRqg4M10GdfRvrmmf5GbgH4bw0Nz/3d4mKvgzS2Yz2Vfz+TRIV2jMSVDdntC/TNpBckJc+H9dVRjX47Gntr0UcuF44B1D6vbic5D5b29mKuU5KUOBimLiz3ll028s0V2SYuUW8Q8m7KHy8iQlvt/sAvQtaYicXhyPga8f78+4JE2qReCHJv91rZ2cyU56bQMwij+TIdkSDzjM+EsSREtyze1W/Bx1NuWkKW4uX8tG5HCYWmSunxY44D+7/dQ8cAG1gESM4mZFu4JxEaYxc8QDqDiDPq/v5mXleM3dpRySKAE+ecwjyuVgVr2D1im5zFVjPiidXPKjmEwJ4TXndfDGvlRZvn7FMDMI9bVX7aD6nHDezszNYXVmTo4JRcpcuXUVQBctVESzqgGJRbSyi8U5Cgu+fwpFytY7x0WE88v5HNL65J+NZ0KtpfUQZlf8kG3ld+X2KFXGdKr58VwQVRYXq1iDgz8gu68zw8UWeuPLgtCdwFMFDUYtLQtC52YHzHC/2ftnRY0JBA99JYph4xvomKEgwlbCBjybi49mN14D3kO5xnqMNSLVnUi4Zd+7nv+VZkK/DboadP9eAUktu8FGoithzY13F2x0D7QQ0EqNw4kCSKpzDhS1YlIA5TYImlhJI61Tj/Lw8o5lwcDtqzDt1eIblF88NXAdETDjSQGdgAod0h7g+BOIkvSglR2IIH+Bnd8CuB5n5PgnYc74lAbQ9DxiAYmkVVpAtctA5FrxTyD/nfD2ee/mPFCmm8l6+j21CS6kW7N6obfdw8Bry7CpigffE9zM44LhdryPLLqBuR/1YA0MjikalaMR8WG0J1Oje57zK8cSxyNdiggRdI4b3hHX+ZKxtr39TCRJcbxgrZoSaUjCc+8Vixwys9+4MOYW8a8zti32fiQSzro9Uf+aihCjQ5PWRY8vHDfJ6uhQOrXnEFIhlafHbjlHjr3lmZfQux6fdaxLihk1RfOk/j+KT3Dzp3+9OvEWiBke0yJXnEkw8ucvPL5ElS+V5PYT/cN9FjM33D3oBoBGqSgARPsb5nZ+D5LZ9dg+N95T8zomkfb9zXfnOBU/E87P6z28kpu+3cK4sh3MpTtm5nkTvK43BngNzfgQ1nhhjS/JQOJSu+XbHkYSfzoXIp9N3g/j7+PLT22Xaj3zGSuo1BzoSxa9LWiMFOPLs4zpnXZTitmuH50NzAxrBytezVBViP5yT1FHENAP3Xj3pIFKaOGIv5tOef+/o4c8SAe8i7myu88Jru4fe8Wf4nfWFibzi3/XwQruGnijl+qZ4Mudi5LMgZ5pz1/F7bU0mueoirN4jKt5xWn7vNz8CV+BEyjIffZ6pNjEOvNMGl5s8Z2W2SdaYTv/QeqbSdxx49tuTE1rGtMg4OZf1xDi7rWY524A4+5RXZhDA1uRAJYPLZty2Ypmt1TagtjGRgsZtHqh6E+uufEUrzvaFTZxICKopUsrZ5TxR4RcebQJ94bUjWrgYbRca2aIm9pMZimGqWWyRpYqGoAony15fhluMuBESs8qNkGNJtX/SJoSbPdu4i/ypmyKiwUxtEUIEpEyxq8OAfuZ23qBIJS3KlkmrAxE3OYrRCmnDwOvAA5O/trbxjEup4ll8vwkguKp4EMWBGBHC1+ekSnDUL6De+kYGmPdZGY+0SFO1221LIc6oI/4dyQq6K3788z9nC5ovvdZG0jbbVN8yvmJ9bV0/i3FDitVSDIMdJqleJRDN908AmkB/obila7hnzx4d5vnz+d+VK1dw+8YNVEsVqeF379urWBOu6IyB4oYuNzAoZ8Py0pI2sIoNyqQUwcTmSJIVBAl4TTg2fA4175bU+FzYpMKISAXI7UG1VpH6anMzj2SC8QzOZpxMaCPE3M+trS3FDfH9M9qKvx8fHcXg0IDiZKjoX99gQWQUI0PDUiTXm2U5Ki68eRbJaFwRRfze3Xv2ID08osgMnpt58OH7MKIigm6bsVIlsDiYSmkWfHMzyecvrENswwBfV1xNMkMqQN1Xy7LXYc5Zg7U54uIaTePg4SMYHCJwS7cVAUweJFv4o9//T9haX0cum0WUoMAOtSIiLO8L27xDJ00kajFGyqQmMJyUeoW/Z3QSr0E2m1OGeSSZRW5oWJEz4VgC33/xefzOf/ptTO+Zxkd+/GO6pxxbJA84VjgOWGJKNwfBev45/6My3m8muMFnBwZJL0Y/9Q/06x7xWf3Lp/4cU1NT+JnP/yPs3r0bpXIZm66AnKonxm2RmOI95IH2xo0bWCSwEotgbGJczxjz9e/cmVG0zS/+4i/h+IkTup4bm0v49te/irdfeRnhRlNxaSySNvI3KILCyMeWQCtGP63mCwJgGUdAMIdOCWabc+wxE5mZ+BFmnYaCUkPxWRwdG8HJM2ewVSiLUCBR0WA8UhciOQj+pRIx3J67jdn5RTSqLaQiYTxy32EcPTSF8ZEJxEamMHzwFHKDU4iGEupZaYXauHT1DlhGfuHCBZEg//jnflb58aVSFRtbG7LpHjx4ABcvsKNiFHundoGp8by+nXAC596+pXiFkwenkY6F0RVREcLLb5wVMHjowAFcu3od//zn/zk2VldEVHRaLJsjScEDNAk2U38GO20Mp5MCKU8fPowjuycx0t8nBwQVXK1gF4F2V44AxoTouQQJI5ImcQQjcWyVy7h65y5eeO01fO/lV3F3aRndUBi5gWGB6N41NzI6pjn+sY8+ip/56Z9CgjFSbuNIRwWz6GXz1mHDqVwdeGRbhwBKlTrylRIuXr6MM8eOYbx/6P+Ho8IfQUSzOvUn/88IbMZQsRi3VGngN37j3+OF51/E1tYqiltrqNKJ4jbRtj6aosdvsDtdWv3ZHdBGMhzAxCg7QvoxPjqIsf5+DPYPYdT1Igz29yOTSqhbpsNYAanrYgKcQ5GEQBwd4hkxwfm/3sD6Zh4vv/4mfv1LX0J2eBBPPPkZvO+RH0O12sSjH34Mub4h7UcUPZSMoS+bVnyTVEciLgO4eXcBz73wArJ9EYQ6TYwPZLA0P4PJXeOKQjp7/gIGRg+hVKpr/IQ4T4Simtu3tpglTpC3gUvnnwNq8/jUYx9AIjeNawstFCp0SbYwP3cJwAYe+/EPY2G+iHYrh6sXXsLuySCOnXgfltYYJZFEsdKQnT3bl8bsrRn80e/8Ns6/8TLKrSIrxBFsdzGSSeHJD96DPVPjGOijAj7zAuqYAAAgAElEQVSMYrmCIg+9XUZIWUQL9zkkGXj8LxXXkckkcPjgERw8eAjRcArL62u4cXcez7/6msrrL1+/LVfLz/+T/xmv//CHKGys4XOf/jSOHzmCtfUtfOVrX8dzL3wf/UN92Lt/n4q62UVx/PA+HDm8B1P3PIxO327U6wkEWkGkkwlkcgkEg5FeB4OfH7nOcb6ixZyEEedPHtrpAKSDTNnalRrefP0FvH3lZURCJRzcP4Hd05Nau2KpOOKpDJKRIXzn6y/gztVb6NQLyKQCclTEwglsFYpYWF0VUcnejkK5rH1GXyoiEpjryOggSZApDGb7RF5z5xCJp1Am4Z/fxNtXL+HSpbfQ35fBBx+6D1PjQyIqtMcLxBBN9CEYTaLcCmAjX+YChu+98AN88smfQq3dQZ0xF4mEuny4f6Jimv9PooLqW863W6W8PjN/rgEhBvwKiHbRTzz4EggjKSqiIhjG4uoW1taWMTo+pJg6uhYY/dRqWITC4tKC5mGuXeyOElGRy6FSLaHarGr+pzqZBC+vPwEodmhwfBeLJczcuSOAg++H7gs5aBVBaXtKaW3YCyLFKV24MdQaTdTrTe3zKaBuNWyuUucb99bNFlbWFqWa7+8jEcq9n0W59JSDDhyyOEyLk5ufndfcEk/FkMgkEUswBsWEP0ZUtE3w4DokeI1JuvFrdXVN/889HglRfs3NzypWkcWUIhjCfOYyiCW5NzBwb+3qkkU/hRj9REA+LABMp36KjFzkhldse8W0H+M+tk9qbBeNJNBYJbbufOHU6l5lyp8uJ7RTyVpxsI/ScYp4163nwRqJoVzMbM9GsYOo0DnGkSIWaei+X9d+WxDmwTrfQaEziftr3zHAxURj30XMGhBv4iSSjzwfCVB10bkCttRbYApzfjYDR61MWn/tABZPdvA6SpHtnCn+LKbr6+KYLNqCIFVH65scFQ6E1phy4jK9Vxft66/DttjNgC4PAunPffGuew75eyuoNvGcL9S1OCynpFXkUFj7er5vU85aV5Otg+aOVJyJXPcNxKNUN7ewsb4moIhO8LnZeYyN71IE4uWr17C5WUCAYhjn2DV3ANX4dTlfeS18NxQB7wcffBDT09Pak2vf0G3L6cH35iipngDOlL0U//l4Fe+epziMAKaVwfLy6AwmIMs+m66JU53z2nm1vMhV1xOpGBHfTenidvgsq48hHNbenOsywTgBp42GnNx835z7eTY29TSjnMxBJEGjuh1sHGgNabW0JnuHhaKM3FlNJIZz3UgZ7ABfvmfvGOE44v7ekgzqmm+4t+Dra95yMS/8Nd+buansoVD2viOieJ15PzmH89raeTsiESOFGlKEO0W2PRJ0hFoRci/azb13/r5XsMy9E68Fv5cKdZLoxZKB9hqXBj57xT/HqI+OsdJnr7MnxuH6ZXQ/fA+SZe5bvJT1Q3K98K4Jr8z365KEIiJh2LVkBJERTXZe9SptkiVco/iMUqRmhJIFH3ZbTeQy7McrYXllTS5Q9jdxrPMMxzM7hXd0LNCdJzGaK6s23MLOMrof7v2opNphJJzPvcNFjhKNme15Tp9d8WS+LNrItV78uBdeOmW+fUYjdHx5ucaQ+/x2P63nx8BqA5L9vGIkiQl1bY4ygkBOF9els33PiAKYi8PHxjkzjnNUWAeU9sHO5cDPbryZjymySD2Rmc7FpJQLYmBuvuOo4LVkpBfJLH5595qec0c82323IvPtWCdbNfx6LTJEhCsdcE58y4g9//ncGmEkvZEgXE89xiWih2uSWwvcktEjjzwup/VJzyvj2UzwK7eJUhZsHTKi3CWt+Ngn9574968906fPyi86KgxHsfdvXTb2XChpxEXO8Xv9a2ntdi4O7yTUvfYPmuZDH2/o7rMjat4hHHBRjzvXHz8GRJLscEvsJDc05zhRrU5r7r1qfvMXzq07Rri7/Zdbd33aiRc68DV9h4lhfFbKbiaS9zoqeoPlvV/8aF2Bk2nbgBgzaQyfORFtobLCOGOJ+TRoY0KljFP8cwLXZm4HM+2vkJETRlT4B9lP9KZssJ/bK5hxbK8HmRV1JLeH5V33Fge3iSSTqMVPhy6zSHMDpMIbsfk2GRp7aWouqQ5cAfXO96RDps8SdJtqKl144OTkQUWbop6CAW3elCGYIpAaRrVc0d8xo56HWV+axc/GjZDy8alQDxsLz4nZjA22gdNusUsyZ5uF5UTOz8xrbZZRm8x1cGB2ONUB8IdF/jweqCx71VRh5oox9tYmYNnUqWytE9yzhVgbmJ6Sy+6/L37SYs+IApeDaCy3WaIVBUFihosrrd/Oui27W4fAbV2EBa+1ERUtERXcRHz08z+ne+mJCr9x5vuIRkLaEPEQRfUnFfwW2VFBpVyyAm1eb2bFp5IYHR3Te+DrcdKenJoUOM3Pz3tEIuDs629gc20dk1NTch4w+oNjhPEgXPQT6bRAX+XJlsvYKhawtrmBeCqJgb4BMdYE21KJjCnSvP2aCgIqsake2EFUcFwxPohl1ASa6Q6g0kSOilSKofXoqKS2IwU6iYpD+w8o5mlhbhaZPoLoScRiSQwODGFhYRn9/QPauDZbZSzNL+Lsq68hFUvg9OnTivCZmp5GP6NFpEixnFduxHm7GFdTLGxIBcr3a7EOBkaQyGKcBg+HtFGzILCQ38Ke3bt1z+xZbBrrz42eOwQRoKfFs4MwRkbGMbV7D7J9OcRFypiisdMo4pm/+briNaRep7tCkWdBdJi/q2iqpB2c6QqIsrMjhXgyIQCOEC//jp0JqRS7PwLohCLIDIwgGk+hE4wgEksgXy7gN7746wiGA/joxz/RG1dePUNCgoctkkb8eRwfVEATCPFZpASfCZCwu2F9bUVF4yJpmk185c/+TETF537yJ1SGyOJlOmP4c0l+aANZrWBhfk6fb2FxXgTQ6OiogC2quPnMzdydwTf/5lv4whe+gPvve0Dz4szdG3j6K3+C2YsXEWkyJq2OZqCLBkF4Z7+3gk1gcNBee62Ql3J2ZGhIEWHKG6biJ5VUXMxQrg8xqs9LZblnxsZGsW/fXkxMTWFpdQ2X3r6Gc+ffkuq60Q7gxMkTcl/M3LyOyT0Tig+bnVlArZjHYx84g3tOHMBAth/JXXsxcvheRd4wx35yehcCsRC+89xLmJudE8HIr5/6qZ9UUfftW3cQFCEVweTkOC5euIjxoSERFaEuD7wtdMMJnL18U0Th6SN7kIqxpDiMejeIH75+VlFNB/bvw6//63+Drzz1p2jT+cPybFcWz7mBJIUBUl3EQgGc2bsL9544ipN792JiIKcCbJKPdJl16LgIkeRJIdTlODTQpEvSmgBDJC47M2N57i6v4vuvvoJvPvc8bs0tIppMi5CjardQKqN/YEA/d2JsFP/45z6P48ePuV4Rc3qRqOB9Czsnnt/Abh/CAiiU6shXi7hw8SLuP3kSYz2iQtrZHZqod+87tg9y7/4bRugUSlWce+ttfOlL/0H3plhYR73MKKuqPrOAtoYVTb6TqGjTi4H+RAwnD+/Hgb1TNHujlN8S2VupNPSuhodHcO+pU7jnxFFF7ARiSSRTadSaJDSJNccFIvPwoHxdljnWWyiVK3jx5Vfw61/6d8gNDeLDP/4RPPrYR7F7ej/27z8shTjV3YzwmZqe0PzliQr+rFqzje889wNM7p5E32AWoU4bSzN38NLz3wE6FTz+xKNIpGJYWiPBzE4eZtgztzmOWr2tUuRohCqtBmbvvI7F26/i0x//MPrHD+LGchvFagytehsTY334m2/8IT77uY8AgRgKmyFceuuH2DedwrETDzmiIi0yKJKIaO2/fO48vvzb/wG3r11CvV1GEw2EugGMZtL4yUfvx+5dIyIq+jJpuVDYgbC2UcBafkuKeJ78LN6Ge6IO+rIp7D94ELsmp7V3WN8oYJHxT3dmka9VUWHfRiiIfbt3o1GtaU146MEHcebkKZSrDTzz3e/jO889h3SOzql9FmtXq+LU0YM4efQAJk8/gNDAfpQdUZFKxpEeSCLY5RpcNpWrA+A9UeEEk1IXMiKArjIStyxoz5AE6FKBP4Pnv/s0NtZnMNAXwt5949izZxh9fUkko/145YVzuH31LiqFMlLxBHK5DDpoYWFpESurGwiwRyeWQJLERiKG/r64IgwJ7mWS/C8l8J/rBa0J/P6F1XXcuTuD1dUlNOtljA4N4KF7T2F8bFDPqBzDEbp/0ppzyk2WmVdFTp69cBkPf/CjqHDsBiBwnG41A1coLGEUU0WfNZXJYLOwqbWUMaQGDLioGZXPWgSCj36iWvzdRMXI2IC6V/gaLKPpkC3mXmBpQWsT1xVPVFCEQKKiTiK8r09EBWOgGD/C7+P7CwaiWmPu3p1BktcmFNK1IiAiosLFfPiCbAL+Ko5kv5h6swjssHCe64jFDlFUqv1/q6VryvXFop8IUtCB4RXSDvxzmcyeqFiYnTfXbDIq0QedFVQ8kvhgDwkP5bYX8Fna7yQqOD95RwWvMa8NxQ4s1yawxZicVJZikpTUrRyn61fYFcX7HEWUhdoREpRGIpgTmHFQ7owjh6ypM/1ZRNFGLhtf7g+RBXa28VER5pY2YF7loA4w5FzqVZmmEHVxtVRAusJklTfTXepypdX1IZDDCCRPoEh85ctJXUwMzwFWoukjDg2QVzQSFZfuZ+ocs4M4M7WlnQvsvOMAe6fO1tnKnZ0M4PHfZ7/mz1MMEyN3uc917hGeQUQwUOwkoMx1Uwjvs3NGry/Pxbpa7I8RFRYlZX0nAgVZ7i5VdlIRM/w76x+ga4LxxHaRuGfm9ykOJWqxL/7PjSTadqX4/HGL0HCFzd694WNanMsnELCiainO5QK0s5ZigqoVOcdWlpdQLZX0men65lxQKpZRrNS0LlVrDaSyWWxuMRLJ1meen8z9HhIpyL02o+rYE8MeLyrbGWE2NDSEiV0TmBgfkxBC57aOlSMLlHckkN0rVxDr5NKK1dL52Ap6ORY0PrVfb1p0liNdPEklcM8JykjG6j26ThD+XaFg5dISvznEk2IUXg8SDdafZ+OOz0QixrnIeiCU5884pwgB+5qIHV5LzjNcM8zhxhQFP04cCK2ODNd/I7W2YRIijERsmSNIAivFkYWMOLHHoKfGl3is1XLzo7k6TFjVUfSjIg0VnUqBin0vQXZzg9BRaq44jX2pmXmOTyjqimOewh6KHiwKiGukcygxCYLguEhx66wxXMHOzQKeFZFDFwrxFeuA0B5MPV6MwmVMVl0/O5NOu7J4i1zj+7Rn2eXSO/GYd6wL3+Cz6MRfEtS48xbPH5zzPSireDwJIhkfZNdcZJUDT/meKR5iN0W70UAua+QSz1BDI2Noge5W9lCyY4PrJFMriLFYLKFXvpv7ahtH4nNhLjZHJkTsfVA8auSazdn+y+6rmyfVp2EFw96BYMSrCV+9a4z3QMXOxDIoIuQ1kxDU5hoP5Htcw9wYrqOUgkyHh/F7FT/uop6M3CBh2e7NVYq+BjGond0DNgeKJHWR4po3HR6jiDBmaLr55t0EgO+1sOfaekv4b/lcKg0kxDForhOLlbOkjd4aILcTo719IbTrPt2BBxlRsJ2U4vd5vQ4j3TPXheKExZ7w1jrlEjrgRMbWccJ4SbsP1i1lzq6eC8uJoI2osOfZY3re0aZ0DxeZxWfi1R1l2g99qthbj7xbyTscjKjg5zZRhr1X64qxOdHe1871wc5jlg6xM7bXruM2Fqef7TssXBSfXFn17UJzc45Z1wT/vU+C0bwaNsegYauOTGAvJyM4iS2R2JXbx/A0YV90PXEOZR9HtYoUY9DVkWRRc5wDNY4dOedfV+/9PUfFjxZI/96nAU5nuRharBO/PGAvNQ2V886t4CdyUxNwo85NKsU+toh4BZC3s9nD6nLunBJDNlG3YbQkP9tsexLCawl66hxueF0Gn+W0W9acd2hwQZKayGfJ0Rrn2OWe+sdZn32+qrGRZkn2C5KUJW6C4eHFrPIhIxciBOK5YQybNTfKCBEWKpkNzBZA5vuau0NxMlLWsTPCNnLG4LL82qmItGJtK7Fsc9Zyh2NTihCI17V0Bw9Nqk6dJMszNwNd22R5FYux+px8bZLeybJqgdamvKliZ2UpBqxcyqyklm/HCU9Zf+7wYXZ9s6J5woqHB/69lQfapl6WPbLsUrI01aWgHOQ2eymokmig1mSRVxOP/szne0SF1Gs7irh5CCXAzwWOlnIq/bSxVDE5gZGiyApm4XNDp9JmKuhjURFHBJQJEHuVCVXyF86ew+bKOqZ2T2Pv/v0CNngI3X/ooHJASVQQINJmngfncAir62vYLOZRrzKGzK4PPzMBGh7a3I5HY3Jn9BMjGUQGNaoosaAbQctNVRZj0BSRKslr6PtYQMwFqVGrY3p6SkV7t25d0zjfu/cg+nODyOfLSKeyOpxX6wUszs3jtZdeVhTG6VOnVdBHYLhvkJttezYJsFcrZW2OTZ0lo4JzM5lKj2oHgvEcP7zHxWIBm+urel+HDx3U+OWN53Mit4xXWPD/uWFsMvaqK+X0+PgkhkfG0dc/iJgKPkmCtVEpFfCD51/ACkH8gJUbK2c8bqXpXmXEOYCqM8ZAsWeBP5NEjcjBQMhdww5awTBGJqYFPDIGJkRCIxbCzTs38cLLP8DhI0eV0U1QiYc/Aj9U+VNxmi8Ude/82OC4ovuGgAhBAI6VleVlrK4sa1xVGc9VLuGF734HR44exccf/4TIDZZp8z9uKng4paKTJAGJtHqlguvXrykmgBuJXlF7IICbN2/h2We/hV/+5V9W7jwhlPMX3sBXn/pDbN65gxSfx3oVjSAj9mwjZM+GqU5yuQFFP5Ee0gGAETLFUs8SzXs8PTWCaBDIsvujA+yenMKpE8dx5OgRxDMZvH3jOl4/+5by3C9ceBuhWBJPfOYz2Ds1iRe+8y3E0lHEkmlcPH8ZMzeu47EP3YMzx/dhIN2P8PAEhg6dQSwzjmAohr7BPrQCHbzx2gVtnKmCn5ubw+OPP66D3cLCIg4ePqjrzjLtC+cvYtfIEPZM7kKwwwNgB51wHG9euqGy3vuOHUAySvIghEYwjJffOK/ujI2tAv6PX/vfsDBzE2jUEOgSDDd1J11AHMsRzX0tjA8O4NHTh3DiwB5MDQ6g37lnIvGk3BJUu4UDjMpKkIoXeRjkQZqAQMSRyN0ASuUaVjbzuHrnDr753Pfx7ZdewWa5ir7+AQyNjKJYqiAcjQmwJ6DwiY99FE98+gm5arhecOyNjAyKqAiZHcAprnyYk23288Ua8uUizl84jwfPnMHYwLC52PSsei2pKcDe+WWOKQcnOQUafyavKuORuvizp76KL3/5z7C6vIJSYQ3NakGOG0bWKVKN6i1+fqe45NzNf50IBXB83zQ+/uH34+DeSYTDjLKjG6KI1fVN3Lk7i8JWHlNjI3jwzAmcOHIIyVQ/RscmpIrnM7G8ton1zS1Fy9SZaBwMinzlGL58/Sb+9Re/hGx/Hx750Afws//Dz2mu63RCGB+bdAfidUwx9inQ7REVhWIJ585fQrZ/AKMTE1grbOLQnn1YW1jAd599Breun8WhQ8P48KM/hmK9D2vrJcU8haNJxf7Uqk0UihUEA8y0rqBamcGbP/gaPvXjH8SufSdxex3IV0PoNIOYHB3H5UsvYatwE594/GOYnyviwps/xKF9gzh67CEsrrbR7CRRrjSRSCcQi4bw6osv4su//VtYXbyDFmqoterqrBnJZPDTH3kAk6ODGOzLYHi4H319/QhGYup2WVnfQH6rJJUjo6IajQqCwTaymRQOHDmEgcEhOQ6qlQZW17cwM7+AKsULEUZR2Bjk3FkuVhRLmU5msJEv4flX3sTfPPtNhOMR7Dt0ADMzt6TuvO/UUdxz4ggmjt2DKJ0ntTgC7ZDIlnR/Auy596ChwESu3w508XGHVOwXyyVUy1WUqxUHuKUMuK13sbGyhna7gquXX8Xayk2kE8C+qV3Yv2c35mcXcOn8ZayvbiGEqJTx3RB7DWaR32IxeQ6xKMmJlIiqbMqKlQeHBtV9w5hEugvp6OH+g0TE+Utv42+/RbKqhYE+kofDOHPmBEaGWQ4eVe48iYpQJIl2IIpqvY1KvSVH1/WZJRw/cz/KtQa4SHEvYUWcYZFHXPsZY0egikKDjcKm5iuuJV6t7PsGfEeFyrRJzO8gKpZWt7CytoSRkQEEg13tOdhPIcyi3cbS0oLWF/5HooLrUEZERVH7JwKjdM1xnuNnzuWyGtMsoidwSqIinc4IbOXaJpUz92FOnU+shOCFd1Q02Euhgk/u+7poM3HQUksRlECIisi23nOz3hBRQRUu57ed4LgnanY6KjxREU1EkCIxlzCnpO+o4P9TSCRHpcDzdxIVfM8ESn3kzcrqkq4ngTO6KuioSKSTAnu5dnOGXH17Ufs5XvuIYh692tKAGlMiG+jAGEqvMvfRRwLRfUE4SQudcywSwu/DDSw1cFxgci/2SM0+BlS419KZyfUe8HrxvujLxevQ+eYjHXZKPAXsyclh2eveIaD4UN0rr/i17gIBsT3XhKlDvRvBC7WMJDCA21Sb/szGva3LTucZxfXVmVPEzkEUYZA0sGghU/MqDtZFZ/pOAN4HI3ssb90TFQJBHfCr8wG70uIWKSR3iQOg+ZpSxLt9p4AuKrOpSnXl1hYlZWChV/cTqPWOCQ/+2nUh+L79b+3aGwDF9+9dHXzepcB3kTy8F+acttbZRDyKxbk5jde9hw6ivLmOZDaHwuYmLr99FasbW1KXJ1IZVOtNuV5PnjqtuD2KhF555WWsrq3ife97BJPT01heXMJrr77Wi2Dk2xKojC4+9cnHUSoXLWKN3XEOmPYxzHxWfYm5ZZPbeLJ5yM6a3r3pY4YlO3TKbA/I8VoTbOdnFxDriCsPmm53HZqDRcCrI9l8P49ICtebQUKEY4OiPLq4SV6rG8htWxity72wJ090NnX337tgeNYjwK8zvgp77fOop40ONHffmRBARFIRUfy10gTMQeFV6vxelUhLiMd9oj2Xfh/Ge805QEAfY6aDJMpYOk18wX6uxqUrcvb4B+ddnpN4JvRgqZ7HHf0EitMiwRK2+U4xPt6R7uYL3gcDNi2WiveuVqUAzzrnOO55TuE49MI4D0ry/vv4Gq/mtufL5hNF0DgS0M60Nk948lXXSGPHYrI5r2hO6MV9GdGgHPxwUI6KvkxKz+XS8hpiiTQCjD6KWKkxyRquuzoHU/BDiZkjG3aKEO01bQ7yCQ68vATfFS1Nu7wj/g1zsG4l67JxY805/fw4NTzIA8mGe/ifYZ02llLh3V7cg9rzb2crqfOdaNJehw4dA5R9kofGEsvJmT7hItWMGCARyIgrkmAcT0ZuSTjmHE0cZyQjOd8Z/hWQ49mKs80d1Lufbo7j+/Lxb7pWVNo7q1s8wUQMi2FTjyjxNEfw8dqLoHFOG5+44fco/y977x0l93VeCd7KuapzBtDdyCAIkiBBSYwiRYlKHgdZ8jiN7fV6HWbsObMe27Nej8MZT/CMvE5HchhbGnlkWVmySAVKogKVKIokQAIEQABE7Ebn7urKufbc+71X3ZDp2bN/2oct4aDZ6Kr6hfd773vfTbw4XvHnycUe5PX3hcdH0EhrrMv5sDwqsxNjz4DWZeoLiABLZYypRUQJdtZuvf6bA5dtTJobi4ais4uzUHtbr9Rkd2QB/TeAZx7r6217jr3JiIZeveTHgAdodC42HfbWOFv/bM63120p8vhzrzzz45H9Kd8P8eCDVyV5VZcHhfy6Zj0+W4e3EwV4DmaPZefl8698P9Dv4Kwe2crn4c9Zu3FcmFKtqhrWPz/sSVpelY1RCUlUQzlV0CtARW/MvPLNP5ErcChprJTvboSoaHTSQz1oblK3R8HLTU3FYAqGbYFfUmAY8z7AhY5lBL3oxFKzIlwyOaLEDg3XhKL/2yKncBzZQtnEYq+xT9dD6n5PExsb/U5Wtv22eLsp9oncqtTz7PPotrwu3bl5xYC/Gr5YELLMU5IAxCYESfVcgJLJ7HjcJvmW4kEhUjbB91BUJyFUgeaBEXfcZLlb8WIsJc+M8ROfX3x7CD1Njsm8bjDU2+S2WiS0sbAwo60JlhsCL/0z8MMvTAZfayq3osndB3n9KT/DACux6p0nJ/9bSL4C8WxD5TcVktwFurJ44h9aZjVadSlDyBZnEfe6H/rhnvWTv19eRcONNNURtLrhJoGAhVimLEgYyE1pbpeBpJuYn5vvsfFptcTXseBh454NDdlTVKp48fQZFDc2sHN6GtOzexSMyoVzdGJcC0Amm5NVAjc82uQnEjp2FuQEQ9gcZjCwId4xZNNZsRW9z678PgEVIwIipDixrA3aGZj0j4t7EBkqA0IsjmiBUBXgsmNqCpv5PObm5i0TomN2X5FwDMNDY4hFE0jF07IFanVKWLp+HSefex5D/f3Yv3evmu283+GIyaVNxmsMDwE5DFrXWGyrKaDNpJqUVpjp+NodFAp5LBAAqlSwY+eUfMEtjNJYlqaaokLKilqBNNWWCq9cblC5C/2Dw0hnclZkxoJSqjDz4fh3voOla1cRIiAXMa9S2U+w4CeLJkq1EUGnmJhy3PTQ/94CvMzXkveC/uI79x5EMBpBsVgVc5JB0dFkDPMrS1hYXlEzRwHrxSImJicFRBCcLJYYpEZZd0zAozIsymWNq2jELJIWF5Zw+fJVPcfciHNMfOULn8O+vXvw8BvfhIHBAXQdY4pBp0EX7MoirlkzhvFLF85jZWlRzLOR0VEpsHie/Pnjj38Zv/ivfhFTU5PIpZN47tmn8KmP/i0qK0uIB4PYLJYQYfigy20hAGD3ClJPcFx0w2FsslnmiueJiZ0q9plbcPuRw1hamFNhjUYTu6d24tXHjuHwrUcQjsdx4dIlnDp9FotLzCugZD+Om26+WYaKcKoAACAASURBVKBXo1pGgEV3IIhnv/MMvvT5z+O1d92GfbMTmBwbQTfbh9F9t2Jw6iDqnTAWVpfR6jYQ6sRkl3L12jWcPHEC9959D2Z3z2pyTyRSYIN5x45RHD/+PCZGhjC7YwcndI2rdiiC46fP6Tk9etMBhWnTCqcVCuHkmZfQaLTx4b/9W3z0wx9Co1xAt2nB9Sq6u1SUWSg0f0bbqCMHZ3Fs3w7smZzAUCatQG02r2gRxj8cU7Y5ozUBfdNDAilCHGcKBQwLzOPnbhbLWFpbw5PHj+Mjn3kMJy9cQjiewODIKCKRuJiRw4P8PoiZXRP46f/tpzG7e0abDGaXDA4xvyQgyxUvsXZieltvmWGzWUKxUsGJE8/izttuw+TYuBXZYtXyb7OFEfDvZM9WjHPD05aShL9rLCwtCco9KFdqeOfv/zG+8qUnkN9YQ6WUR0OhvLTkgxqfXTK5u0EEu0EEwoL7lbVDFcprbjuCm/btRqtVl30X5+3+4TEpkbhhZZZCvbSJkb4UDu/fi/HhKezcNStw5/LVORw/9QLm56+j1mwglkkjlUnJOoZA7+J6CX/+nvci2ZfB7a+6A9/3/d+He+6+H7U6VTYBrK3npQBSmCTX1QCUP3Tq1EkUNku45757cPHKdezaM4sw1TflGk585yksXDuFTosB3Dncfux1WF2vYKPQRKVBD2h6D5PNTJZsBrVmFc3qAr71pQ/gTa97DXYfvB3X1sNYK1vux8jgKCqlVXz1qx/HQw/ejVgkjie/+SUc2r8Dew8cw8JyB5UGGzNtBbKHgl088fnH8P73/hk2N5Y0NpmlQRb7SDaJH3n4bowPZDHYl8PQIK0Lc0gkqSQIoNqooVKpoVKsClQqFDaQSIRl17ZzdhcymRwigZiAbgLn6xubWM9vIBTtirHOPAUqR7rdIJIc66Ewllfz+PKTz+KTj34a3VAA07tnMT9/BfWKARVHb96P0X1HkJ68CYVqDJ12UEqUgYEMajWC3FWx8rcDFawPuI5w7eQcS9Yt11xubNm4T2UJztLKKIiV62uY2bULoXATF86dxKlnn0JhdRmDfWn0ZRM4/+JpVAtlhUkzYDYY7uDq3DVsbJbQbAXRqJGgkMDYUB+mxvs1X+7asVPz786du3R8/X19ApY5Nk+ePo2Xzp1DJp1CpZhHXy6L/ftn0defMbIJ67AQmbQxNDoBjTX+HYymsVxsYsf0IWyWqwjFGGJqAZNkcvOact2n93yx4ICKzTUxUWkx6usoNZPsybW1mw11Wnb6rLVAGEureSwvL2KYYffBrtZGqoe4DHN9W1leFtuY9k9Ugi5ev666hIqKdruBZCaj+iIUMSXs8MgQ6rWmAAYq7a5cviTmHddO1oEEiwmWWZgpQQHzZ6f3Pf+bFm3Wa2d9ToUVVZjWFCJgqeZ3p6MwbRIeqM6LyMvccsd8Dd5rDEltQQVnU4A1QQ5aPjFMW0BFL6OCLN6WrJ98tgEvAi0S+cWMCrGcZW9lSmCqHKVScUAFmeqJVELXR0riYADrZ5dEcCA4JCCCIFEvf8GsIThfCgDw1ku9fY5ZfPmGv+od13z0rFbeXzVktvlX257EGoSUkvHfrPlo4bY+LNQqbJuj/X7D2zCxrmY9ab7ePpdvC5DQ+JVimcx8IyN5ZQT/tjBWAxt4LN4uotfAsVaN6jWfc8ffs9/fyt4wYlnIFKO0cSEYEecYNRsVP+Z5nMrxc7l1JBT5RpNnr1qoMOteI5f554Q1JBvkVC2pQeP3UG6fpPviQBcev66JY//662aNni3lh78m2mf11BzOIoTNwEik1/jl3tHvrfzew/ZnRrayRps1W0WUcqrka5cv4dJLL2F0ZNjskEJmm1OpNbFeKIpcwfw0qhkJ4E5OTMk+NBwK4NKlS7p/tJ5lTcj9wuVLVwQu83s2o9jwJPh2/733OFU8AYmGxjv3kXIdIDs8YLY/vCbcZ0pZoqB2V5NTecM5R5kVRqYzOySurQYeWVMuYEQvMc8N+JIKQyoyAphml6xGrlMF8HdFoqN9cL2umoRj0yt/tR9y1lA+C8EHp28P06aVq1jx3E96tr1Tf3C8cWzJesuBNH6/6sezNee6vUwI7v5ZtPH4OVeTYOity/hs0G6M50/QU9ckGNLcbfaqRtDzY9xbFPl5gNeb7yeraMdylurHXVsParDeVni5t4ZjMPo2Oxg13jXXWI4Mn61eSLqyikwpYGooU65z/rI5x+3LXZ/CGshefWJ2V7ZOGwjIdVO5kfL8N+KixhCfA/nvm1JFjH1Zctm1McKkuVHIPppzYLOOFC1sR0alKFpb20Ay249uIIIAx5XbE5KMw7n/hnyPnm2RW2NcPoQauM7eSXtRjT9T1Vt/x+Y5m6+Ya2MZP2ZZzbHvADmnSOC+lveSr1cmjRtXmpJdoLc/N14DUyrYc2AACD/H+lfcy/psCTXTSR5xRB5jc1ozXuBgr2/URaG4qZqO78V50TJiDLggEZGkBnuOCdiz/uZ4MAKrB7rMysfZCG3LONVx0U5Viic7boWG+96VzkIpEfblsuYIVBjgY9fWg+gaKy7XxwMWBr47sqrUagaS+d6WZWmYOlE5tu5aeZKrjTf7cD4nvnbQtXJgugaI+/Lrhf9vm2Psdf57zsfPfG4LqLj94Q1rVTmwT4oMp3o0YJXH9Q8rzXtgiHNZMUB3i9C7tR7Yd9se395x+zVo+9qx/XVbAL09d7xPAlRl22jnr/Xqu8K1t3+Y3AH8abiD8Ioxb6lvfbotFY9/gc7xFaDihvv1yn/8E7gCBxPGbHbzW09qaYitTYq+SaJnJ+gCveS7asU0JzBNeK2WilDKKE2KapOxAgYpeWXDTnLaSO97FR9ucvPop0elPetfLCInx/NKCHm8OTsnyu4kg3aAyrb5ugfAeKDFpHqOjeEtfFzIlWdam/TYmEd+8bSzcAxWNp6cHRN/LoTTofoqjCQ3NPaUGD2Sm7ugPVdkswHqGSkCAJR2bai1UH3HmuJ7yCrKWWDZpG/yaXkIu9wJj8CTfc4iSk33cESLOyc9L/8WO8VtULhYcQLlxs7ifTwjx21WXXifl6J7xJvHS7ZMkd7ULCIYuqzgIpOnctGq1ivGYgjSL72hBdysn7aACi9P5vGYFNSYYRw3LDw69P53zBJu+jkGGDLN42SmQX5jHesKq2ZjgD6XlR5bik1qf60219fRrtewc3oW0zN7FQLW7DQxOj6ia9Noc1MZU2jewMCgmow8JtlduHwR5kWUyiUV97wOvM/JeLLHAOP15TXhRoTPDtn1bFqzgcuEWz4XwU4AmVSGvVGpYQqbm8qlmN41rfv13IkTuH59DiOjDI7eiZWlFdTKbBAMYWx4HM1mDc12QR79ZCj157JicBOYMMWHlxw6th8542zMRRmsa6oWlRoma3KWCAx4NO42mbFslL1w+gU1Jg4cOIhdu6YQj5o/peYIl3nA54nFdL1m2RX0yd41PYvxqR3o7x9SkR0kIEGwIRJBfm0Vp597FisLcwg0a7I2oUyUCopEPI0omS7cDLAZEQzL1kMNF9dU4DjbWN9AIjOI3YdvRSAelZqgW2vqGgSiIQSTcawVigKYeO+YxcDxzbwAFu+drsWJ8nqwycH7RWuypeUlLM1f0LjdWNtEqVLD0NAY0qmMNj6f+OD7MTExhu/7/rdhaHREDU8GftMGiL78yvZoNbGZ39DfZNGdPn1a+SrcrHJMpxMpARVfevyr+MV/+YsY6M8hlQirgfeFRz6OyibHcRj5YgWJdA6VOgOjmXuRlvSawas8+pGRMWQy/Wi3q+i0aggF48jmhhGOxxCMdDA2MIiygtorqBQKGE5mcMfR23DLHbchkcliZXVNSodLL13U+Y6NjGF8bExsN55XgMBLOIK5K1fw7j/5IxzcPY3pHWPYtXMYgUwSU4fuQHb8AMqdOK5dn0OhvA7UQ2iHAlhcWcaVCxdx36vvwoFDB7FZq4jdXdgsYnpmEidOPI/h/gEc2rdX4AIbZp1IEMdPnUGlVMOxI0cQj4VkfdUMBnDxygKef/Y43vUH78S1i+dlb6P5kOACG/KdCrqBNoKdIKJdYGasD3fcshv7JkYxNTyq4GeGxZMhw+cwEucznjLWlzZrZhPCzQt9pskS4zXg8+tDXzcLmzh77jw+8tgX8aVvP41Ko41kOovh0UmUyzUko0n09dNCLIAffvs7cMexOwQ2BaNhNee5IRbA2myoOGVzjqw8zrmczxaW1zUmL5w/j92z07KRMhVjQDZFZF4ZuMgGFjc4FvZIpg6feY5hUzpZZWuMU9oEbeK9730PLp4/j/zGquaMpoBOKgE439YRYKO2k+AWEcEoJe4NgWV7dk5h7/Qu0MH66rV5rBc2sVEqY2BwGAf2zmJ0MIexvgwaxQ0E2g3ccnAf9s7ux9SOWcwtreLi/AKuLixiY7OAeDKOkbEJDA5mMNDHxmMSX/zKU/j9d/0ZEn1pHL7tMB584H4cO/YqgWYEa0PhpCz8AiGuhZx76lhdWUC1XNQ8yZBmNudjmUFlfATaQZQ3N3Dl4nHM7Ezhya8/hte99m7M7L4Zpy+s4OJcHqFwGtlcv1hxwXAcjXYLm2uXcfwbH8P9dx/CLbfdjaXNNJZLATTbAQyPjKJeKePS+ZMo5xdw952H8e1vfxE3Hd6DXXvuwNJqAIUyg+46GMikEGi38OjHPoQPf+R/oFLNix1ItRnZ78MDcfzUWx7EcC6FYdrO9RMYzyGRoPougGqzLL/0hbllAcXMGhkcyGJichQ7pqeR7etHs0pGaRyRIBuGDdTqFVQbFbSo4ozT2iwrsJcZF81qBasbBXz128fxkb97BO1gGGM7JrG2uohWdRN33noIt9y8G8PThzC46zbka1HUWgHEExEBiZVK3Sw6CIy6GpCNKQWT0n6rXhf4y/WNm0UDKmpIZ2ixxLWnKxu9KQcSV8pFXL10ERtLC5i/dgWl/CqK68voUh3VaSFHJUcyiqWNJcyvrGNprYpCoSE25c2HZnDTvl0YHx3D1Ni45RmFIyjk81ofOLfQI7pUKQucIAHg+sIcaGO1c2pMOSe0qVP/PUi7TDYXG8o66QTDQDSBUHIU2dwMVvMlRGJdJNIMmzZffhFPWl2BkszjoDpgLc/8LFO9Cuh3jGQrOIyFzw28/1v1sQOPlpcWMNw/KHWhrC87Lbo/yYJkbZ1rQBTDQ0MobRZw+dIl5b/Ua2Wt3emcZTbQRonr8PjEKPFedNsBbG4WcPH8BREW+B4ELDO5DJouO0wNHkdgCIWNDNRssFltoZDdVgcthnrLotLqPzXoux0sLy+Indzfn3MNLavxxBB0rGeucVL5Msaq3cHc1Wuq4+JJZlSkLExbFoVGOGA94S0aPFmGpAO+39raulmrKn+C4FcQG6sr+myGE8v7PRKUipEKEgJxVDCvn16ULR/3FyGGaW8DKtgE5rwvprCbO716gteLzSQpBHhHaa/EBpojIHmwjrfXB27q95za3BOi2myWubreWzSZ5YddZ++bbQ0herybok/1ulNiay/miEoiOrHWdpl75VJZ11zsY6dy0nV3TTZf73qmtvYJjthlKnUHMETNf58rhhrIjs3JMcFajcG+VAbLL51gAZvSqsNMfcvP5jjcIp0ZeczYyWZD5Bsv3nLL7+nMx30rZ0/BuVzTtvuh92w6DOjgvet1bnoNHPtMv+bZ91b/+uvgm7e+GUfmN5n/1gj1oIaRe2R35pq9HMOy/JJNalD2c1xHr1y6JNuxarmMVDqrea/ZBpbW1tEJBJEbHMb6ZlEALwkwfD/aw3EvoByTEEOcm7I7JcBo7H4PPrWVofXwGx5yZDWzbiVYwuYyX2ONWrMUMxtilyMocpjt4XsOB2xaO7DImt+OoOTGlncFsIaYgVh+r2/7fWc17Nj4tpc3VajAB9VOZo/H4+E1JfDCcU4ww/vmsyHN+2dggylkenbDbt/PMco9LolbaiT3FApezbFlw+L3gwLuGKwei2locO+izAXO7xUbvxzXCuf2SiJHcFHT2qkJtCyI7WxNco1X7qGd5ZP1FFgrGuGQwFIqnbKAZwdIcuyoUc7nkE1JAiY+k8z1RXogiwcHnXOBGtiywHEuDzp3Azm9tbV6Mb3gbwOtROTsmsUO5y67ZqYurFYs39NAKOewwHmP85kjFfp53vovBnzZDd7y0WfdlYiGUS7kcdstt+AUM+gKJQyOjMsylrWyPctmW81xRoKVqVK8nbgpPPgZ6nPwOXAse1tbm1KeGNhohyCmuFdJCPwyMM6r+NhzsXuyldEpgNMBNt6WUE10AZcGylq+5nY1h507a2q/z/RzCmsfZWS6Zr2U0T6LyI6yp2Zivcb/eZcJ39D3/QyObakQ1McyGzqtBVI3OlWEGxeauxwhVJlJbo5zomw3txGUtNwZAzb8ddtSPxkg6+Zi++ee1dNWM92eZ7vetp/wQJmBxGax5oRI2z7P994IsPtAegM7dfwMu/Y9Kwes+/HI++2t63oKAAfW2Bx1I1Dx7DZFxdEeUGHHaeubuQ3YM2i5rrYqfPeXs1i0C2FD3YVa937Tqy+2/c7LvE1PGW+jYOv9dO5ekemAnR5BzVntyeatN6dsA1WcgkTtQTcn22fbzd0CTbbAnq2f+7HgQJxXgIqXHQGv/PAf8RU4mIzdAB2aDNEmPE64KpYUBmhWIyy2bEKwxZgPHgsPIevbgnJs8bXGsykNfAjOtrBu57Voi4499vYexiwQYrz9WXYTSy9YSaHUhoL7Cd2/S+8hd7IoP6lou6DZYGvx96CHZxd4X0UL9HJBeozGZKBzICBpq1hlLGQdim8yW2OuGRPAJHHyRnZMASNfbfkkejaHfpGsdSfh3i5P8+oKj6TaAmDAjdgILkDMS5r5Gb544fvoXvliU4uk+fJ5ifZ21JiZAFuh6FpXe4wavidfI/9PhXF1kEwxjJg2ETUVHCxIVfByg8X/MRyuUZP9QLPNn9sG94G3/1CPJeHHhfcVNdYOCwQLeNSG1m2geN5s+HFcMUiaLE4WjmxaNFt1JFNx+fGz+OPGmqqLa9euYWVhAa3tQAUVIe0mDpHBnUljeS0vSSdfw9eKtUjWDS1+FOpMyWddGzZuFir0rC1XtdkxkMQ8I/XaDMO0gfz6mho6STaancfsFlDB+9dEfmNDxRBzNhjSt3B9QVkl9UZJoc3xcBRLCwvottqYHJ8wZUOH7B6GAUbl8SxAyrGrmNFgxZs1i6zIMEYV7aYIFMkcxmdJORsB3YMAN611bWbJhjx37kXZJU1P78DBA3vUmPJAoJquZGUzjLdtYfYMWR0aHsOumVkMDtLHP4FOMCAbKPqu0gIlv7aMc6eeE1jRrhfFNE/Q4iOeQoT2XlSF0IYnaI0Gea9K+mu5Kqsrq0hmh3DTHa9BKMkNYBk1bgwJhqQT6MYiUg3kNwsCcq5eu6pz4qYllc4gEks6qNEyRziO2Yjm2E3HjeG+vLwqJjjPlWGttAj61Mc/jomJCbztB9+hjBNu2Qg80ZKFBSjHK9UznCt5bwhUKOA9n8fCwnXdq/GxcVw4dx5f/vIT+LV/+yvYtWsnauUNfO3xx/DNL31OagHep1K5jlgqi81SXs8igYoOny1u8qpVzMzMYHZqFwYHUkglyHrhRiAsS6NIPIBus4EqNy4ECCsVBKsNHNy7FzcfvRV9wyNiAHKcLy8tC0jhsaWTli/AsR6XdUhUx/6Hf/Df0G1UsXf3TuyZmUAnGUVkcBLB9A5sNiKYX7qOQnENI33jqHXaWM1voFOt41VH75AiaY3nFIpifWMDe/bM4szZs5jZsROToyMI0cc0EkIgFsOJM2dQLdVw64FDakA1qCpi0GsTeOTjH8EjH/sw6uUCWo4NRxY9O2LNdgXdYBuBdgCpYBhH9k7i0J4J7BkbwsTQCHL0tE8kTaVDO7E47cQ4jm28828yI/nvbJIHyOhltooDTs0OrYhrc3P43NefxCc+/zjml1cRjCUwNj5Ffpwae9bACygb4Hve8lYUSkXUWg3lczDnhl6/jWpd6yzHNMcVn7lKrYbFpTU1fQqbG2KWk6mu34tENLf5wpf/LWaqY4zyHjdaLWTSGT2HspdzjYlUuh+nT5/DI5/6JJYWrqNYXEe9WhVQoXOTzUVDQEUIlMLTSqWJaLiB0f4cDu/fg/HBQRQ385i7vohWMIi5xWWpCh567f1IRILoVovIUv1SK+PmQ/tx65FbMDA0hnNXF3B1cRXPvXgBV6/OiYE9PjGOwwdmML1jFLncEJ45+RJ+9bd+B9FMAgcOH8DrHnoAhw7chMHhUZRLFcQSGeWdcO7kZLWxsYpdu3ZofSzmSxgbm0B/3xCq7S7qDVpYAesrSzh3+ilMjSVw9tRTyK9dwg/9yI8jEOvH0ho3bENoNshgBToh2kW2MHflBZx+5lHcfmQKd93zEPL1AVzPs2kcEAjZqFVRXF/Ei6eexvRkPzY2LuHwkb3YOXMUi2tB1GoxPU+D2QxalTI+8jfvw6Of+RBq9QKaDbPFYxN9ZCCOn3z4tRjpy6A/m1bQsykqslJJbJQ2sLCwhIsXLwu8TacSGOjPKnSZViEEzitFNhnhQp65DtYkIwrK9jApWyPzsG8JYFnNb+ILX3sSH/zE36khPzI5gVJxHdXNZTx4z504sHcC/VMHMDxzO0rtJKpNgl4RTI4Oo95oa+7nemaBosYK5FzXZNO+UlFDhGuXQHna0dXrSGU4lmyzRhs42jBy3eC/EwBPsCFcKWv+X5y7gisXXkStXFQg+thAEq1AHdeXlrFZbqNcomVCGWOjfRjtz6I/m8NAX59lELA5G6AVXk7ZFZFoSD7v3HRzHl5ZW1aNNjjYr9wizmcdBNVUrDdaqNBWksGhkRiCyTTGdt6My9fKCEaSSOViiCfMGoKNArMHCUqlSkUFwcfV/KoYocpQ64UnW81MUNFCPLlGG2DhgYqV9U0sLS5guG9AwdBqmjCnhw3MVhPra2tqUA0PDEktd/Gll5DNZFGrldXIyvTlrNZIxUWbGR0dFkEg2A1jfX1DihLOA1QksngjqNIOmAJGSkvV4STOWG3/ckCF3+V7Bjz/Xl5Z0D3MZtNq5rOuYy0nhieb/15RLHa8KcE8UBGLR5HIpqSsEHu02e4BFTwGX+tyYY5FzFaIQAXrLDKXeT78PQMqCP5YTRCNMtCd61ZKhAiiuBtnlgRU8J4pj8KNFTWVpCYxwg8rI1kYOTKKBSabFUuvoa7unbNWkM+4KYu9mlsNd1ffeyaq5SRZE0V2JAJjLA/Ndxt8m8HqXrNa8o012/MEBRTwQlJRInJOtWZ2RwQKHJNfGQpuX8Fnz6sW1Njn2OI1Yc3AxpBr0Ik45Cxg1SBXc9LyDHyDm5/bU5I72wqzwzC2ul7nGt/MaaGViu+iiGUrSx0GM7tmkJpfpqJX81I+74545TI2vJ2KgDun9OXnyEbXMfptz2Y+836vxz2XFHfO/93scKwRyrnJW+V6IIbHKXWG2+P6997uR25e6dY45xnQQpV5EufOnEUhvyGggu/DhixVbCvrG9gs19DsAnU1YiPoOOY9SThkpHOe4HWpNaieMKslrry+WSw7MjKxo2E8/PDrHUhS12cxQ45NcdrB8RmUhaxrgvk9JpvxvCfbs094Dbz3uprozqLFjwGSCa0RacBi73nv0CbHGn6eEcwGLP+bn897ybpI2YvaLxiDXI1DFzzscwHUuJe6vt5T4Khp69UdDhywzzarJr6Gx+qD1sXQl6WzKUQ4xrzSQwCLG9+8x5Z/4FjptNOqVG2/zhwJNtH5XAFOTdFAq2l7aPU53F6Iv09SE4/FGoEEYEgGaWpsmkKFKgtTq/hn14iAW/ZEyuRSOLGpTvw+RjY/fB5JaHTzg+ZMhb9bJgKfNYKTdQLqBFVpQad1yPZanNvpVMD5j88+9yJ9uZzUeXy9egE+11NMdQNhAkGqkG1e4tqmAHKX8ylrLzV/zW7bgJW2LJ/yqyu46eBBnH7hBZEYBoZHBVTQKpHvIXCQRErtQ82qjvOVB79473xNbcdhwJlsfwnQuHnZQBXrAnkViQfNOc9zv+ftrcUcd7bTmnNFBrXMUn4Z098In16poN/zTWp3bz3Y4TMt+GxLHaDslZaIAgLiBCw5EYRdTesjSZRMwIhAsM21vAey7WoY+Mf9rwdJNG6U+2njwMCPrWdQpFIHbmmsu/NgL0SCPGc5xc81y3bfO/MdLltqeJqyLHfztlfTGZjs7QENbPM5jfwAn1drChSXQeoybni6HtDgfWC+FY/fmnTWb9Cc7Midqo2cqsc/H7yWvbnJhYv7HCgDSH2eCdVAHRz/fL+dEIDbHt6w6+32QHyudI+3kSiNGP3yX1vAiFuO1bPbum43aDHcOHnZd9pChnr/LLBHz6qNMa9AsXXLgUTOWUbj0KuN3KByGOp3fdyNoIT/R/v4rX/zh+PtHV9RVPwDA+CVH//jvQI3pU2+rj9uofDNYxU6rjnvnJysCHTsFx+WLakiJb7OJ5FXQ1JCF/Qm314XMGcBOuZ/Kw/RbaikBys808mzEBRk58AOTnT84sLBBZobJ1kQuY3DDdPOti68Zw7oPNWksgmlV1B7eSibpUEWIhZa5KWxsYjPl7ANnwVgGSIvVoAsdswywAoQbtqMRWKTkpvIJa0wloPJ8Ymam2ehijHnneiLJ89iclNrb5PgN8gqZNxGiIwxa+ybJNMKfysEFEJGuw83wSk4zTGIxCJRsWALjkkKTS5KBi4LG8tZsAAsMgm5CJMJwbBoAhYs5jaLBTGAKH02sKKlZj03tVQwsNgjM/DBt/9zvRdZPZLEOU9OjisWcNykkjUqz0wH+tAmgdeJ10dsuxgLOdvM0mJgbo5N6TJmZmeUUcFrziYjLRROnjiOzbW1nqIiRL/dVhO3HT0in+NyxWS2vOdqijfqCjfleyTTGaSTtNyxuw7anQAAIABJREFUsWAFUlCs/Y31tR4oxWKYodk5NlNCQawur+jaMQCzIWlxs6eoIJGTbBWpPjpdMbM21texa+dONGoVLF6fU2NisD+HerUsJj19cgVQsJBmcyZkGx6CFNwsqogPWFFPIMpYKzbQ5S0bscAzsRBcAaFF1CmTWNnQ3orNKG7O6JFNkCefX8POHZPYt3+fPMM5frgJVP6IckTsOSZQkcrkMD0zi+GRMSSTaTX0yfJNJTPGXKmWUCtv4vL5s1iZv8gkciQiMcTZMOIGgE03Bd0xoM6aGPYcdDQmFpaWkMoM4fZ7H0AkndbGo1YoKrA2OziANi0x2FwLBnsh5cwAYV4AQ7DZoCXARLYbD4g+8Qz4pEQ2m4yoccF8lKtXL2N+fg7r7v4+8+0TOHjoMN7+jn+OXbMzCgxmMTrAZiaVFJubekao7KjWSrou9LGlwmJ1dcUYiSBQk8dXv/o1/Mav/wZuuukgVhav4LOf/CiOf+urujZqUtTbiCbS2CisaxwxUI8s6WgwiPz6Ovbu3q2Q6J2jAxgfH0YinkOnE0OlUUelWZT9FL+vthqok/FcqmLnxCQOHz2C/rFJdALWjFEouoJUm7LDiAmkSIupzgKUap/3/o+/xML8FRzYO43d0+NAKob0xCyyYwfRDGaU6dBq1VDaqKEe6CoMt7iex32vuUuNo6X8ugCi+evXcWD/bjx38hT2ze7GYC4noCLQbYOz+bOnTmN1aRU37z0g9mIwQXVMGi+ev4K/eNcf4/ypE+jQa73dVDOLQBbHaLNTUaQbAcB0KIy7bjuIfdNDmB7uw9jgMPozWaSiccuwITuXgESMoewGVAi3DQal+qE3cCiRkvqJc7sx9tiELWNpeQXfeu4UPvh3j+CFcxfQQBC5viHk+gZlmRKNhZHrT6uZ+gs/+3Nq0MbSKTVu5Z9MtpLzO+Y4EJPY2aCs55npUMOFC+dx6OB+salV6Dvmm0fqPdvISAMBKQIYpOutAr31jBlFhfD+D3wYH/3oR7CxuopSaUMgV6POhqeFtLc7to6GugmEAlTVNZFOdHD/HUdx9KbDyKUTaNaaWFhdQalex2q+iFAohkP796PTrKBVKiAVCaBTr2Df7hncdPgQBofHcXFhFU98+zl87NHPoNJoYWZmlpoIxCMtvPH1r8XMzD68cP4afuf3fh/BVBS33n4LfuBt34+pyR3o6x8EffNHx6ZQKBbw9a8/gVqjgMnJMdx8+DDW1zYwNjyJiYldsuRBJKgG9MZaHk9/+2mcO/0M+jJBzOwcwTe+/Bj6B/vwlh/4fnQDSaytd1Eqcs2Ioh1qIhwFXnj+25i/8ARmpxJ47UNvRiM0gfl1BnYHMDAwrOe4XFhHfmUOL509jlSyhnvvO4qp6VuxtE6gIi5Fx3BfDuWNdbzvv/8pnvjaZ3XMjTobxOIzC6j44QfuxthADrlkQlZRuVwfkqmsAo3XSxs48+I5rK2syx6LdiEMr5zaNYGpHTswODyEapF2TA2BdVrvmUUUiyCWyiCRygoQ5rhu1mtqcq/kN/CpL30VH/3ko2gFQxgbH0elnEe1sII3PXSvnpPc+B6M7D6GCrKyx4oRqBgfod00NvJ5rfnmfe2AClkstDV/+iYixzGbOgL5U5x7Dajg+uGBCv7b0tIqouE4EqyvCN/U61icv4rj33kKl198AQPJNrL9UWwWN1Gp8HPIvicZoIVUJKLrQitC1nupRBL92T7ZKA4MJXScrA+ZX8XPKjPoOplALMm1hM0y5otR1dRWyHi1TkZyHJFEDNHsAPYfuQ8nTy/iye+cwE23HMCu6XHZrnDHqyZTgHUOVR5FNYeW8iu9MF/f8O2RS5wlKdczU7VuARVUudA+YyCTQ4J1KzfltFGlSrnTlqKCjYWhgUGpx166cEE1BTNLWHdl+/u0rqeySa3Tw8ODiMdSCAejsks6d/asairaP0mdS9Z71GpzU34Yq5oNK9tYm02Gmr/NDtoNa9J6Rqs1pBmOvqBaJZNJyQqIF0Z1KZUL2xiq1hBio2ELqIjEwkgR4EhaTgiBCjZr5CfvLJQ0EVEdFrW9CIEKXm826pW1EQljfWXF1NgRa0hyziWhhPcxmqQXfgBrpxcFQChfhBZ+Dgwy65OWQAFec9aQtChTE8XZ6ugQvF+5s0ixRpTVe/zSs+CY2Po5m6NaR6y55/MsVHVJFeDzJcw731tOad51eyWvtFAAsdQNVEjQ7sQ1Rl1mg4EPEa0jRoqy4+k1R90xWoPJ7Fvkmb1ta8r7zLXQ237I3sc1FDlW5efuGJ36Hcdw9ddAqhxZA5n9Fesv77/vG8XWBPO+8sZaNZKV2QHLhqlpRCTZenL/4/I4fEiuwohd81phqM4GxWcwKE/QZex54IOnac0/A+FMNePWUafS3h506vMXeT+91QsJb0YqMzUF7zr/cM459dxzAq6pbDVgJiQLyPMXL2GjWGacLtrcUzEAnAxw/W05XFSPcv8TjhL0JRBAqx/a7VmzyWoBMtGDAiqoGiLAoXne2XlxTLDGNwDOVOd8zixvwIVru6a2eeW3BXjJgo7H4kJl+T33N3wPPYMueFt2Ms62yWoUyzxQiLcIFv5Z38pr8Y12EaLomFAuKwzZ79u1RyWxsWUWU9Zk9BbEZj+juUagFPeXtldVI11ZBMasV58g5HJDuI9tGkhAchhV/QTUbW/ogo8Jpsgax1j63qpGz523ZvuuMOsQ1XPeaoxqEgdM2n7a5kG/5/aAmU0Ptse3vaF9z7HJ6629ooiOti9Xdg3Pj/ttB3JwTKqG83t415PgGN+yLdpizSs3JkDlQk37Fq9sIwBGK1eq0sTidj0GfW7PMrQtUF/1H/s6XmnjGsSy0W5ZHpXImpzn23URyvbOzuLC+QuoVJmV1IcmFYlU6ytbwlTkbMAbuGUEVs5XfJ6M0GozEa+HGuJdZ+Wt7rCzoet60Mgs2DzRlWOGwIUHqPza4TNmVBs7oMI3o9UjcqCmAcyOme7zJzQ2DXT0IJ1veMcSMWUTmvKHVt4WqN5zHnF2QQapOMcQZ93HuYL3hjaGauYrZ9C5GDhFjnpjYA1uRN6tNr+RgNnTMEDRCEvai/j9g7NpNxCGz+82Mq/r3/g2Nq+fAdi2JpgVlTlqmO3YVras+gLOJoxjU8oHB0r7n3tw3t9D2Yg5sJzkR9/T6wHXTrkm5ZEDUr2lnEi0qksMePRrim/4+3nhxBdeHqjYUpS4cSUloiqTbS38G/uyRhS2Bc7Oged/4+/cAFa8TFvXwwMvB2pYT9ByN/0589rx2mqed2pJAy/MBLj31cMdzEJtC4j47iO68Qi28BSzEJNC5hVFxcvcuVd+9I/6ChxK0V7Bnt/tAIFJ6VzItJM1iG3kJhwxtl2z3+MBPYaBC8Ti74vRT4mo/P5M9usRRz+h3ZCQ4f7dgyfSWLggmh5zy3nSclHVxsGBAP5G3PBo3zApuMlJHuAe6QzIhsOzM3QsASsmuekTaCMk1KTqLBLUrFWxxEYqiwwr6sVYc0FtXKR1jVyxosmetjMs+BREbFZHnnUnnJjsEwEktsn1sjF/XpwItdj7TYkL/rZr5RQwzk/Upjqi+5QP0x7Cgs2UNaFGh6HftvGyAsI2PSYtFUPGXVmCEWT3eCaUB6b0GtkO2aLrkXF6etJqiH7oBJMITpA5wT/NTgsPOaCCTQCxZ1wjRDZiDK6iUqJeN6mkCxqK0T+VxV2rqaZ1Km6MetktJZLYyK8in1/X+c3OzoqBxN9j9sPxZ57GxsqKMhR2ze4T64mL/E03H8TA8CA2i9xwmQSXRS/vCYGDjfyGvM19wcn7z+LYe3fz8/gZLDzIuOQVJzuar5efbzyBTC6LapNNxZY84dlgoV0Nfae5MSXrhxYas9PTCn5eW15CrZRHYXMdpWIe6DYlv42GyXwLIRqKyj6KhRA3BRxVZGwoWI/xVgpkMcaKAAt+z/ESNl96yUodMy0gSayNAd5v3meOa55vKpV2Nl70dDUpMm0lWOTyuG1sMpDbNul8tMnunJjagbFx5kL0oUPFRyyhDX2pWJY9SoQNtkAHF888i+WFeXSqDaQTFqKdSDFImyxes+DhpoXHw+NnMPmly1cwOjWLO+9/PcKZFOrVGhqlEkhnywz2I0AfbD2TITV/mf9B71gxpGjxtLqsIoAMZWZHZLP96HQJvDZQLW8KeFpZuo6lRb6uJHsPsuGfeup53HLL7XjTm9+KfQf2i0lEqfng0IiUA9p4hnmPyDpjgDmbWpsoFTextrYqgGd9dR3X567j6aefxa/9yq9ix9Q4Ntbm8ZXPfwannv4WWlUG/zIsvY1InIGtZmmW5HgKhZBJJLC+uoqZnTtx2/ROTE8MYWxsBCODk4jF+lHmWGoVzYKqXMR6KY/SRh7dcg3jQyPYd/NBZEfGEYxSLcQ8jhbaLKKlwKIag+qhlAq3wmZBzOS/+eD7Mb9wFQf2T2PX5CCi2QxmjrwKozNHEYj2C+QDmrh6eRHNYBeX565h8eocHrj7PkTiYcyvrmBm9x5ceOklHDq4F889/zymxsawY2KSw1EhySzHnztzVv78tx08hFQyim4kgOViGX/1nvfjfX/5l8gvzQMM33bgKzt7YjmhpqZbqAUMpzJ4zW0HcOuhXRjLpdCXzmIgm0WaAe20IuQ8wyZfmkG2ITUG2ehX8yROj/8kIqmsWV+5OZzzAechAlEvXrqGT3zmMXz2S19CodpAKB7DyMikMa4DXWRyaaQSCfzg9/0A3vTGN2J4dAR9Q/1qFIlc6oJTNX87RRO/L1aqWF1bx+nTL+CO249iZGjIr7auTeJnfwO6e2vB31v17F/4Wyurebz7z9+LT3/6UeXDlEt5BTW2G2y0UE3BddPYtbFwCqFOANFAHXt3DOLH3/JWHN6zB7GwKdvKDActVbHOjB5leACxIBBn4Hu1jE6zhh0T49h3+ACGxyZxZWkDn338m/jM419BNxDG7ceO4cDsLjz5jS/iwL4ZHD16DKfOXMV//qM/QWIgg3seuAc///M/J2XPS5euIJvJIds3pHO5fv0K2p0CUqmE7kEoGMX4+DQmx3dheGQcpSrVLvOYm18UUz+TiODK+VN47X13Y+n6Oh77wqdx0617ce9996JcBVZW2iiWwghwjoiE8fwz38Da3NPoS1bw0JvfitTQQcytdrBZaWN0ZFKB6pVCHrFgA89+5+soFy/ie956PyZ2HMZaIYpiiU2TrsCHwuoK3v2H78SJ576BerOIRoPWgWxCBNGXieDt996J0b4ssqmEFBM8TwIVzAZaXF/CtbnrqFcbqJVp61fA2NiQFH+ze2YwPDKCRoUbyQBa9SbWVteUJ8K1JZXNIZ7KIJ3hhi6grBfOXcxW+dtPfxYfe/QxJNIZDI4MoVbaRLuaxxtfdw/2zwwgPbQLw7N3ohrqR7VFj/UIdk2NIRiIKMOGa6FnHMoyhU+cC4ulksdvvAqFglMPmsKS68fi4iKmpqaUFUVbKwIVwWBM6q0UQQI2OktlAcKf/ugH0SnNI5vjWtVCs94Gyb50lGy0qgi1gWQ8rrWTOT0kDuQyWYEXfYMM9TTiCDe+BJB5DTjHB2JRgROsaep8z1YHm4Wi8irIKKZdYHpoDEfufAPWC1H86V/9NZrtKg4dmlW+BkO7RUWh3UmNdljmQ05FBWsrhcW6r15zjtkWDpwQO9j94Zyzli9i4fo8BrN9SNK6RXfRLDk6VA7l81q7+rI5dJttXLp40TGXywIH0szRoqogFtY6x+cik+4TACSg4swZrXXZTEb1JRtHQdo29sKXrbZlI9QIB8auVBNJYdq2nm8xD22+WVldVI1CaxqGeXKWkULDWV75hobVh5ZhdfXKNSkB46kYEumULKBICvCKCs/890xLrUOsZ7pdqUMIVLBhY6qKCNaWV3QNuFZZllUEiSSfpZRs9qSoOLvs6ms28ywMlGunLJ+8cauzJGFjVMCE2JiWp8f3tVBgjhtrTvlmvYGDZl3lWbA9pq5rWPoG+fYa3ROkVG+7poU171kv0WLMFOZs+DO02jf0TUkHkVBYA1FVYcoHFzrq3s8D2L4Z4ptMBpRY28bv69RwdpkQXuWhY3bMbp4XP8efF2sa2b05n3PWjdzXUMnMxrk1lE2F7clkyuRzIaVqNKrJy8a3NdqlQo5ZCO/W+RjxzM81RpoyYE0g23Z2q5tfNGbdnqXniS7feCOB8XWmZGjbcxsOK3vOshLMNcA3wXvsYBJ/XE6D7El4v0WGi+CF508qMJjqZpbTzLjJ9g3g8rU5rBdKoKN/hCoD5r64ppSOi3u6SlUqqHqrrr0V53Eqkck+p4Utj4PEJJKT3/CGhwQYt5sNzXkEg8yexbIL/F7JNzP5/HI/wvNiQ5X7DxFRnL8/92dSQLt74puyVJhWywRAt/IPqGLmlyeucc/igRFvtWTEMrN24b6hVuU+hzZgzEas6tnhh/E6cjxzbq7T6lXMcKtg+Gxx7+fvn9XP1pDlvfCZOhpbzo+fx6XmJi3aSFpz2ZhSdDnvew/yaX/Ca0DgQ1aYZjct4qQjOorE55jiPCoBEgwQ3vZ+nAvsGH1mpE32HkDwDXMBKQ74EUAoxZk1wn2OgBwHqORX0LbNN9bA9vt5Z8HnwJSe+ss1xZXD6fIW+D7cY9DBgJ9L4JfHbnka5nZhBEkDjg3wYQA3czXNronzmLHnzWrOq6R8I5d1HmuXerWEaDiEPTMzOHnylMhsqdyAMipopcjnjft6wXtSmjSRpIrYXWeOd696EcDqVE1SFfH5FjhlgBSPxf8+rw37O9xz81yk4lQQtl1/AV8KSfeAh61Vvj8j0NWR8DQnOdCVY8DPa3yFJ7gqj5XPQogkxCKyuaz6C9xnW1Pb8hs8eL3VDTeogs+Fskw4LzpQRufgHEmoOlIjXcAb50WfH+JUGk7Zw+dYc4ScPwwIY/2STJp601QqHjh0RAOPAAo2cY1sXmdHMvEZNyLEunwam0/svFQf9LJoDEji53JNEiDiniPrg2h1M8KjIzXoOrvn0/dK+I+61g6E0FFtW7N0PV3j0KsoejWUm5P4+pcDKvhahU17AMeBJVpfOOZfDm3w2R8OLDOCsvXAbthZ+bXGZZD0Crx/4JvtH+WBP5EyncrDg+V+nvVrm2qobfs5G2B2LP7e+2vtLp1vl/aWw+3KCr+e6XdfASr+v27bK//+j+0K7I+bLNDQYfedPOOcKsAzrqVisEBgFfK0felNXE4q6xQGHgHn+0niqEXW0GM/jxpSbIiq/3ST/dlGjx3FnsRXM7ZNbGIAOc9Dsru4MKs4ZUHsFn97sK0Y8IvV9nNTKzdsEjM1xy0l21QSsELaXg/Zb1C+zkBnFl6SylG+6xQeXJx0vG5R8QF6YmC45pS3ktLCqIKc52iMJ03W2idysWMD0Rbn7ZL6LRDB5Tg4f1lePxbfPM8bA7e2RqGKFrfAKdND9zWsDbeh/SxojJnFL15PnospSWyjw4apGCKOweMDp7wNk3gFAq1oxVG3sCgGadN/GWRHMky7Ibsl/uxVD79Z708wwYLAjdnt/RvJBJJE0PkI8lrwGPgafqbYdg6oMM/ytMKFObzyedvkEqxg4//6/Dyee/ZZZSQQqJie3YdAKCKG0+69MxgdH0e13lLoNY+BRT8bNNyYc4zXGbrZaKJULqLmpLgszCm15Qa6VCyYDQQVHmxss7nHph5lo33mRa5YMz5TjTZy6azYzHw/2mIV8gVM79olayFZZFy/hnppDZsbqwrBDQc7SMVpuwUwcD0cZsh0Qs1vNrqYhcJNtzYx0jAYUCGWk1QJVhCSFqPrL39Zx+Jggd/LB+no2lGBwiJkdna3WKlkIrIRa8+eqRy4mWVxQ3af5I5sbqgoA7L9/ZiZ2YP+/kF2wNGml2mYwddlxNlkYAEUAmKBGp765tcRandR2SyocZOWlUMCIfnIOwm/886lwuX8hQuY3XczXvO6NwuooHVRq1xDq95AIpdBPJsCRSTMZ+D1poWVl6nzOS3XiihXqgIreN2YS0L/cRZkIQaRd7tYoC3J9TlZTSSiEXlgP/7413Ho0M14w8Nvwp79+1BtkJ3LjQ2fiw4SZOTHImIGco5gY4vjYnMzr8yRoaFh+d5+82vfxPFnj+O3f/N3cOjQPqyuXMOnPvIBnPjWE2jX+Tqg3uwgnEhhdX1VzRjOO7FwGNlUEquLS9gxOYnbdk5genIIYyMjGB3egVRqBAEGbnbpFV/BanEdC6urWFtcRKTRxvTUFKb37Ub/+BRCcVpJtbWpbTDIMUTGXRSxVBLBKNlRHeQ3NhVe/IEPfQDLG4vYuXMMM5NDSA32Y8+tr8HY7O0IRgfEoA4EWrhyZRGNIHB17irmL1/FXXfcqTGzvLmBQ4dvxvHjx3Hs2FE8+eST2DM7g5mpHQIqWFa3Q0E8f/ZFVApVHDt8k8nRI12cunAF//Wdf4jHHv0U2tWSQrSDzjdeQAVBt0DdWI+tAHYODeK1x27GrQdnMT6SQyaWRDKWBAFObpxow9RudZEUyBeVbRL9ormpIEgZT6YQy/ZpbvBya84HfJ7JIF9YWcfnvvQVfPgTn8T86prsdAaGRgTI1VsNxNNspOZw5OAh/NIv/ZJyUciEN5TCW3/Y+kaGpepSBFCq1pQbcub0aRwTUDF4g6z3H6onfEn73f/O93zpyiL+6E/+DF//+tc1h5SLVFRUxNLk8y5gkRARrdlCCUQ6QDxQx9sefi1+8J67MTk0hHQsoeejG4mi2g6g0m4j3y6jUiogRIUcG+qFPJq1MoYG+rBr/z5MzezBcr6CUy9expW5JTRb1kRJJWLgMhUJtZFMZHHq7DX8lz95FyLpON70vW/Cv/yXvyC7uKeefgavuvPV6HTDePTTj+Lw4QOIhGoolQpaGxhgPjAwipcuzWFjvYDRsWE1d9nAzaSTiIU6eOG5pzE1PobB/t1S2T357S/j/tfejQM3HcHcQh6bRW7YYwgijGe/8w3U82cRaM7hwTe+EaPTt+P6egBrhRbGx3aiVKqhmM+DZPD82jzOn/0aHnroKEbGD2K9EEOpTMC7i2wygcUrl/HH/+0/46XLJ2X9ROVBq0XyApBJhPAD99+OIa4H8agsybLZPgHNzEu4NHfZGgadgMBIzj25XBoHDx/A3r0zUtB94XNfRSyWxBsefJ2yeUqlTQwODaBvcACJdBbJFAOpI6iWSihtbuLi9Xm89xOP4vGvfQt9A4NSlRU3VhDp1vHGB+/CTbsHkeifwsDsMVQjQ6i1QsoH2jE5JjB8YXFR/uqe2ea93evNFlZWVzE4OOjsgxoCkdh4TGep6rDBvbS0pDWNQAXXQ1qIEdSjkiQVTyl/KhqMCGz+0mOfxvPfehyxaBXEPmlJxtBwPiiBUBsJNrBVF4W17mdTaVki9fflMDBMWw8+ZqZcEMjYIHM0ii4brwQuai01UMhgLpYMbGDTvR0EhnfO4NDR16FYT+OP3v1XuDZ/CQODaa19nGv37d2LyZERVKplFDcLsphaXV9THaWmnNug+xqN4v8tcMLyAwRchMNYWy9gcXEB/Zkc0vG4sTEDDG0mWEGgYkPHTxAm2IE88dmcqXNtCBCoyGh+ZFeI6yPrEAJekVBcKoQL584hEY1J1SmrCDZko9b4ExtepPaALDK5nteqZivzvwYqulhZXVI9xM+LMx/D5V34Jpy/Br7B7YEKNrKT6bjs714OqPCKSV9rUy3HnxF08YoKNmQJTqwuLal5EmcttM36iZlg7PCySZA/u6y62ljHDqiQbzkttsh25PgwxbMdc0iNFNbBvA6s+1gneLa95UVs4cOsf8zSiQ0+12CUKs/ZPblwVplPsAHiwknVuPfMeNoiOUtd4uRiuNfrjrVudTjXHdYkJD2wacXx45u7MpNzwAKPTTY6MiezUFp5/DswReehQNyGxosFHdv+SlZXavaQYduWQpi/b9fb1B1qBKo5ajUCf6YGoXvKuf+Q0trZ2fB6qakuSx6zHfF2FHy9QmzDjj2rRmhUc4MC3h05yrz3LeuFwKkHWfzPZYHo9oC+881z8Gxea8SbWoAnYI1Oa1SqsSwVjAsTlsqAbH3+jE1fgvNmXav9BmtqnmM4gpPPnUCL5CmSJZiH12xjaGQcZ85fQLlB+7YIGiS9aH/nHAZkv0VVR0D7HjpWKtOhTvcBU2rx2Ana0uefv/f61z+IOPdErbrqW/6M15ivIbiuBm8goOfRCG0R1BwAxFKDjU4SURR0vq1Zz7mA14HgDet3qrhIWuD11DjyGRV6MCxEWPtrEkKkGrW5jvWtiFjKyYjrefVB1J4Bzz1zOpM2C7OgZWWQ9OezApoNZ0mja2OECJH3+Fw5twJjJJsVtJroCttmCDvVE6xfSfJjLmFT5ZXPtvDscb7GW7l5xRP3sMl4whrn3OvW6qa2dRk1FsjbAbNgVDOSfCiAjeRB6xfQOYAZGB702w64GjhkFlUWXG3B3VICsXkp8DMo4owpNWxvRiCfJyFlYMAyNgSExxJGcGNjVsoEs23m+LZ5ypQeHOfct0sJ4+z3LAfASID22bxfUYGM/NJnuXtnahcjY9q86BvszF0IoFWrYd/ePXjx7BmpRFOZfjSZreNiCbSuODsy2XA7O0QeD3s4IhtyHnZ9Fh6QrHdpB9e1PpPas67D3AOTXEi8qbWMnGTghQFqdj3MmlvPN0Etdw/YdxKR1eV5iigkezIjQ8rhwKlr1O9w44/nzn6PAJkUiVjQ3Mi5yq9TBlZY5e3BVQ++8px7vS0H2PleGV/H8aPcULWcrOfSA0vceZEwyHsrZRStvZ0dtgXU95z2TCXiWcKebOwa4LwW3Nc0qETv2HPP++BBZd9I94o6zZMO6DF7MHPkoDqEJEJ+KeNEJgxG1OU18QRnmzasj6benVNoKJSbY1gqDvsM9QzcNVePZ1u2g+pNZxH494GKfA/c8KofdxPP0zbwAAAgAElEQVR65GcTTTgSMi+Pa/wZIOHD0E2B4w71hnvp91MekLqRHmZgS28B3IZSGDhhWS1eOWm28G7scu2QesQsybSGur91DbbfRwdS/T2gwh2cjRvryfjn2wjRzqL/FaDC38ZX/v6ncgWYUeFlhybjYiFsK5CX1qn4c+oK72lnRZ/JN33hyN9Rwey82noTu/dF9Q+ak3Ruf+BtvTX03y96nrFHdjQ3zWIpiEFQN7mnY1uoueVkbGoIOxa+WRVxore8C19UePUDf48PuBqOzYYKFiHgPdTVrJnMg9HZY3l5pysQjE1vTBJeJ4+gakF0C6gmqG0+jX6DpqLKMYlkX0XggtZLtG7q+Vf6JrH9zCZy709rigPehy0GkTG0bBGnZZZ5THPG7nRNbt+bKN3ixmOQpyLZQCzSnVcsiw4vW/SsPMvF6CIWjsl71LOSeNGabITZnRAwoRBt+lq3yTqvW4HZbmHfq15jRWciIbCCzSx+qXhgc4F+2JJeW3HNMcFwZZ4nF06x7WJxMR54PrlMRkAFrZ8UZFcqyeN89+7dul4nnnkG68tLNwAVhGAmdoxrYe0bHJFHPz+TdgO0FKBHNxtCwTAVEuYjTDYPP5vnzIWfzQ42/1jIsKCgTQO9NGmbs7C4oMJJDZNQWD6pyUgCfdk+NJpVFEqbVjxGosqooGKFYdGbqwvYWL6EQn4VVDxQzUBWPe1AWKxy88Ygv3iCn5U1xYKKYYJ7LIQ9UMFTs5+roI2F0Og0wcBHC+e1ok2LncIM21heXgKtkqTwmJ3Fvn37dDe5yTeGmzVe5FfOzSltI9psAPFq0kqCJJuo7F4mJnagzWyReBL5zTKCsqpibG9XIb2hblUhqieffhatKlmzbdmCMHxXm2r5b1pTgX/I8H3xxXM4eMsx3PX6tyCaoTd/A10Gc9ZbCCdjSOYy8m1nQUvrEfqk816xKGeDBWFjkxeLFYUN02N4564ZKSOqTSo2XsJLL56TmmCwr08+4tVyFZ/59GPYf+Ag3vimt2D3vr1i5jK8lT7nskxyrBveI957Hjj9xTnvsFlKv/tcOqcA67/75KfwW//+N3Hw4D4sL102oOLJr8nrX7LpThCBcFSBrWSvchNL27P+bAbXr85hYnQEt+6axPTUsICKsaGdyGYnxOajkVKtWsaVhau4cPUygq0OBmIJTI6NYXTHJIYmphBJEOBpyhqLDQ02xdiUi6fSCHAOqDNQfB2ra2v4mw+9H41AHeOTw9gxnEN2ZAj7jt6NiRkHVKS3gAqGX1+Zv4brl6/g9ptvwVo+j3Y4gNtvuw1f+fJXcfe9d+HUqZPYOTmO3Tt3ya6LYAZDuJ8/cxalQhm3HDiANMGxEPDo41/B7/7H38P5U88j0GZgckMKDGOtOjltiH68XYQ7Idy2dw8evvcY9u4YVjMxGUsox0bPjAtY4waFCguBtMzaEbsJ2tR3qbJgPoX3uHa2CN5eY2OzhBOnTuODH/s4vv38KXS4kYgkMTY2jk6IYFzAfPSzOfxfv/bvcOgQrZAG9Wx611Tj8DjRkypVoFSrq/FrQMXtGHZABWX3Zoz4cl8q7be90fbfCeDr33oef/iuv8DpF06iXCwIqKgTZFeANp/3DtrBprzdQwgh0Q1iZrwfP/djP4jDY0MYSJmNFefEQDSBGiKod9uotkoCKjY31rCxsoRmpYJwoIuBgX6MzuzB5PReNDpBrG9WsLqWVwOQY1chzxHO4w2US3VcuLKK3/vjd2G9WsA7fuyH8NM/89MYGRrBY1/4Iu581avx5a98Qxk9r7rzdjQqG3jqqW/hxfPn9Jzu3rNfYddUb01N7lSj4fLVi3jhhRPKfAl064hHw7j16L3Y3CyivFnEhQuXccedd6ETjGNts6RzZnbKd775BOLdJZTyZ3HXfXdjz833YzEfwXK+ganJ3SgVa9hc30AyFkKtso4zp76IB+8/jIHRfVjLM3Q2ijpVcqkkzp56Hn/83/4L1tavot4ooFZjaCDvfQuxaBfff98dGBlkkz4mdRTt8GiRML+whEJhQ4B2inZ5zIco0Iu3hfHxIc0To2NjUlSUK3VlvHDdu3T5IhLJMEbGR5BK9yGWSKuJUa9UZDl38sJFvOcTn8Hxky8i3Z/D+Mgo1pauoy8ZwpsefDVu3jOMcGYMuZ1H0YiPotKOaN6dGB+VHR+BCq+o4Jhlw4oNPDboqOgYHx/X2irV4uam1gSCzHym+XMCFXw2+vv7BBzPX5/XverL9gsIaTDbo28ItWoD1y5exKc//kHk1y6gPw3Z3DWqDTQ63AxD6gcFLXPzy4ZyNI6h/n70D/YjHu8gGo8ik85pvuSax8ws/umEQwqOJ0DJRl+pVNG9pwIxGOqiEw5g781HsfPAq7FaCOPdf/k/cfbCGaQyZm9ESwuuSbt37cD+fXuVHUGwfXVtVU0Gy2vwbGdrZAUiZPBac9nXeaawCCvgfGV5CX2pDDK0rFSgMm1h2grU3tjY0DpLC0HOj1cvX9E9aLRqmizS2bQ1XoO0dYrq+zjzSYIxWVVevviSrPEIIvE6SSkZswaXhQzb36l0Ug3kStka9P9/gAqC5+Gw1cWe3KImBevkGxQVV9WY3g5UEK7dbv3kWa4CeUgQkq1fUIoKqWZTKdVNrEeXrl93CgOSMrg3CSjPh02/gIKKQ8ifW1YjUCxYNu22gc48d1o/8bVsHKmJ5xq1ykWQwoE1tgFa1sS33zPLC7PDYc328Pc8gHtfdye+9vi38flHnrB8OdXtVodrD8JGj0g4lmP3M7/049g5M4mPfeBRHP/OSWdt4tTMLs/BM6x9mKr3Ref7eY9+qcu31fA9gEwsVLOb8sp2NfQCplSwxojrsTiGsTWWDXjwexjmubDO9aCfD2yWfQ0bzq7RZkQq439a45T1fNwxnM1GxIflcgyb/ZiFKasJJ7sbt3/ZFgq7/XpLUausCatqNV7cufh9j2cpy/plm3qdjX9/Pa27Z+cuJrH72zfTzBKKz62xdHUesjxq0yRSbPGzp15gMaqakHUT9z59g0PIjg3hP/zhb6BYqODuV/2whf6SDOYsflSNs67geh0icY48Fmu2cpzpe90DsqXreNMbH1Y9RqJTm5lyAovaOHLrAbzlex/AtSsL+J/v+YTt0QTQmEWOATSOXEZQX2oYA2IEqhEgcdkTnMtJ7lIOg1Gdtb/3jHF/zz2444l2Iq5ZWW6EwkhYCiQ/Jvm+/Fxj89szwPGnpqy89K1foOeLxBrlMriw5SAB1KTIWrIqcu4NIhJyz6/3pqqe1kIkFG4HBw10FECgMW+1lW9uc48upZeyL/14p9I6jompUfzsz78D1Uod7/y9vzQHAgWtG4NePQKp1L2Ns7M3ahroxTf+hV/8EezZuxMf/MBn8OQ3T/Qs4Gze9cod24dYFobt0e1YCTLUzYKLll9ScbiGqAiDlt3Bc/BMd4aWG7BIWyI7XtpHmdLA5jDvusD744k3/GyuGfYcmCJBgB5vke8xi4xqWZvBQAfVcgnZTAq7Z6Zx/MRxtLsBpLP9sn5inhtB6RDB9mbdsqBY13s7M0dONbWE5cvwfAkCGgDjCG5ygTB3Bq9G8L2Un/yp78UDD9yJj33sC3jkU19185g9zFJgqC9FBYudm2W4GLiq59qte5avY/0jfoloJxKuxYaaW4BzrHA9pO0s9Z/6qe/HAw8ewyc/8WV87KOf1/n4XowdTBc/9/M/hH/xL/4Z/vp9n8Jf/PlH8H/+8k9Infmev/okvvqVpzQPCOjic7ddJfZdJb5/prcr9ERrUhfc96LsRQI7HflUKha3VvB6bPWJbPLfskffUpT5tVv2ViLfGrDLMWQ9IQN0PPjE3/frkzlyWL3nFRncb/G42cMh0Mtx6RUbW/Owm4y3rUk8P698sfXKdk3Pb8uoOPIGq48EtPt79d3XTmuRWdvdMP/38igc6dm9zqz/tq7rdiRIY8bZKGqsOos9s851zhTufbZyc7YOyK9Hf+9W3wAuubHs7cFsprEhZYO8t3Drp9uVHu57my48IP+KouK7hsQr//lP4QocJENKjXiTpfmHSxOTZ/44FNtPWCziveTOJGK0zTEmTG9B4sPDAlMLhAv5dcWHR6FN6mmoo9BNIb62SGqj6IJ+xDZ0X1ywuThbQFrdrIrIlnWsMYENbE5K9WFeqGSwmiRzKxTPP/DGmiD6biF0YifRq5K+8vRuVzZC2+w6HDjRQ0IlJ2Rj1AKwbE7ZmrgpHfbFvP27lzhuQbF2zezkpKpwCKzfxFXKLKjMw1/WT062adWFvZ/5y3KidzLenleh+ZfymOQH6wKTWWAq06DbQTJhsmErDKz45OLHyd6kbFYYygfVeasTORazgawjMuyFFls+ApkevF2yfnJ2T41mXTZQXPwIXtz7lu8Rc58FmLwYu12FUNNOIp5OauHl+1sQkzG02PDiNaBqQTLQaEy2PjypXDYrhikZaLQCGBwcwOLSosAKMnmuXHwJhY11zMzuwfTMXgu8Qxeze2fFRqL1CxtFvPZsYpBVxs8gq4I0KPMMbomtsR0k0oaZ3qlUXJSKWpSzuT6US2TuUzYaU0N0fbNgxWQwKn9yLsFUP5Ctbxsi86JlA6q4voTyxjU0KiVboLoMHY6o0GeNHaP3diyBVCqD3MCw/mbDXDdXAZfmy2oLHRsKFj4ZikfF6uImS5tqt5nuhUIGglhbXcWlS5ewtLiocX/XXXcb+9LBT3xPNgG4WSdQIXZ2w8Ao3iX6xnMTMjQ8gj179iGYZDBzDOUqc0osEI9+p8waCKEh0CIVi+LiqVOIsgChxRQZQQGzElNoXKuFSrWGxZUVXL58GYduexVuv/dBxDNZC/NWoHcX4XhEigqqkji2aD1CJryYVWGqJ0IIxwPmYU2D+kAI+XwRi8srSGdzKNaL8uEma5YMEoIPnEvI/vrwB/4Ge/fswVu/53sxu2cPyvUGNgsF9A8MKYOBAJ+Bvaak4Jg7c+as5LrXrl3FwMCA7MleevE8PvfZx/Cbv/HvcfDgfsxdO4cvfPoTOP6tJ1DeWLOmCD1RAWxsbiKRjCufIhVnY64PVy5dwdjwEA7voKJiBOOjoxgenEAuO6YxzMyIlbUlfOfEs2i0m5gYGkWzWMJArg+Tu3ZganpGTWM+0wQjjj97AlMT4xgeHkZuoF9B5Azw21jbwOLKEt73N3+NaDqGsclhTAyl0Tc8hEO3343JPXcA0X6FHQe6TVy+tgACFdeuz2Hu8hU8ePe9Gu+b9QomxkZlQfTWt74ZL559ESNDw9gzPaM5ucsmHbp4/vQZlIsV3HHkZhXyi+sreNdfvgfvfe9fo7C2gkC7KUUFr4XmUOftTM8njt90NIFX33QT7jxyAImYsaposxbqBtW4Ixg6ONiHkdERZNX0pHKN831UwcEr6+u4dn0B67TNke9qGOFgWAqfocEBjR8y+ZhN8sjnPo9PPPZFVFptKX8IQtE2q4U2+rIZTIyM4qd+/Mfx4AMPom9oQA00X3Rqc+0oPlxP+FyValWsrKzj9Auncccdt2CE4IYKUgI52yg7NxQbDqjYJsX2YkKut5985At491+8B5cvXdIGkqqKZqMmOwmCPWJWBdvaGAfbQCoYxBvuPoq3v/kBDIQDyBGsTbBJmDY7rFgCHUraO2Xk19awOD+H1aVFNCplDOSyam5nxndiYHwK4VgStXpbDUmCfGpeBsJodxto1svs9WBxtYp3vvtP8dz5U/iBd/wAfvAd79Az85UnnpDiaXp6D3J9/ZoPuy3aqOUxMjaCW47cisHhESSTWRRLPJYi8qVNdDoNFMt5bOZXsbY6j/W1Rbz29Q9ifm4Zo/07EOjSPoX2MHEUqrRz45oaxZNf+zwG4mUUN87j1qNHcOj2B7BcimNhrYldO/ehUKxjcz0POu2UCst46eyX8dADtyA3tBer+TBKFao72+hPp/H8U0/iXX/wX1CsrKLerEh9R+o75zqq4h6+5wimRgaQSyTEpmd4O9eFq3ML6MtkpdCjKi9CO4VOE5FQAOlkDCPjw5ienkYqmRUwxrWgUizgwoWzqNWLCipP9fWZV3yTFkUtFAslfPvUi/jvH/47XL6+iExfBpNjE1i8NoexwSje+MCrcWT3KILpQaSnjqCdmECpGUUgHMb4+IiemeWlJZFDWAtwfabFHcdNrdGS8m5qaofqAq6T24EKs6IPYHlpWQBLf58HKua0lmQyOXSaXUTDMakCO822lIbPfOub+PLjHwcaG0gwJFxZWW3Ek7QcZLOaDGcSdAPumc4gx2DywZQpwmJkKJOBGECxUEahWEaTTT6C7G3mKTVRrzKgNoZcLgcE2kAiglvvuh99o4eQL8Tw39/7AZx44TgiCcHzzqe+ozWLzcSpqXGMjw6rdiLhgIpNhVczd8OFXlKVsgVUWA6YaqpgGGtrmwLQ7flKmoI3THC6zZ4P8sw66rQFWLH2mbtyDfEkWbW03WqLhEGfexJOGGzNNZ/ATCgQkbJo7soVrVmczz3Iz4wK34yQTR6BbzZCOy1UK6xnnOUIwUtaP2lz7htBRhRZXaOigjabUa2jDP2lQnC7c4FYz86H3hQVV1VrJNJm/RQjIYp7DNpwNUzZ2Tsu10jmfVaWUz6vmpoAFWtfjvnF69dVl5PtamoGoK8vKyCDSkA2WZZPzml95z0hZZzNA7PRMAWKAqjVkO0IrCYo6JtoVJ9aI9NYiarbCcSxScj3Y+3DZ69axVu+70Hc+7pXCah47BFrnvGCy3qChBISn9x+QnVsKIif+9c/IaDikx/6LJ5+8jnnI++U3+5C+ia8t7jV3sXl88nuRd7nVNcaIMJ6VSpjWV5Yw1p2sgTQpITgeXBPZ/W7rjftQJ0/v/If1Di3JqrsrpRVVkYmk9X+yhr4Ifzcv/4xjI4P4W//x9/h3JmL+hzeQ8uZoJWMHQ+vp/Yy2xs5LsDVFLlmReQZ1t6CSvsjR3JT5pkUq8Y+9VYYWkdd2K7fNFk9bnOUJ9PI1gZtrSnWfLTGnNlvuGwGFtOOpGY/Nwa2t7DlsQbY8GQjuVrB1YsX0azWBJbS4pMV/MDICILpOP7Tn/wOSsWqgApl4tBbXuPN6x6DaHVbAiVtD+iY0G5f1nF7AOZUPPyGN+D2YzfhJ3/6n2FxcQX/z3/+K80Tt/Fn//vbsLK8gf/4m+/SuuoJhVvXnCxqU4bzD58FZVmw2e8sWDyIRRCQigLr1NrY5T6H1nK6fq7Z6xvh6gf4RjDvr1On8LU+lF2KHUcYFLNfe/KurimVurI90bbVVCHcd3Iu4hfV3iJBSR1CBYXVPv4Z4Hsw94P3+NDh3fjlX/0pzF9bwr/71d832yin7ub5qz/gcio8K916C1vNWuVDhiOYnhnHr//Gz+p4/tPv/jnOnrnYs97pNdiN8+2Cfm1+tH2QgQS/+Ts/jzuO3YS/fu+n8OEPfsbujXsOeg1eb7fU7oig98v/9idw32tvxx/9wfvxhc8/6Yh7VLqZvY9vGPt7K0WSMgks64XrLs/NmP6QtS2zibjv9OokPmemZDJAi/fY+iNuP6/Q64gyrWQJxXuugGqeFyPASBAMoVmvYu/ePXjuxHOoNJrI9g2i1Q2iTkmYGwtUzZarNUQTBMENYCFZ0StifE6F+hoCWJqmYtAzYmPoLW+5D//2V34CX/j8t/C7/+EvNB7+9b/5UbztbQ/h4x97HL//+++zmdY3nW8AJl3fxQEiBoG4/oEbSwo4dg4DAqGcZR3f069HGndtZxUl1r3NHf/ml38cb3/7G/ChD34O//W/vteybLSX9akIXfyrf/Uj+NEffSve/z8fwbvf/UH8wR/+Gl7zmlvwp+/6EP76fY/grd9zH379//4ZfO5zX8dv/9af3VDRb/+PLfDRwLY3v+Ue/Pvf/D/w2GPfxG//1p9aG9utTz5X5QZgmfN62+XWOGKtAFinqpAlnSOweqDBnz+vm80bBvj48evzfXzfnH97oNSrE/hsKn92W5/LgwC+L7hdOeDP2YQhPivEek6yE2+3cfKLVJjb1+GHaHlq1+Tl3kfrgwLdjUTt3Uvs1X4v5dUM7k1VS1if0nqIlqerce0ARfUFnXrB9yK3wH97v+1Ajq1TW1aPJCzqlm0/Yf877l7q/XpqDXeM7n39urZ9N7gF9dgb+88TgPaKouIffLZe+Yd/pFeAigrPrO5ZXjhLJhYA/iHeAh38g04lgjHHfACTb677BX6rKLOL4ydFeeR7lYVCgazBbk16MjEoDQ1rkeDn+vej9JgFkEn1vITK2qhiQNFCyBXP2lSUK+Z56YAWFp9WwJn6Qc1WL913PoP8bC7m6vu6YDpuENhA8yBGT2LlJzh3/PYauz6cnORDqBwNW4g1aTs5GhlvxkJzceLf1ZMyJYdZHdn7eemnXR9uNggESFqn4CXPCJPRkGMmmFTUih++xiZLWtUIAXfHwAKIE7ldZ1sEFLKoiZJSSQsJ13XXPTJWiUkJLYeEG3ttlLrWPCQgwUKF1kEepBBw0Wnh4R/+59oEEQwpFoqgxzXfg+/Fxi/PiZtW/i3pNNmLytgIqGHCjRRZWvKbJVCRy+l9qgQq0imMjo3quJeXF3HuxbNYmp9Hu1HD7MwezMzspu+PmCG7D+zXJnojvy42xsDAkDZolNxSflkslcSn0sbP2WdZOLnPgLDlxyTxVlQbCMTGfFuMwFCYlmFVNdXZvLLF3QAhjvFmu45YOIh0IoZYMITzL5xEfumqGly86PTH5bPB+6cx9P+y953hUVXt2ncmmcxMZia9FxIggYTepPeugAh2iohiVwR7BbGgrxUVBaWKCIiiSO/Se+81vZGQnkySSWbmu+5n7R3Q43e+7+85l3lfLjDJzOyy9lrPeu5G6buR1hVWBAeHCLBiNvvJ80DQhUCNfj/1sc3jZWCwCku8ma8iGRPCFlQyUzbqs7OykJ6RisL86+jWrQsSExPFIobHotRJRrn/AuLw9Q3FKBuy0oqVZzipWTKsoXFivcFz5r2TzYEw4llwE+gywGjwoDw3FxU5OTDxGTR5i68t1QmUnNN6i82xDOZNOOuR0rYdEpq1gJ8tQGylFGBJqTWDzynrrsF15nxUVwvLlNdemh1sZhiZ56GafbynPBYCGsUlZfAYyfqm73y1BNy63V4CaBGEW7NsCZolNcWIO+9CXEJjAV4IzERGRSurgAZPUo8ocXj+tJ1iY4fKGo5Jo5c3rly+hB1btwvjPjGxKa5fz8SuLatxdM9OlBUWweRjFkseb5MXSssZhGiU0FWqKiJCQ5CemoaIsFAkxUQhLjIK0WER0uRkyCztb3ifUnMycejYUbFY8fU2Iic9CyHBoUhp1gzxjeNQU8tQZReiI2Nw5vQZuOuciImJRmR0BCx+NlTVOFDuqMCV1FT8tHyFgBuBIYEIDWXTPgCtO3RBVFJ7GOxhwqxy1tQgJ/86ar1cyMrJRk5aBgb06CnNt+KKUoSEBGHLlk24a+RdSL2ahrDQcCQ1TVQBg9wTwIOz586LdUmX224D2WKnz5zBezM/wN49u+X9hUlNqT/nQNoDiLLOC/XebmlEhlqtaJUQj9BAf2kSs41ABrZYcomdiPJlbxQbg1bNm8NuNoC25j7eFhSX1OJiWjqyi3Lh8TGK17/dP1CeW3+bDTaLGTVV5XCUlyE4JAxHz17EwhUrcb2sAgZfM/zsNgE5iT/42c1ITGiEB0eNxtCBg+AfHiaBg9Qt6NO7it9TmyjOrxUOqr9Kcf7sRbRv3xKxsWECMJKNr5h8fylJtSpDgdK6pF41XxTJgIG/P/20AitWrEBRUZHMScVFRQ3KJLLk2LjyGJSdh8fpQKTVhMceHI52SY1gJ0BjssLPZBXllsUeCF8/K+oNtH+qRUF+Hs6fPifBokE2KwLtVoSGhsAeFo2AqEj4+tvEtsfL6RblhlO8pHlGStnodHmjqNyJ739aijXbVmPS449i+B3DBWDbt38fYmKj0bvfQGRn5YM2QxzTebl5aNO6tWy06KtNtQobBcwccbnrUFJSJnZQ8uwZa+B0lcC7vhJlJdWIikiE1cr1gDJ2F8rLK2WzHRTki52bf0ZMuBFVZXmIjY5Bt559UVIfiIyCesQnpKCspFYUUrSUqizPx7ULOzGwXwcEhqTgepk3iitq4e3xINgWgAN/7sD3336EWqdDwHSqQBXQxLW0Hl07NEHLhFhEWP0QyOB2XzOuZOWgoLwKfj42mI0+8qyzURBosyA0wF/Y/Fa7GQlNEuEfGgYvHz24shJ52WkoyL+OoPBg2EL8BfD1YqngMaG4vBbbj57FgpWrUVHNjA8z4qJikJeRifgYG4b064yWcdGA1YaARslwWxuhzGGBweiHwBA76F9eVlQigC3nbMl/4JquWQcy94kh32Sh0qaCmTacBzn/suHOcViQf0PWYc49XN9z83JFcSF5MSQeWNQ8LLWZl7dkM+3esRXnTh6Fp6YUNhNVm3UIDgoAvBmKzfHD1YXkCBPMvgbYA00IYNaHxSrzea2TFpJuWbcdBMe5VrHWpK0Jvc19fMSujsQWB1wIiotB+56D4PKEwlluxeKFy3H0zCH4+iv1DxvtyhrHLUokzjmcP28U58No8BbVUWhwEMLCIxAZFQm73Q6rjZaQtGdkCDTXavWH811FiQOlpWXSUOKapH9x/aJtX62TVim0ubTIDEELJJPFqjIsQHCC4dFGUc2xSc9GrDQVXV4oLStHdlamNPOoqBB7FlGNqSaVYkWrOlQCqVkM1ivLUNV05vOqanHZ+Grny58Vl9yQ9d5sps0kz0ez/9GtCzT/b6XIVkHK6ekZQv4RRYXNCl+LCrLmnMBaSKw9JbtAeYML05Z1KUH64hLJBhDiCtc/o1HIE2qPQLIBLZIAu90Gq90GHwKpcCP/dLpmw/hfFRWcc2WMWv20Jiv3FyqUWMAAza5HrKNEGVEvRCCxwBVvedWI5weffIMAACAASURBVDEMHt77H4EKvcnN3+H58bj1htBjz40ToOK35Rtw7PApBQBq7HTVRtFWCAGfOAxUXaOzS/n70uAn4UpTgvDzRFVKaxi9MSwghDp+RVxSjHqC77IHEyYxFVLK65/PIedNxdBns5gBuMpyRJ2zqmeff/VRRESF4acFv+HCuatSf7OxQ0IXB4w0wbQauUH1wKa+tj/RGfCqwaRqUH6WnhVAdRlrfe7fOIY5LoUJr9nPKja5BrI3WMso5EIAEs0qiMfO68S9l279ovv3601v1sp8b85drMEVSHWzKUeQic0qrpMupxMBNitOHTsuczQVmVwT2Fi3BQXDHhGKmV9NR3l5FXp3H6/mCgG1SB5T+ykWIBIia+L+UzW3uRbqDWTaSSkveicGDRyI27q0FqAiL7cAn82cJ7W9sklWFllsUuuWIjqQzM+VcF1NGaHv0/i+eiAv90u6HRLnBLG08SH4SEcBqlMVwMT3J0itq8K41xS/fmb+UEGhBUezluY9EUW5yy1qcr4va29eBDl3LxUWzf0Ux53VQoCE+yBFUhSbFA/zhdTYvnVfemtDUt9/8dq1a5+Ml157VGqEV1/8VNm96UqLW549UZno1lJaVgqfAQIF3Bfw/rM25zVko1//0gmZAthqNnfKMUBXYqlweDoLiI2uNPc1YidtMTmfu9X1EDWIWLuR5KX26vx68aWHMWBQV8z+ajk2bdzXoC5RTHA1V/HeSc4OWen1tCAm8MB6Vj0LJEmwRyPPheayoKtn1L68VsgPMr8o9otm8aUcAfhZYi/nxfWYDgWVqK2uEjKdo7JKAIoAq1lq8FatWuLMmTNiTesfHAZvkwUVjhrZg/LkSouLYLHZxAatpoa5Jcx20Jq94s6hsk30Rq/eh6nViIo8vGEj+uDVVydi29aDmPb2bLl+tKqiMrchh4WWi0a1JvA5lXmCIKdkhKgwddVrUsAYx5UoBTSyq35vdUcQ/g7HocoG1cLXCWhLNqm6brqyS7caV3ZpCoSU8aqN3+cnP4Rx44Zh+YqN+OKzHzTQm9WOem5vH9YDr78+CZu37Mf0t7/9x46hrkaS51nABQuG3t4Nb739ODZv2o/p78xp+Gw+CzpArMi29ZrriFIv8dwI/LF3JCoqu13InQLY6BZ+mkJBAdoKsGkIxdaBYS0EWoirWu4Gf0+ugxZ0zqshIdJii6jWdf0c9H7J30/4VsCFNtIKMFbEYf7N/z57C1BBRcWtCqV/vIBaT053e9F/RwcW9P2UTuZsCDS/xeVF+o6akOHWdUsH3+XaNoDyGqBKBYqmFFJqP2UxyGvNml49fTclJNL/1AEXDXSSY9T6oeqZVVkhCvhTtUcDC/UvwMdNoEIqiX+Bin8cGv9+83/wFWiqsTyEnSOyQCXR05UBwsbWJn+dtXBT0qQmJL3JrE9IOgIoC4ZseLTFQ2MZ6Oif3mhRsj/NZ1AmQOVjqp5utXliYaxYEtzoqOa9MNc0NQYXc27M9I2F+JBrIVP0sFcFh0LydXWFHiYlx6sBmqK60EKr9ImEG1sWJFwYpSDRw9jIiNEma0FUNY8+AQ0aJIeKdaCrVvhakWhrmzO1cN8MMBQUWCtElOyMxQ3l0npomPpdfl+KQcmDIPNKLbi8blIMC8ijJlTVZFaKF567yPI05piSwav3Vki4khjKxkhC9NSxCztBA24UisNigAuLUqGIbJOgBL3jPS5VRLj4bxbQSknBv8kGHPLgg1IYqEJYMWvYzCDYQOaeBAf6GGUjSmsk+sxTfcAi3FlfJwUmN/rCqIdHGrVUNBCYstosiIyMlOYkr8W1a5dx5uRJ1FZVoknjpgJW6EBFYnIyzHYraqorhaHLBkJUdIxsdvleyt6HhbyShfI6/xWoUMwoFr1ih6DZDjlqlJqCY5aBiUo1ItwMZSFFdioZjbXVKC0tQnCAXUJMq4pLcP7UCbiry4WRpTc5OH74OilGySz1Mcox+vsHyOfQwsiP4Xi1dYph2HDf1QLHP8y2ELmrPE9KTaOeUyUb5HjifSjIzxegIiczU5QpvXr1gq+Fxa4CKsjglCBF8QN1wsutNjgSdyEsDqVAiYiMQmxSW5QyvFS8kVWQoz5HGAxuuA30vKyH2elE7vkL8HbWSqPL16IaEbKR93ijwlGL/OISNG7WDAFhYfC12GAyk1GqQBvZ7FCH4OVCcXGhFLecY2hhRXambB5pO+XrIyxYvUhXKiOOW49Y1hQWFUvYqsfA/BjhUMkGZs2KH9E8KREjRo5CWHikMOvZzA4KDkE1rae0uUr/TF4bMmdF3VHCMG0LfGDApQsXsGXTZrwwZaqEtVVWFuHc8b04eWAvSvILRXHj9qqHl68bpWXcVKqNMZUm0RGRYu0RaLcjKS4WkaFh8ifEP0CAOj+bVQrya9kZAhjwXpYWlyEvJx/h4RFo2qQpGjWKEd/3+lo3WjRvgVqHE5cvnIPF4itAhT0gUJ75amctzly8gLXr1yO+aRPxGw6LtCPY34aklNYITWgJjzUM/kHBqKupQVZuPuq8PcjOzUFBTi56d+mK4pIilFZVIDDIjrycHAwaMBCXLl5BSEgomic1V+GG3Fx43Dh1+oxcr25du8u9XLNmLT799GOkp11TTSXOPpR2c3PIuU3bJNQbuJEDooICEO3vj8jwUISGh4jdTHBAiGyKCazJc1lbLeHmASYT4qICERURjABbCMoqXUjPy0dRVQlKKx1i5UOFYEhoBKIiIxAWHARvjwu1FWXii3w5IwdfL1yM86kZYunma7EgiL/DsE6bCbFR4Zhw7wO4Y/AQBEVHgmZsRrAppr4aGlKaxLeiugoF+TpQ0QJxceENQIXCtbV8i7/UGFwDWNhrYDeZ5G63WB1dvHAJP/+8Ert37xbgkfMG51bZuArozcYmbZ8scg9Q50BKdAjGjx6ChNBABJlMsBr9xFKGLH6bfyDM/nZ4vL1RUevA+XPncObsaYQEBknIIt+L822jhKaIapwALz+TMJVrSqtElcLXuT0KqCGjtNblg0qnF1auWYMfVy3B8y88g/Zt2+L8xXMyz9Iqq0WrdoiNbSwgcXp2tmyuGlNVYPHDxQsXBRhJaNJErg3VVzU1LqSnX0dpaSUKirKQlXseFUVp6NG9N0ymQELz8PIiS0xZGDmcXLc92LZhOeKjbXA7y4U52Ldvfzh9o5FR6EJco2SUFleLOsHb40RVRT6uXNyFoQM7IyA4GXklXiirdArrNtBsx74/t2PR959Ks5lrm6OGgKdq2nPtTWkSji6tUxBl80O4nUozM85evYa0/AJkpOeL+io8OJATPfx8fRAc6C8KoKCgAMTGNkJEVBz8/YNhYmMNtSgrKUDqtSvw+BoQFhOKILsVvm4CHX7IK63BL5t3YeXmHYChDhazEVGhEbienYXkxAj06d4GzaOjmNQL/7hmcFvjUem0CVBh9feDr8WESjbUaSuoMcPqNPIBxxGBAN7zqkoGd1dLo5M1oMVqlnvMcy68XiTzDtn9CqjIE1s/qg/4vnxelFe8l3jA1zvrkZ+Tg93bt+DM8QPwdjtg9zPA30aCAln8bIby3H0FxPOzGGEL8BV1DZsxbBpxjS0rpe0Waws2iX1ETWEU60gfqdVYy7EmcXh7oVW3rohKbAmXOwSlecCC7xbjUuYF+Nq5zrGWdCnFBweOxoLm2lnlKENFWSlMPC42TXx94UswnI1fP7vUJiRacC1mDcB1Rpj99R5UO2qkUcbroDb59VI/1LtrxTaLhAyDgb7OHslBslptEopNdV1gUADCwkJRX18LP4sJIcFBovgjOEOwKCMjXT4nOCREWdBQ+ajZbwhQoci4UqtwLfbxqPBVpTxWliyiVmPN51K2JQqoKNQAf19pViqGoG6FejOo9P8NVBiktmZd/neggqAeVUYcDwRzaFHJUHDWfqwT/wpUsI7wgt1uFaCCuUKs6cqu5MoYYKObSlLeF2meuBi+6S1qCI4BaexLRpxSk6gGgGpO6F/StHHTB98Hw0YNQKeubeQe8P5lZ+YJ6HCroqL3gC7oM6gb/ANsSoVSUIytG3fjxOEz0rSY9MwYZf20fD2O7D8h479P/25/eU1RYQm2bdiLIwcJZHjh8efHIiomHEU3StEoIRpXL6Vj3tfL0KZDMoYM74vQ8GA5XH7W2lVbcfbUJbmvKa0SMXh4H3ktz4318rGDp7F21RZZD3SLDd4DknJ4PQYM6Sl2VgGBdvl5ZnoOfl+xSd5j1P1DRcmir2CXzl/D158uarCvkYaqjw9CQgMx5uG7EN8kVsYO5wCOL96nHxeskvF779jhyEzPxqyP5jU0tF6b8Zy89YfTvpbxltKqGUbcPRCxjaJUM7WqGrt3HMK637fJHoYZDqMfvB0dO7cRuzfOSbwnq3/ZgrQrmWpsMfJHa97e1q0t7h83EqlXMxEdG46AQH/5nEvnU3Fo/0nccWc/hEco5m7B9SL8umw9Lp+/KgVoZFQoRj84HI2T4lUIeHUNDuzYj9nvfwVHbR2imiTgw9nvoKysEsOGPi3nm5TUCNNnPI0u3doKIMKf/bB4NT788Ds5/ujocHz44VT06dtZ7GP5GloGvfX6J5jx/svoP7BLQxuKjb/NG/bgel4hHpwwEump2fj0g/lSv6e0SsK9Dw5FXLy6TlVV1di+eT9Wrdws15Zj8aFHRqFNu+ZyHNwXXrqYhp8W/4HcnAKtaU6gR9nD8np179kBd90zsOF6ECz5eel6HDt6HhMfvxv9BnTBgX0n8cWni2Rf8db0p9CiZVOsWb0Dv/y8Bc2TEzBm/DA0adpIyF+VFVVie7Nw3q8ChpJAMmxEX9x5d38EBwfI83flSgYWzf8Nly6loW+/znj8qftx+VIaGsUz48hfmtGnT13CvO9WYtToQRg8tEfDc8qf/fLzJjn/u+8djJ07jmD2l0vlWe/UqZUoL7Ky8jFj2rfo2bsDnn7mAVy6lI6mTePk+P5YvQODBncXW8AnJ72jKUJuEkT4LPfo2R4TJo5CfEKMPJfcK27ZtB/z5q6SPdknn72AZskJ+OLTHwT0eW7yGFxLzZb3b9YsXqq+9LRsfDlrqfQg3nz7cYSGsi5RX+npuXho7OsNPRe9qernZ8LUFyegV++OMk64Vz918hJmfb4EeXnFAoZQqfLc8w9iyJBuAl7zHl65kikAyKlTl+W/x44dhtH39EdERKiMGypNFy36HZs27pEMlqSkBDw7eSzad2ypALyqamxauw3zZy2Aj6janejRuzuGj7kTKW1T5BzLyyqxcvl6rPhxPZo0bozMjHSMmTgSd44e1HAcly+nY9YXS3HyxEU57wceGIIx44YhNDRIjiMr6zq++vIn7Np1DHPmvInbOrdquCa0bvxw5nx07NQSw4b1wg9ip/SrMN/Z56E6X79Ok6eMFTUGxwrPl/eX1/r4sQt47PG7MfGRu7Bu3S68884cGbOdO7fGu+8+jbS0HDz22Dt4991nMXhwN5w6dQnt2yfL+k3gcc0ff+LTTxbL3vHtaU9ixIg+WLjgd8ydu1Jq71demYg7R/YTAgF//8KFVLRqlYhlyzbgqy+XYv6Cd9G6VRI+eP97+b0uXVs3nF9VVQ0+eH+e2Fk9NGEEHn74ToSGqeuSkZGHWZ//hK1bD2DxD++hc5eb14XP+Pvvfy+vG3FnXzzxxD2SIajGUZ6oTnbuPCLrnyIl1kldQkCZdQdJlQLAaEeigxb6HlkAH50UqQVui7uBpnpQvSCdkKveSQcYGjKJtFwj9rj4+boNmSaHa+BeSd9IR4Ok1aeAXR2I4zp05m/WT3wP9v90oOXmen1ThcDvKUKk5jDylzP+q6JCVy+qPoACmXWAgS8T9UmDNeHN1+qAiSIbK5WmrgppUEBoBFMjN/Da162qCr221r+nAxEC5t9ic3irekT/2d+2g3+pW/4FKv5ydf79j/8NVyCJ7GWRq6pmtpLH3ZRfKVBCy2mQyUSTaPl4CzNCl90qeZTaCOmoMH9XLIM0No+8l4YUNqgrbvHYFIRYZKo3w7yFHaQ1AhVrRm++a5ItbaOhv6+wQ/Tmu6500D6T7y+MBQkPU96nbHTKhKaxDRQSrJgK/OI1IYAjE6o0jdR7KObDzWKYEz2ZO3pDX6yrtPAhmdxv2QUpNFdN8hpOIf8pE6Lm48gJkpO8sPmF9a4kj/rkxslcmABs7nLjKF0RNSJ5DfXQHgI7vDa6fO1WL0/eV2ESCGNHMcdEni8sPG9hDenghx44Jz6l4t2qQoIk5IxsH7L+KNcja5/WPa46yaaQjIr6Wu1v1aAfOmZMA1ChLyg6Y4SM2cqycmH1SAaJ5rFJ9o7F6tcQmqbLGHnvyCBkU5rMHrI2o6K4cKtrxjDjo4cPobK4WICKBkUFvJDYPBkWWijALbkENbVONG2aKP7h8n4OR4OiQpfVi5pFu5cqusQtm3hRSfh4SwCdw1EpYBBBBDYplNehAgT0BZYMwJpahwqqLC0S1m49z72kCBZaPNHKQsuE0OcZCYGThdFHNpjSxJAARKsoQRhey0YMx7AeOKaDFmwC6Mx/gkVKukl2j2D78j7SlCi6gby8HGSmpUswc8+ePRARFa38WLUcCo4bFiXV1VViyaOUNbwW6tng8dAWqXFKR01RUa95zypbBF4/Lz7jBtqWAcaaapSlpqO2pJhPHIwmgzQW2LBxewwoLK2Aj58NLdq3Rw2vvzebDSxUGVKqmkSOmkqkp18F3E6x+pG5pL5ebEk4llTBBAk4DwwIVMcg4eQ+6llnsG2tE3n5BSgqKZPPJSDEe7vu15+RnNwMd44cBXtgkDRF/AOoYggUppiSySqWCscNQQKORSqKmJ1CP2A22i+eO4+tm7dg6vNTBIRzOEpw7cIxHN+3GwVZuYSA4DG44PGuQ3klZdpGCf/zcrsQHxcrFmZsjCXFRkuGRnhQCMICQxAUHCgNG9rGZuVlS1A7mxPq2Dyw+/sjKCBYGM78E2ALhNVkk2bQpfNnxNqAzFdaOYHjwMuAg0eP4OCRw4iJi4XJQuApECEBdsTEN4UlrDHKPWaxqaqpqkIV1wGrGWUVZfKcifUTVSWFeaivq8b1vDwMHDAQp0+dQeOExkhpniKNPDaxaWpCCypaxXTp2l3m26+/+hqLFy9GRTnD0wgXeYlnO+cxzgeSXcP76+WCv92CZjExiCWzOSwURrOPPMe1tS65ngQf+SzR+okMsfL8HLRp0RTtWjVHRFgMcgsqcPLiJZy7dgHpWVnIzS9ESHikBMKTEUzLrV5dOyM6JEjYwFkFRZjzw4/Ytu8gCAd7G40IDAqSTYDZbkJIoD/G3DUaD9x7vwAVvJa0oPonEydRVFRXIT+vGBfPXUK7dimy6dAVFf8dUMEFSZg7wgZWuTGpqenYt28/tm3dLuw3jkE+AxyTegAesw/4/BvNVllPzAY3WsaFY/TgHoiwmRBisUuQttXkJwAox7kfbfF8fVHhqMLZc2dw5twZaahW1zjEkiUyOhod27RHyw7tUFhZBrPRDE8V8ynMsPjb4eVtEUTd4+1BtYumb2as3rQBi39ehPET7kNsXLTM4a1at5MA67z8InTt2hMZmbkoLi+XuY0h48wAYgD8xYuXEBsXg+DwIFHyVVe7kXrtOhxVLhSW5OJGUSrSrhzD7bffDoPBRL2lAJ5slLD56wJZil5YMOcLBFg9CA+xIMBmxIABfWEOSkTG9XpExyShuKhGGpNulwNVFQW4en4Xbh/SFfbAZsi+4UZZJS2aAJvRip1bN2PFD7NlreOcUV2rwmh5jznPhgda0adTaySEBCE6OBAmXzMupqahoLQMR05fgsnPF717dkegjRkyNaiprJDNJVlwAUE892B4uQ2wmn0RHGBBoN2MkpICVDrKEdskBkEBAfClJs1tQnphKb5Z+it2HDkJL0M9goPsCA8KRXFeHtq3ikeX9s3QJDIM8PNDcEJKA1DhbbTCbPOFj8kX1eWVsFuYbK2IK7XuejiF7KCAed4vqlOcNVQ4OpRHvdUE2gvpQAXBjLCwcAHMCFQYTVy3zKJUUuo8AuQq+JhrF0HIwtwcbN+0DqeOH4DRQGazCxZfH9htPrDbLaKm8HL7wGT2RmCgGW6uEbTi8CFDukaCULnGcN3lnMFMCRtVdGLV4CVEhypnNUJi43Fb/37wCQxHfZ0/sq6UY/53C5FXmgkfM+tMpVryaEolehcqhiCtwxisXQqvOjeMBOZ5DlzXfKgGVEo9qY24cGuMb1mPGqxKbwZ/8/t8XwHdxPedDXSyjCVJSjKQmEvF5y0oOEDAZs5zIcH+CA4KkmdYBypo9cavkNBQAUhYL7CpoysqWFeLKtigGLSoo2JRqTzlj2SUqRrz70CF2G1S9Sl5WX8FKviZ+ob9v1dU0BOUTN+bigq9/hOgwsjxY0BZWbmsTVw3abPDNZpWZDwungPnc86NbBDJukcagI8Pii9mS41FpQn/FisbqeeVkkSv0VnDKZCCIcFaRp9H9+lX91nqbU090W9QN5SWlmPfzqMICw9Gx65t5Jh2bN6HzWt3ov+QHhg0rDcqyipxYM9RaWh3791JrukvS9fiysU0THpWARWrf96EQ/uPY8CQXgImqNcck3PqJq+px68/rZcm+mPPPYjE5o2l2XvtcgayMnKQn1uI+8aPkFpz366jslfr0fc2+Z353yyX+/Dwk/eJNdi+nUeE+MNjCQwOwJZ1O7Fl/S6p7fnssUblv3v264zhowfAUVmNA3uPC7mga8+OyErPwc9L1iImPgo9+3RCSFgwtqzbhYL8Ily9nC5rDutwpQaox9MvTkDzlKa4eO4qzpy4iJZtmwtownP8Yd6vCAkNwj1jhiEjLRtff7pQxi6fsWkfviD3duZbX4vV3ePPjZGcqT1/HpaGaK/+CkD545ctAliMvGcw+g/pjoy0HOzfdRTNWzRF+04tpfk++9MfZN0je5tjn03Hbr064Z4Hh8kYOHn0HK5dyUCXHu2R0CRWmnKZGbk4euA0mrdogtbtU5B2NQOzZn4vCqIpbzyJqJgIHNx1ECcPHkefIX2Q3K4F9m3Zgy9mfgtbaDA+m/u+NCoJVJCgNm/hu+jctQ22bt6PQwdOYsIjoxEVHYZPP1koDddPP3sJI0b0w/btB7B9ywHcPqwXevW+Ddu37sPO7cfRsVMrDL69KwoLivHn9oMCGsU3jsXYCXci7Vo2vvh4kYzDyS9OkGfgz22HUFXpQK9+t0mz9udlG7B101488/w4dO7WBiePXcDRI2fQrUd7tGydhBPHzuPTD+c35LRIlp6PD9p2SMakJ+8T+6dtmw/IPEFQgASIWR//gOraWrzwykRpNBNYsNn98ODYYUhPz8EH78xBWEQIJk8dj4jIEOzdfRxpqVkYOKQ7YmIisOqXzfj1580YekdvjBk/HJUVDmzZuE+AoL4DOuPa1Uy8/eZX6Nq1DZ5+bqz0FfbvPYHLlzIwaEg3JDSOwb69J/D7r1uRnNIE99w/BPl5hdi4fi8uX05Dv35dcPd9g7F96wF8NWupPBdt2jbH1JcmICszD2++/iX69e+MZyaPlWfn6pVMpKVmIzU1S86BoPukR97WlK43Vaw89nc/eE5AlbV//ImiolKMHDUA4eHBWLJ4DZYu2YAvvnoZySmNMevzH+W9n33uQZkDCArt2H4Qnbu0EWuoQwfPYNpbX6NHzw5yLJ27tMbyZRtw5XIm9u87ofq4sm9RKoH3P5wsv0OQhnZI/DdBk5MnL2LG9O9wo7gMTz5xNx4ccwcyM/Owdu1uNG4cI6BFbm4hpk+fiw7tm+OJJ++Ve/jHH3/KHD5q1AABi2fO/B4Xzl7F57NeQ1KzBKz9YwuuXLiK4XcNRnKLJPy+7A+sW7paLEJfePcFNGudjEO7D2PPrkO47yGO6Qh8+N63WPj9Srz65hN47Okx0mT//fcdAtAMHdoDOTkFmDbtW3TokIxnn30QBQXFWLlyM2JjI6TxTzvEV176XICxNm2SMG78cOzdexx/7jgiwMFjj9+jgIrFazB37i8Nqirdfvypp+/DQw+NELDn11+3yucStMjOvo6XXvocI4b3BnMu1q3dhWnTZss+lnZM7777jLzm8cdnYPr0pzBqVH8UFpbIsXFuv//+ITInf/31Mvz44zq8O+MZsW5avHgNvpm9HI8/cQ8mTRqNvLxCeU18fLR8LoGeefNXid3T/Pkz0Kp1Ij54b568d/sOyXIs+/aexNatB3H8+AUMHNQVzz8/Bvn5N7B06QYkJERj1Kh+uFFYiuee+wgRESHyuokTR2L3nuOiNjl2/DyaN4vHjBlPS53z888EJoGxY++Q6/nsszORmpqr2d6pfFRdEchaTrclk76W1s8Ssp1GwBVymChUqHRUORi6OkaUE1r+lrKFkyJH+ggNlnZ6wLnmoqIWU5W9oIdb/5MyQHZ4GrlHGibwwtktCoznV5vBJB2qNUNI1Rp4Im9/0++6AfDT7cqlb3grC+GW32cfQvp4dBDRsnglMFyABwVU6D1PVc6p3p/+PWXtrr64nrGeVb+n3lfcHjTrJ+0HfzGh0t9HrxUbmqgN7l7a8UmNqJT42v8baG9/19z/C1Q03JJ///G/5Qo081UNSh3NZIEgDUnJBtA8NZWJnBS1unUL/9bRWuUJ+dfgT9VQZwHLyc4gnvic1WQTpE1gOvKoh2PpMnA2wnUbKja6ZXLQm8PSHFfSaglT0nxxlRpASQv5c25WdKUHGXv8ktAhhk3JxKVmT/FSlM0cCwRlpaRmHW3DJjZVDHGkd5/aYCp7JwXg8LV6qCJBDx3FFtsnjbUugITmrar8Vm++dwOyo02Kwtx31snGVP0eL5+SCfPacSFUUn21mVabNxUgqYfZKZmjQrr5pW8G+T2euwo9VF6bukStupqbFgXcKNm1FjxYp6Tl/NIRauWXSbRcU71IVoOS0av8BcrGnaitqxEVBRu2SHh/UwAAIABJREFUtH/i9xRQMVbOkfdYyWbVBpnXnxJA/ozSf17bqspKVJZXij+vhHt7sYmv7A24Ged5BAUFCYOGGxQyrGhlw+HIYyy4nofDBw+gvLhIWT8lNIGbihZaP6Ukw+pvh9Go7Ap4jek5z1BHNl/4nrQtIZDDhUttcG8GclFWz2NnY5r/ZpEqC5UBcty0qSLooRZ9pbgh249e4IrB4EZNdTm8PXXITb+Gwtxs+HoBZrFmUE1/nqveBOfYqRUfWErLydb0kzFI66egoGBRnLCJxNfozRIdVGOuhYIJxYxECx7js6Xswbip5/WuLC9HSWkRMtPSkJmZgaSkJLRp1xa+IiEmm0F5/ioZsxP1ToeynVHKfRk//FkoWfwpnWj3KcevAriVN7XMFVRBGPk+BhidNajNzUNZdrYEsxl8aBnAyG1623ujpKoaKe06weTvD7eBNmAWyRagLRTvI4GJQ0cOID8/GxFhgYgID1djS1NVkNHLe+R01siYiYiI0AAkxaYUhQXnCLLSGO6anYuCghti28Ofr//jN7RskYIhQ+8Q0Kbe4yXqA9pv0W9bf874mRyD/MPzrXJUoKKyXPznXc56XDh7Fju2bccbr72OxKRElBTnI/XiMWxb8zsyr6bBwGYqOfg+9QJUUIlh5pziqkd8bCxysjJlQxkfFQa72YLggCCEh4QiNCQE9gB/CXHMyctBbS3HgEV84HkvmJvCsULvc+aH2Cw2+Bh84aqrxdUrF1FVWQ6evq/ZLDYaBqMJa9ZvQGpmGkIjwuBr8kZkeKAoKpo0b4HQhNZw+4XIc1Ry44ZYctUZPJJRUVNeIYqKmNgYVNVRxVCKY8eOYMjgoTh3+ixiY2PRIqWlPAsMpOZoJoCRnZOLPr37IC83H9OnT8f27dtkDpB5mNJXTX7M8aPyHRhO6SUKhnaJiQiSeduFS2nXUF5ZLSxaqn8GDRgkc1NG+jVEhoeguuQGunVqje5dOiA8NAbX0vOx78RJHDh+QBpTefk3EBkdix49eoltnKO8HN1u64jWzRIFNCp3urBuxy7MW7pc8iwIHLKRHhAUIIqKAKsfRgwYhGeefAoBUREKzLjF+unWuoHPcWW1A9nZhbh88TLatk1GfHyU5NHAo4VC/l+sn3j+OihO1Rb9pnNz87Bnzz78tHSZ5LlwDHINFOu5euVbbTBQOUeLNVqguGDz9UJKTCgGdG2NUD8jQvwCEWC1wW62yvn62eyinDFZLBJOz+ySnNxc5F7PR2lFGcorKuX826W0QqPExkjNy0TzJknwrnXB4PYgJCIcPiYCHSbUGVxwGkxwelmw+Ofl2Pzneox96G6kpCQhMCAELVq0hbfRgrXrNqFb154oLq0QiySuUfFxcaLQEEZjeblYqoVH06qPoaAEKm6g2uFBfmE2yipy4HGWIyQ0RNQIBm9mDEGOtaLSgRoXLRF8sPD7ObCZvXBbh2YoL87E4EG9EBrdAtmFBL/jUVbhkgYgk1RKi3ORfnkfhg3tBr+AJGTkO1HuqIPF1wi70YZVK5Ziw+qfBASS55/qFbXoKztKA9CpZRLaJcYjNjgAgTYbsvKvo7LGias5ubh6LQ2tW7dAjy5dERsdIc8+N5T24ADxgzbCF/nZ15GbmYUrl89KfkOLJGZX+KBxYjyC/APh5fJBTb03jl5Oxyff/4Ar2bTLccmzG+ofjLKCfHRq0xSd2iUiPiwE8LMgKD4ZXvYmqKgjc98PJquvNPRqKh2wW22iNCWoQJCijgG1BCpqakSZxuYtwTs2QznWLDaL1CT8EuuniAiEhoYJUMwwbSraOFdbTLRtrEaA3V/VJ7QoqPfAXccZ3wsZqVeweeNanD93Au56B2xG5jP4IMCfwdFmGDzMXWI2mgEugqXVtaK85Hjm/EjQgkx8u8UkKhw/2lAwMJhWk1UVqPc2oEvfQWjatj1qfcgytOD88QwsXrAIFXU3AF8V4Erllp7F5tZqHSqI6p1VqKE1hqNGlLZiySi+VGQr0CpSWVHo9bNu08K8mIaaTqtnGzbBmlUKQXhRqQqpgYCLRXKF2PgSNYrVjNCwYLRqkYLY2BjJzmBfncrBa1evSg1GRYUQF6jepApYs8qjwo8fS8WyqIprVR3JdVvuMdeyerUmGjQhl4BON/Ll/lqtSh1CsIC1tl4LSS2jAzLa8WRkZEj+FseEyWqByeKrPOq1z+H76bWpgDWSF3ATqKAKWhQVzGTw8kJhQYH2+2q9Zt1i97eKlRMMvgJU3LiQKbUbCSIeN72mdZU475GynlWZdMq+lMxhsU4heCOWldrex63yF0gSev61R+EfaMOqZRtw/vQVIeLcdd8QdOnRATu3HcDOrfvx9AsThKX/67J10qDn6tR/SE8MGdEHl8+nCoDw5JRxYr3424oNOHXsPJ575RF5Dd/3zMkLcm79h/bA4GF9QMXCwm9X4InnxyEuPhqrlm/AiSPnpNZ85OkHkNwqEds27sGWdbvlfj844S506tYW2zfuQXFxGe5+4A5pbn/5n/lS5xFY6TugG86fvYJNa/7UbKWo9VONl5feekLUGb/8tA5HDpyS+/rMiw+jaVI8fluxUcCBqa9PEuunZYtWC4giRCotDJn1T5fu7XHP2GHC/P/28x+08eTEi28+geDQICyZ9wtCQoNx94N3ID01C7M/W6SF2Rrw1vuT5bl4/82vRNlB0OfU8fP4ZekGqTHvvGcwBt7eA4f2nsDSRavx/KuPIKFxLH7+cS327zkmte4jT90Hq9UPa1ZtFSBEKxfkXAhKPDB+pAAo875ZLnvAlm2bYezEUQJszpm1FIV5NxAeGYonp46T9/vhuxVIbJaA2+8aiBOHT+LtZ96CVexoffDB/I8RFhWGhV//iAOHTuCL72aioqIKQwY+jkcmjcaLL08UhcQjD70uz8udowaI8uD8uasYO+YVbNz8nQBJUybPxN7dx5DULB7T3nlG1umF3/+BPn274KGJw5GXV4DPP1ooY7FP/y54YNxwaa5/9ekS9O7XCSPu6o+jh89gycI/ZPyMvncQhg7vjQN7T2DBd7/gg09ekGf2u29W4Mypy6KOGf/wnRIYPUtjirNuJ0OZtesLrz6CNu2aYdXKLVj3x06ZPx5/+n706tsJG9bswvKf1mHIHb3wwNhhSL2WJe9NwGThvFXY9edhjBk/AiNG9sPO7Yfw7ezlMmclp8RjyosTRen24vMf4ePPXxVwYu7Xy7Fn13F59t5+92lp6M6ft0qAoyeffgDHjpzDRzPnyf4+KiZUro+vySiqBdZzz099SKyfXn/lc1Fhjh0/HPfePwS7/jwitju8723aNMPLrz2KnOzrePWlzzBgUDc8M3kMzpy+jDde/0Ku2W2dWovqgvu9Jx57R+2JtfBgPutUW0x+fhwuXkjD1Cn/gZ/FD3373YaRd/XDwYNn8OPidfjPp1PQomUTfPHZEpkHp7wwThrlUyZ/JESH5smNRWFD699JE6fLfoFZDP0HdBHFwbath2Tvy7Gu9nvAgIFdMOWFh0SJ8fKLn8lr2U/56OMX0KFjCyxY8BtWr96J7757S0Dnd9+bhxPHz8v+65VXJmDQoK747vtf0b1bWzRvHo/PPl+KLVv2y3M26dG7MG7cCKxfvwuHD57GlKnjkXYtCw/d/wz8zCaMHD0Yr70zFedPncdrj72C+yfeh4eefRinDp/E4w8+h6paF+64ZxhmfPQyzp6+jAljXsL6rQtEOTX9nbk4dvyczCsz3nlKlArfzlmJFi2aolPHFvjiiyXYuHGfzEFzvn1Twqb/859FWLvmT2n0v/7GJAFl3n33O5mf3p72BO4QoOIPzPv+N3kdVe68zgydX7Lkffn7lVe+wPnzqVKf8DW3394Ds2cvh7+/XdQKG9bvwYwZc+VZ6tKlNT6YOVkUFZMenY7p7zyJYcP6YNYXP2L58o2yvx07bhgmTx6D06evYOLEt/D++5MxQgMqZs36Eb/+8hkiIkPx7oy52L7jkOxHXnl5Iu67bygW//AHZn+9DPPmvYO2bZpj5gfzsWbNLtw5sg9ef+NRsXAieMOvTz6ZKkqSzz9bIr/DBXrhwnfQsmVTzJy5AKt+3YrRdw/Em29OwsZN+/D2W9/IPZw9+zX06tUB3875RcK6Wee/994zGDmyLxYsWI3Z3/ws7g9ip9aQ9aLlJ2l2W0KiJJmY/SSX6vmINZnUCIrwy5pDkS6pZFX9PKlZxMqVFoGK2Kz3h6S/pudPaf0+1rFCwGVvUfppWkdJ+0t6gqJoUOsun0Gxlff2wemNAQ1bplYDixt6IaqPofp0qj2pChbJchWLa2X/JcHbtJnT1va/Wz+xV6XbeInLiJafwuOVHsLfnERUH1KrV4SArWUjaf1Qvof0A7RQc14r2bNqIKQOSAi0o5G+GwLJte+xTpL7omX66kHdch01srecrNZL/QtQwZ//a/106zb733//b7gCVFRIc18HEbSNNR8W8boXCZJ6+FggqKar8pfUG6jC7JQNiposJASNjV8NydTDcpSaQfkpyu9pSC/fh/8WP2QCJGxea+CIbC40BFOkvMqrpiGwRyYn7b+Vlxu9BVVzS2/I8986CMINkvLZVfJxfnGDRryXbGWZWMSLUqkF1CQmPjBSEAiaK76tymeTm1ROJPw3m91685xqBDat1bUxKN9Gvl5j5slmkMfKBj3BGF4Pg7K80XMuGpj7YgUFKdQoPdaBD32CU0FjDBFTCgiVIaCYhfxdfbLmZpTNSJH/aZ6ZPF+yr7mhYciwqGB4r6myYSNe84VVwJGedUFdNa+vutYqo4EBYi4BJMQ718VGDc+NrD4qKvh9ghZ1GDb2IWHySWCdlomh+9YqmyT66CoghZtdNplZTJOZyWaZCn5TTQ+yNtkQIaigs/7YJPXxUSHnRUWFOLhvL8qKi9C0cVMkxDdRGQQwIDE5BX4BNskSUACdUgNQNsn7RSayi8xGrXDVw9718cjhoX9PLK/EN74eNrtVNs70dZVrLiFwXIUU8OAlC7wCmuprK+HvZ8S540fgKC2GL8ek5iutWz+pZ4+bbh/U8TO4kIulDa2zvAVECPAPkJwCNuX5eTyfBrDC2yAND44FYR54sbGglDP8WzVE6AtcL36kZOQX5ufj8uWL8izf1rmLND/EC7+OjEP1vPK1TqdDGnFiG0FGAT1vjb7i25/YopPYOdzqV8l7p7JFvKW5DW83bLTNKi/H9WtXJfPCl00oPjswoMrphiUwBE1atgNbGybah/j6is1VdTWfW84HHuw/sBf5+VkIDbQjNiZaxobY3ThVpgk3gQw55zFHhEeoBod2PXhPOCdQqcJgcioEGK586fIV3LhRjGNHDqFjh/a4Y9gIxDdugrIqBwIDg8VTm2CdzubQFRUcwxyLpaXFqHRUSJi2q9aJs6dOY/fOXXjrjTfRvHkzlJUVIPPKKWz47RekXbyM+lqXXA+XlxNV1W4pwM20qqivQ0JcnCgTePzx0REw+/jIxjkqIgrBgcEwGL1RXlkuDSuyfIMDQ+Bv84fZ1yRNTKpveM39/YMkgF3UWHU1OHX6GMorSmAjm56KBJMVpRXVWLpsJZweJwJD/EFnjajQQATa/ZDcqh2adewDv7B4WGz+qK6sQGFxGVxGL1y5dhWZV66iVVIzYeX5BdLixo3U1FT07NYD586eR0hQMFq0aKmebaqxPC4JHk9Ly0C/fgOwe9cuvDN9BlKvXmVio1aYKbBQ2EACqrNhykBUbzRLiEObRgnwNxrFouRKVoYEOttsAbBbA9CmdVvJecnOSofFz4Sa4kJ06tAC3Tt3QEhQBLLzSnEhLQ1nr17Q1jUjQkIiEBkdA6OXAb4MNbaYJI+BG+LKOg+OX7yCDz6fhdIqh2Qo0Ec2ODQE1gA/BNutGNyrD16cMhXW8FDUCZ5yM6Pi1pqBU0JVbTWyMwtw+dIVtG1DoCJSU8f990AFJ2A9J8hgMAowWlhYhH1792P+/AXIycmRTYejmmoi2sMo4Je4Pv8QjOIzS6CiWVQwerRNRDDtdExW2C022C0M/LVIQzogKEj0acUlJfJM1ThrUVxajqpqh6iLOA9F04osNgZFVaWIj41DTVEprufkIjQ8DP4BUfCh7Nzggsvkhyq3Ee98+CEcdSWYPPUJxMVGobLSiYiIWASHhGPnrr0Ij4hAbKPGKK1gPpQFsdHRao+hFfeVVZVIz0pDQuPGMHiZkZ5WLIqKvOtZKKvIQ3REOC5evIC+ffsKmEmGenlZlTBfq+pKRHl3PTefEh1Ehphw8vhW9OjaEk2bd4Sjzg8GnyCUlrvEEqLeVYsb1zOQl3kMI+7oCZOtCdJya1FeXQeL0Rt2XxsWzp2D3dvXCFDBeZ9rusr2UQAuLacSIkPQrXUz+Ts6NEQa/bQPKa2pwdlz5yRonaGVnGviomOELe4b4CfZMQGWQBTmFWH/nt04fGQfGjeNQWx4EGxmIxKbNZGsGme1GxVOH/y8bRcWrvwDFdX0ancjJjJY7KlqiovRoVUCunRsjuggf7jMJgQmpMAYlNRg/WRmZpnBg9oqWi9xzlC1GEFQJ23+oEgiVHqUlpTLPaH1E9dLq53KGUUmoO0LAePgkFCx7srOzRW1HwkGYqNZVydB28JyZ1AwlS4uwMfLB2XFJcjNyUJebjp2bt+C0utXKf4QCysjgQpRUXA1cMLbxyTHyOBlExvQ9Nv2NQmAxWeWzWrWr/TCpiKoqLwc8YlJ6Hv7XbBFxKAaPnDWmHBkz2ks/eEH1Bkq4GVyicqDw42ZOML81oAKKkXddQ7U19SiqryCS6nyDyZQIWnfXtIcEEWFVlPrZAG3m1aVt1i53RIiKVWmiBtZ21Il6Cdrp8nXAm+jSdR9JMqwruFalRAfg44dO4qqggfKPJrUa6lSj/jzmSU4zmwR5oSJ6ljEcg1kF6lhnIo1KAQWhlxrGVoCOng0JiE8KCzMl/tls6lcEbIQGbiq1yV6nS/XQfYBDNPOEmtIAhW+XLP9lP2V5NbUKusnff8gntis0TXrJyoq6mprESBABdURHE8FDYoKHajg8XCNJOhK3/zC85mwmFReF/M2OBao3BPI2pfqYWUZoWxZxeShwSqWVE9RWXPO9zXK8TVvlYT7HxohgMan730n9TwB4WGjBopN0p7th3Hh7GVRMJSVVuDzD76Xc+K1bdQ4Gg9Nulfe54uZ8wRgICt+za9b5Hf5vuo18zTSkBuNkxrhoUn3SN364bTZePqFhxQ4sPB3XL6YJtfh1XeeFpXAjwt+Q+qVDNkL9erXWeypThw+i+2b9oh6gwoKsqVPHj2LE0fOKNtQTQlO5StrNu5bkpIbY9yjo+UcP54xVx0/g23v6ofe/btgx+b90vwnOMBjWTJvlTT8hdTEXAvx3PfgzrsHo+/g7ji07wRWLPmjYd547qWJ0tBb9N3PYv1EUIVAwuczv5O8MI6V12Y8I/MkgYoGxbHWlKEifPio/rj9zr44uPcEfluxGUNH9BZFRVFhKQ4fOInjR87iRkGJUoWLpZwipSmynAe0fiJQcezwafy06A/5nSaJcXj4iXulkfzB29/AWV0t4PCr7z4tOTZLvlshYFT7Lm3x65JVWPTlAtgJHjvr8Mzbk9FnWH+sXbkev/26AZ/NnSnrSq8e4zDrq9dx9z2DxRppzuxlMncmJsVjwQ8fyjPUv88EzP72bQwf0Q/nzl0VpcGmjbslj4IK0u49umPQkJ6Y+MhIYWt//tECudbdenYQoIL2Vf95n2oPleOhEwZ5/e66eyCGj+yHvXuOYfG83/DU5DHo1LkV0tNysG/PcRw+cAoV5VUNY1Qsa6lO1gLLP/nyVdnjfvnZD0i9kiXHTkXFA+OH4cCeE5g3d6Xcr+dfmoAu3drI6/7ccRjz5qyUf0956WG075Aiaottm/cp1rOXR3LPWIe2a9cCzzw3VtbUF579j9wfzk8PPzoKdwzvjd9WbUXB9WI8/uR9AuB8+fkSleXnY8QLr0xAu/YpmDN7uVhpUbmRlZmLaW98Lc/Ag2PvwL33D8WObYfw5Rc/yl6Vx/LCSw+L9dObr32JXn06CMCxZ/cxfETFjMWCdu2ay+9w/D/26DStQcjwb5dkJIQE2/HBR1MRHh6Co0fOYsf2Q9iz+4SyudUIZx9/NhUpyQn46stlch2enzJWbIBenPpxQwP3x2Ufy88mjHtd9mwvvzpRAI+vZv2ELZsPSP9Bz0nh3o1KAgIva//YKTZC3Aty7hn30J14+JGR2LLlAPbvP41XXnkY165l4YUXP5d9OPcybCzz96mu+HDmc7LGPvLIO0KqosqaOYbcT7NlzP01FdseVx0K83MF4B98e0988MU0nD1xDk/e/xTe/vgNjLhvBBZ/8wO++HAualxAVEI8lv76pVgPvj9jDj7/8jXQ6mnq1E9lblE24jobXzWh/1L7ejz49ps3xSrp4/8swurVO0RhoQMVM5jF4AVMm/Ykhg3vjcWL/sA336y42fvxuNGnz214550nce1aNh59dHpDP0cnYXJpI9gwYcKdWLdutwAVvBY9urfDjHefRmpqtgAV738wGYMGdcMHH3wvv8c1gADKZ5+9KADRyDsni3phxJ195DgOHTqDmR9OlnE4evQL8rkkpkx9frwoQhYvWo1vvv0Zixa+i1atkvDeu99h9e87cPc9gxoAh+nT52i1j7cKX+feW7Mlnz9/OlpTifHBfPz+23aMvKs/3n77cQnhflvLtli79ktZj1999UscOHBK7vd99w3Cyy8/jPXr9+Dtad9I3aL62YowoysQeH24HnA90/t0KuOrtsGaVvbDBm+Ul5fJGiokXiFAKmKv9A+kaa4UofyZkIe1m6z8QtSXml+UA4rq76m+l5Cjtd6KENIMBiGaKBVyvZCDz9+SUdF6kNp/6GuEuFzcsq5J//GfpOvqKqjenoDrXONVOL24lfxNbaHcU7Trxn6YRnDg91SPU8/T1XJaNbBGz6W61QpLfl8DUf7yAKgPaOiR3qrSEBcTPZRc64Pq56zfO75crpWHeTZ6lpXKwfkXqPgvV/rfb/xPvwJNvVUjW2+K60wwJX26mZ3Q8OBqEicuRPoDyYJJrGZEKqEk7GpqUBOkWN9ovlBsNskWQVMm6JOVhBfJBMoGrppUFICi3ocTFxkaUtxom5yGjSAZ3hI4xcVQvY4Tn26BQ7sQCVeiVz99xWkPRfa+9jsityQ7nIUu7ZvEhklNImpiVBOosOo5uYmdlQq7ZrNdbQQ1VFg2cFrOhJeGtgo77qZdlA4GSIyx9jqZqLVZVgAUbhRvYdOqsC4dMFIgkZyT2HYpViKbBaLYoHyf3ugSOKUQcAFGJCBKbaSkwVBZKZsFXhNhtbk9Cj1n+CM9ySsrhQXJxUkfH4KqE2zRNr/64iC2LB4i8wqQ4EZBKStqJUDbpeVVUF1xxxgCFVRwqGa6vqGgaqJOAzqkIaX5QgvjhwCMG2CQZ2VFJcrKywTxJ0jRKL6RFEe0avKzmoVpSNYfN6ZsFu/fuxulN278Bahgg61ps2T4Ws3wD7DLODMYfGRR9jaojWpFZQXqXSrrg+fJJoDOnldjX4FaajEmIKVUOTpQwfNiIUeARbIbvBmCbVGKCvFjdKO+pgJV5TeQduEs/AyAo7JMLB947/RATv3eEWSinRjvLpvOoqoRRYVFGPNsKPKLQIB8jh5yqYVpN6hsvFTOigIq1KZdVwPxfJzOapQWFYmiIj8vDymtWqJZ82Rl4eYxyEaa901C3lxUKqhAaWVxpeYTm80fEXHNERIarqlzbkooad9SVVIFg58RLl/A4KqFze2WUO2igjz4MXtAgj9NKCyrQpuuPWCwBcAvKESCtumrykedgde0DOG5ZGSlYc+uHbAYIUBFdHS0XEMCN8w/kCLFyfBXB6KioqSRo6vAeC5mk1GBSD6+dKdApaMG128UIS01DWvXrkGrVq0w8q7RiG/cFAVFxQgMpg+4RbMu155zLaCQhRzHd1HxDVFUhIYES6PrxPHj2L9nH956/Q0kNE5AbU0ZMq+expY/ViH1wmVUljngYzagzl2N2jp6bftKmCiBimZNm+JGYSFqqh2Ij4mAnUBLnRvxcY0QExWF8qpKXLh4EXm510UxYSPgVu8FX4MR/rTwsfrLnMJ51+RnkSBio58RtZ4a+Nl8YfM3Izo6Srz8T5y6hNXr1iOI4EQYPatrEBUaDLvVgqTmrdC+11DYIpvAbLVLRkVRaRlg8sG19FRcOXce3Tt0QnZuNs5cOi92RnabFa1atsaRQ0cQGBCEdm3aypijnQzzMK6lpiEjPQs9evbEN7O/xdw5c1HNgEanAnCl+dcw/yqgwttDIMeIts2aoEPjRITarIDRC9eLC1HnMSA8LAqhQaHS5OYcy6yQ0uIb8HLXI6lJNDp3aCOKivIqF3KLipGanYaigkL4GIwICCYjOQD+NjtCg/zFeob86FqXB0WVNTiTmo73Pv0cN2gRJhZ89IUPRlAYVSdW9O/eC6+9/DLMwUHMq5Vn9Z/qZ66TDmcNckRRcRVt2zZHXGz4/xdQQWWaHhDIhvf27Tskx+fkidNYvXq1NC51UJAsReZTcE4mHutr9IZHmNsG2DWgonPLBASavGH0scDPZIaVGTu+JmGkWWwqNFMBeirrhkH2LODNFj8VjOztC/+wELi8aSdlQMX1G7h64YIoMSIjE+BttsBpdMPgH4SLmdfx2rRpSEqJw1NPT0Tr1q3hcJDN7YUbRSXIys0Rq4WOnbshv6BMQEGL2SxWSGxyc22w+FlRWk5FRzkCAsJRcN2Bqqo65OSno6wiH8mJidi1ayeGDB0ilnTkIpQWO1BRWQOnp0wsdayWINRUVMIH5ThzcgtSmoWgTfsuKCqlNscGl9sCo5GNTw/S0y4i9fJejBzeBz6mOFzJrkSNPKNGWAwmzJ31JU4c2oG6uho4amoUq0vmWNrx+aK0wgF/izeuHt1yAAAgAElEQVQ6JiegVZNYxEWGSRO8upp1h0fUMLnZ2cLYjIhg5kdjRIaHITwqRPJwHKU1uHzhCvJysxEaFYwOt7XAjYI8eDz1aJoYL898bY0HV7KK8MmiH3HkXKpq/nq70Sg2AmbmhFTXoG1yI3TvnAK7rwH1Jl+EJ7WBJSwFFU6lqKB9k9vLg5qKKjWHaKGSJF5U1zMLSzV3SeqgipNlHfMRRFFhNUsGDudVKipo+xQaGipARt71fAEvZS6UsEpvaZjwDZjHROY/x5TByyie/NwgBwbakZNxFT/M/QQOxw14ezOY0ASrWYGnXl61AoyztvI1GMTmiYG3QXY77P52YeQzY4J1QEVVFUqqKlFnMGDAkKFo26kvXCYbHDDAWe2DvduO4JdlS1HnXQ6Xt1OeA6mXaAnAdU2ro0QVQZDE7ZYcjzqt+U3VsJcPbVRv5oLpDQK9QczQzQaHgltyEaWWY8YS61whIfjC5GcVxZ7JRLtLi6iCxCbL2yNNpoAAK1q2SEa7du3kGpDAkZGeLuu/1WYToJ5fBJgUo0/VrMrukGQWLwEqFCmGTfp6OGvVOi51WYNHA0RRwSY+GeuyESbBQrIO1O/q9aVspglUuNy3ABVmybgiUMF5ks2HvwMVuqJCD9MuKy0Ti7cAf38FjACiqFDEC2gZUx5YbVZYbX6iwuIPii7kNGSGkGxyU4mtamn+Txowmr2K2pKouleMtrRGPq8BAd4WrZth7KOjBXSb84ViS1N52m9IN/Qd2A17dhxGwfUbuJvWK2k5mP/1cpljdVtXggr8jI9nfIunpj6EuIRosYLi59/NrIa0HMydtVRpXMV6wo033lN5DR9N/xbPvDAB4ZEhWLrwd1y9mIaYRlF4+Ml7RZnQ4PPasAH1EiUGjzMpOQHDRw9CTFyk3Gsqjtik/+OXzQJGqcaLt+x1WrVtjvvGDxd2/D990V5q2aLfMeW1SaI4WDLvV7GhktB1rRnF6zps5ABRhOzedhC/r9yk7YtcmPzKo4iMDpcQbluADfePGy6WTZ/N/E7uFa/pm++rc37/TdV0Hji0h9hRcQ2QbD/ta+/OI3ItOA7ufuB2yQ2RTBC3R2yf1v22DSePnRdAVEh2ykcEXXt1xP3jRuDY4TMC8PAdW7ZpjnGPjpIGNT9Xcq88Hkz7aIpkkcyb/SOGjRqEJonxmP/lIqxYsAz+flYJ1r5rwt0YPmYkfl+2BmvXbFOKikoHBg94DLPnvCXM8H/6IvAwZfKHOH/+GqZNfwqDh/SQ9ZXPJ9nwb77+MXx8rBgypHdDmPanHxLIAnr06oixE0aKndIXHy+WtX3osN4YNKSHWMLppDt+LtUN875dKdZM4x++C+07pggwz/0CLZaWLVmDjLRcbR+tshvjE6Ix5eWHER5x02rl1nM4c+oSZrw9W46FNmCPPXGv7IW+/Xo5Tp5QJI8ZH0xGYmIjzP9+FXZuPyj3jns/3S6G6gXaOtntJAn9169NG/fi4sVUPPHk/diz66ioMgSMMRjw3JRxktXAJjAVOS+9qpQSb742S/ZnOlCxfdsBzPpsiZxTy9aJePX1R5GZkYe33vhK1BFPPHUfdv55GJ99uljmMio5Xn31Ucn3eGj8a5piTBELdYIfsy6olGGuBecP/u6OHUcw99uVqHE48cnnU5GS0hhfzvpJnsvJU8bh8qV0TH5uptrfGwxYtPh9Gevjx74m89Irrz0i9k9ffrEUmzftayA0qv6FF15+9REMGdodPy1dj8ULV8v58J7ffkcvTHlhvAAmx45fkMY0lQQvvzKroWGpg6XMW3j7rcdQWVWNBx98TWsqK109bU3FPcLjxujRAzBiZB80SWzU0ATm3Tl64DieGz8VH37zHvoO+b+M6dxC/LxiEyY9fjdOHL+AF178TMsAUs4Vam2AWGU9+8wD6NmzvQSY671hyaL4cD42bdyPO27viVdffwRbNu+X5j6vA0OkCVQsmP8b5s5ZqZrK0h8Bhg/vjTfemISzZ6/iscdmNPQSRO2n5TNMfm4sHn10lFg/vfve9zLoqKgg8EDLskmT3pF/DxnSAx+8/x02bOS9UCHmq1Z9ImPgmWc/wiMTRypFxaI12H/gJD76zxRRNz3x5PvKOcTlwuRnx2D8+OFY8uM6zJ37K77/7i0BYt5793ts2XIIQ4d2w5tvTcLmTQcwjUACINZOU6eOQ58+HUWRol8XjrGbQEU/ASqoRJk2fQ6SmzfGl1+9jLjYiH+es/edEuBG/9LnUL324Dp36/zInpuujlDkAbWmi7JI6x3p/R5dqSB1oEao5PyrHDVo5aw5tCgKoXzp9kgsKdi/4Jeyk9J6XPo6rNky6DmpJJmc3nQzy6XlgCJ5rdiP87PYq9NC0uX7BKf/5uzScA000FoHRPg3M6hkDfuHzZn0K/Ue5i0OKIpkrTp1t7rI8FwE/NHAA319VAqMf8oZVPOuTu7WawAOCgVUKPK3WsKUaqVBUaH3DLUj0fuEql/r/heo+Men4t9v/o++As0Yzqgl2OtNWJ6Q7kMnzXkJitZUDlpxqi/iSgKsLIAECNAaSvxvhWAqZkuDr129vnFSjXRpAN8Ssi2TqIAVWhNbm0lEnlangAQlNyMSrUKpJShIfGnVZkMaqMLQYxieUTYhImnTJk0930Ema41BxOPjJMONBoENsq4k3FMmGmV9xc2anHcdZeHKa19HNBVoodlIacAGm/7Kw1VdB2n2mM0am0GBOPpkx8legqwc1XLM9AImq4ONbwID/JlMrmKdQ7aCpnbQGuhkg/O8uJHSDrfBzotzLt+H10tJ0NRCxCLQZqNXvkMWGTacVDZGvdxzmfjJEiSTXpPk8fVKcqfCzNlsMfgY5JyctHmqq4WbGRW0HCBLRIAH3ot6OJlVIYqKCYpVr2Uw6FLbWloASeC2KnBEfaJ9LjesvJNsYLIxrgczkxVEsIKMVQIL3LjGxkYLUMFis6KiDHt37ULJjYIGoIKJJAQlGjdvJuHUoWEhGmhllOwHni+bG7SnqHEqRYyyhiIzWQFcKtNDIev8N5mW3BRyLDMHgdeP58qGGoO5yUY2+1qEiWqgTYVYq9Wjrroc508dRllBHsy8bk7Kf5UKgWCDbuPEz7H4+aG2vk7YldyIqwwCtzQoBayw2oRhWOWoEi9w9UwqQM1kVgoCYaSDAJwC9XjMLClUEBaEYcN7Vl5ajuv5ubh85TLCwsPQ6bbODaz82tqbQIXLUyf3XhiZDK1ntoMcqxUhEU2Q0LhpQ8FzExBzwV1Zj+vlxfCx+8Ls4wUfpxO+Lhey01NRWZANg1iNeCEkIhZJ7TrCY7HB1+4v49HJoFoPxzCzCgicOEVNsGPrBjjKixAZES7hu2xSs0gjUFFcXIwaGef1Ml4Y8norQGvy9RZFk8nPT2w3mFNB1UZJSQmW/PgjEhMTMXzESMQ2ikdBUakoTFRjRYGovO/c+PBz+DftUEpKilBWUSKsVzbMmJVy5OBhvPLSywgODkJtbQUKsy9j/47NoqioKKsSIKYetahxkjHhLVJsT309WqakoKSoCKUlJWJ3FB0ZgdrKSsTFxCIhPl7mzIIbhbKRTb+agfoaJ4L8AmDzMcPoNsDoxWBuglkBCImMlPDrlh1bwy/AjOr6ClQ6yqTxU1TswNoN28WKhpYNkXGhcFSXIipYARXxjRPRuf+dCIprBrPVXyzZiqio8AYyczJx6cxZ9OneQ9RfOQX58DW6cT0/D2GhYbh65RqaJDRGeHikNDfrvSBNcDZr8/Py0Tw5BW++8RY2btgoXubyRysIvTnva3MSaA3o8cBuNaFjSlO0jItHclycqD/qvN2orqmDx82moUmYfAQ5CQoW3bgh+TEhARa0a5OM2JgmqKv3RTkZvl5O1FU54HQ44SA73GqXRqq/1QojrXBqOTd5UFpbj0Onz+GT2XORV1gEl0EB4sypCIkIgd3ii37duuPt116HOSQYjAKXovwfqgTOo9V1tcjLIVBxBW3aJiMmOuwWoEJZDP5XmpAqSNXS6IUzZ87h+PHj6Na1B35e+QvWr1sv41YHKnTbNQVMMpTYKLZm3IzZjEDLRpHolNIIdhMVZf7wM1lg9jbCR5pEasMSGh6qlGwGH5jNSp3DZz0wMAj+/gFyvU3+NvhYvUFUoLa0HGmXr4g9VFREHAy+JrgsPvCLjMa8ZauwdOUK8W4eM+5etG3TBkFBDAk2SKN2w6a1kovSrHkLuD1mtEhpIcx4IR5oikGZg10GAayvXy+Bw8HmmxFZ+ekor8xHclISTp48iqZNmwhTu6YWqK7ywOPyQZWzTKzb/CwhMMIbtY5cXDizHSGBTnTt3hPOOj8YLRHIv14jwIbLVYvy8jzkZ5/APXcNgLelEa5lO8QCwUwloseArz79DBdOHYSzxiEWQ7KhMShmmNnPihvM2fFyISEiEB2SE5AQHY5Aqw2uOmapeKPw+g3k5eSipLQUIUEhMtczPN7owzBoHwT4BSuLsUA7WndoAXuoFdm5GXC6axEWFiKZUS6XN1au34mFqzeirJ7PDwkcbjSNj4XX/2HvvaPjqs7u4T29qfdiyV3uBTeMKaZ3DIQSmgkhBAihQ0INhJgWEgih914DhG56s8EY9967JVmS1UfSzGg0mm/tfe6RDW/ytf/e32JYXrhoZu4995Tnefaz944nEehNY0xVOfafOhpIdCHp86JixESES0ahI5kJXyATocygzu2uaAcyQhGnuQHqfI33sIDvU7wl8F7Epl60tLQZj4pwAOwm4P7P4i5lnwhUsEO+rqHOGELn5MiLgp3yxmuAZtpeEydIJtmHlrZOtDST5RWRtOAbzz+IHTvWIRaLap6FAhkyP4eLDQxAgEV8rwt52VnIyoggFAho7TKeY5GWjQ0tlP0iq2X4MJxwyqnIzuuPHm8YXb0uJGJefP7el/jg3beQ8kYRS3bA4wkaE2yXOdMJWHD9JLsT6E0n4KXJb3sH6KmluJPz0kOgxXYwMsYwTQBGMtUtGcS9XzYZ5lruTRvTyXh3UrKOBNLCEXOuuz00H/eLTSGwQg0RCRQU5GG/ffdFRUWlgIqa6mp9PDuFGWcwuWWnp6ROtU8Z7wwBFmwgcqSfGEPYRgN6GglYcYAK3kJjUwO6u7knkuXB+NJIe/LMURzuyFzJx+onQEUwEtzDqKDBJ81Qud/2MSocmVKykSPGiJpARSIW7wMqGJgQpLcAC7vJKV9FA/oMglEEgj1etG2sU1zH/Zad4tZzTU0VASPxxK5jXqeRUzA5C+NJycopzjPNG8wxBg8bgDPPO1H6//+48ymHcefG0TMOkW/CnC9+wPYt1fKMaGpswWP/eKkvzh9c1V9MBc6/vYGKN1/6ALGuBE4/17znn3c/be7L5RaQce5vT1Hc+tdbH8Hvrj5X4MCrz70jCSnOwxtmXap9kF4Tlnlt9miPGBob1m3RHOC65H3tN30iDjx4XxkuE1j59+sf9TWO8dkNGTYAMy/4hdhR9Hvo0wB3GPP0AajdWS/pKgtU0NRbhSunoYzzl4yKQ48+QH4bb73yYd80pyxWCZkYT72pveuXM2eow//+u57o8y68+Y7L9fN33PwQDjpsKmaccrgYBt98vgCL5q/A5P3G4pczj8eSBavwwlP/1nPi2mTszzGbuv94TJs+UT4Dzz3+pjwmhGeTCUUz5OmTcdpZxwmoeOnpf2tNVo0YhF+TURGLG4DE8Ve86Y7LtE8999hrAjgmTB6DZx9+AS89/iLysnPAtrCLr78E0487BC8++Ro++2QO/vHEnWLrHX7ob3D3367GSScdhscefkXeFzqjpQLgVm739Zc/qNCt/KY3jYmTRuI3vz0Vxx43HatXb8QNf/wnjjn2EJx3/vHYVbsb9979lD6DJtdnnUuPip24584nccjhU3H6mcdiV00DPvpwDuZ9uwTTD56MmeefjAXzl+PJR143z0AJm2F1HHnsgWJY0LPh9lseUd7OHFPMbHqE3Hu15tY7b37W53/FwIWxPSXF1q/dqq7vm2+7BKNGD9H+Nn/ecgEDzMOvue587DNxJJ57+m18+fn3hpEGo3PPZzFm9DBccfW5aNzdgtnvzzGNd5IwNn5x27fXSuvfMioee/h1J+ZL4bY7LpM3xYP3vyj2imVK3HLjA3rG9L047fSjVMD/x33P63nS6+Oqq2fKv+Hmmx7E/vuPkzn13DlL8Ld7ntHwEMT54x/P1zM579wbdU/qcHdqB1bGRvl/TxLHHD0dJ/3icHkhsEv+oQdfw733XSOPCho484uvuHIm1q3dgj/+4T6tQ+4xTzx9m76PptmcvwQqyKggUPHxR98pnlORV7I1aVxw4ak4/fSjZOj8z/tf7MvPzj3vBMw8d4a667/7bjmuu+58bN1Wjcsv/6tZ9/SJdKSby8oLcO/f/6Dnd955N6uxwKpGqAGhtxeTJo3An279Hdrbo3jtxffw2vNvomrYQDzw1J3YVV2Pf9z2EC644lzse9BkfPL251i7dhPaOmOSaky7vOjo7NJY33HnZTKxvvKqvxkAmzUlx1OUY0pZooOnT8JXXy3Eq699orn+p5svFJPhb399Du+99zWOOmY/3HzzRZJ++vOfH9E+TBNrAhKUunry8bf65J95rwcdNBF/vpWMip244AIDVFj5IO4P3FMvvvhUnHfeifLvIEuDa3HKlNG6HgIVF100C7fccpH8NCg3RYkoYvcTJ47APfdcCZpez5hxBW677XeYMWM6nnnmXSxcuBp33nkpGhtbceqp15r560rjUgIV5xyHF1/6EI8+8gYef/wmjBlTJcCBEk4n/+IwB3D4Fjff/JDWGr/jsMOm4NNP5+OFF97HqtWbcPusS3H00dMw6/YnNcdOOmkvoOLPj2lc3n3nPoH4Tzz5b+3FMoJ25Nbr6poxb97SvvjDGmDbPceaVev8k9eDYTNw3vR5nyYM49HsIaYeaNnMqhPIx9U0B9u1IhkkDp5T+bdAhSFCc74YYMLMC6cBlA0gToYjQMWpqTFy4vm0N1Ax+vAW7RlskjAqFcYsXA27jq/uT5k79iDi+ShpcXt9alKmxOYe2aifxmaEI2wDtf0329xgGjpMc7IFYqzsk2l4YHxhm73/M1BhP9OpMGpcrBcoa3DyELHj4dTsDIBkvld7k/MMzRgYFtPPjIofhdk//+H/hBEYSvqXE9jyfrjZWzaFBR0s3Uqaac7CMTJNaRXzLeXLyAMZPXq+LP19b1qT/QxusuxaYmG9j+7r0JyszNTe3gxWhomfZbS293Tjk4ZOQMAWDAWAqOvTFPjJkBCtjrRgmQIblN8gxyao16ZCzwpH8opJDjcybsRkAbCzWV2DNCkURc8mNpY+bzZ1u5HxnuKxmMaHY0U5AGor8hpUsHXknPgeyWnE432FUwsCcWO1VDsrI7W3mQ+zYoO2Mkk2zApu4sZnwgBC/D3vmcVkahTzXlj8ZiGbxVQ+T+OxYGjyvBbSoSVp5aO2N+l1BjjiQcYXmS3UMub4GBogO1YNIOH2GoNwGq1KDslhVaTSvJ6kpKGOOesch1HBDdc8RwP4JPpYHTL0hgOQpChtZcylY10xXS8DESbNnHssOvPvWLSKRCIoKytR92ZXVyc6OqL44ds5aKqrk5m2pJ+YTMONqhEjkfZAXWs0O2bxjWANk20WK9mlbpkdvF9zKBspJwFYzMs5frG4U4g0TJbc/Dx0OSbLBHO0ZlTQaTUG2NQhdaXhd6XQVr8TKxbOQzrRRZ0JFVn4PDmf+ZzsmpQ2ND/LQ9aHATAIMHFO8vMJjoQzspGRmdEHypk1aIolBMhEuXQ6x2wQYoIWYwTOF5+n/UX2yqaNGxDv6sCkSZNRXsGOG/pGGP8Pdeb5CFKZ97ArzQJavL7MrAKMHDkWkUgOkgYXUWCgIonWVQ9a21q1Pggq0ACRQEnNxlXSU4/1dOPQw49GRl6+OrLZRpuSNB2fg3QydO+pnjQ6OzuwctVyrFi+EEV52RhQXoriogLp3HQmkmgjq0U/F0U47Edefq6KGZQRMWsqpaIQx4mxTHNLK5qaW5XsP/Pc8xg2bASOPvY4lFf0R3NbuyRqzM+yWz2hGwuHM7BzZ41kl8jkqN9di0SiQx4VLELO/+47VO/YiT/+4Y+oqKyA25tC/Y5N+Pjtf2H9iqXojLYjyfsiW6aXz4Tj4hMLYPjQKpldVm+vRlFxASr6lSlpzs2OoGrwAElldHS0o5MMnrZO1Fc3AF09qCgsR2FGPkLeAMIeH7LYzRbyomhIBQorafacQmNTPaLxKOJIY9n6rXjvg09BWHBoRQXS7gSSqTj6FechKyuIwuJS7Df9WBRUjIAnNw89bqg4wudeV7cLNTu3Y8rkiQgF/Zg7dy6KCvOQEQ5h7Nhx2LFjhwpow4cPd6T4ehHt7MI3c7/Xsx0yeAiuuPQyLF20UMVQWzSy54OlFwskpDdNJITxVYPFqqDmfmleNkqKChDJyYWfgGOaiR8EpjQ0NmBn9TakU93Iz4tg8KDB6N9/ONyeHMQJgrt7gGQcSa5lsoEF7gURjITlQxHr6kSsO47WeBfmL1+HO/7+KBrbojI/d3vSYhCVlvVDbiSIKWOH4cabb0BOaTl6vSF5Tvw3RjL9XWpqatUNPXLUMBQU5DthhZFoM1m+lSqx/zdyhGSW0AGDza38nJ07duL551/CBx+8J/k2FhO5P3KPMEA5i0uQDArnOAvRrmQcYwZVYNr4YcgKuRHy+VGSX4jsjCyxS6prdqlI2tTWipbGqNhmKfrUJCkbkELYH0ZlRQX6VfSTrUZeUQ6y8zKRRg/q62uwa+cO5GZmIZCRBU9uMWo7unHxVVcjnoxj+vR9cdQRh6qTjKBw/0ED0N3Ti+zcAqxYvgr5hYUoLilFcXEZsrPyEAxEZH5r6OYM0l0sg6C6ugZbtu1ARlYmdjc1or6hDv0rBmHHzu163lMmT0Ys0Yu2aA/aogkkumOSpImQeRTIQLyjCevXfAWka3HoofvD6y1CLFmE5tYgmto6kUYb2tu3oL1hDY4/8mCkPQXoTATgDdK8OoH2pjbccdvt2LFlnSMZGDVMCjUu9EiWqKmpxZyxQS+qBvXD6MH9UZabgTA78NVJ5kZzU4ekL1pb2+Ql4kIvwh4PykpKUV5Wifz8Agwc2h/FpQXaO5pa6pHo7lIhu6vbha21LfjnMy9ifU2DTNy5nwa9bgwZ0A+prigyQx6MHVGFKZPGobOtHt3JFIaPnoKcivFoSUXgCWchIyusPb6luVlNDDxzOXdMUYvJU0ASAWzWYHMI932CK/w7GtfbLrmmxiZ5RxUVFUn6qWZXrWIOxk8CABgHSYeYnd3sxksYCcHetGTAWpqjyM0tRFvjbnz69kvYsmk10ukYenri8rHiHOBZGfSk5EtFYIKeGoxhwqGgTJiRSEmGq7Ujiq6eJFFRHHHiKWLo8RwlsJPqCSPe6cHLL72Med9/DZeHvlox3SvjD8aPHhipAtOskkCiN45ErEv69kpKHSkAJYmOV4M66WzC7nT5KV21WsVOHG1jbSk+ygA4hWAkA/5gCJFIltae6YE1wAe/z8oa8kAdPHggJk3aR+cUzxh6wXG/pBE1ZVx60j1qbhB7V7JSbvgIqijuNR4cbIThryTBmL3iA8WtvW60NDVoLyFLhRKDlAlhrMZ7tWacivWd4j9ZpNU7q38k/USmjmRm+D2SIIlpn1MBxETk8Iqt4UJ7WxSJrpgYMVZWNdrWJqCGc5MgRSDoE3BigJwAfIEA6lbtQIjNA+oKJQPFb0ZO52mPafZxHotJ8k3BW3E2fUHU0MOYmddk5EquuOE3kiyiT8SqZeu1h8447Ujsd8BEfPHxt5g3ZzEuuuJsFeHffOVDrFhCjwrg8GMOkFk2WQ4vPP4mLrjsTFQOKJfnw5oVG3DxlTORnZuJ1194T74WXAs05T7yuIOwYe1WPPHgy5J+KikrxItPvYW1KzdKrpIyU+x8JnuAbAe+AkG/TJKpF8/POODgyfh+7hK8/9anKphQ+ojeEPSteOS+F0zO4MSlLIZcdu2vZF79ynPvYc3K9Rq/8opSFBbnyXyaOcxFl58lj4OXn34by5euMXmAxs6M18QpY3HK2ceirqYBTzz4CqLtHdobbpx1OfLzc/D8U2/q5845/xQ0NjTh77c/rnh04CAjwcR9ktJPZ/36JEyZNg6fzf4WH737jWLGg4/YF8f94lAsnr8SH777FS6+4izFbE8/8roK9Yz9b7jt9+g/sFyAyLJFa/pAFMapBCpOP/t4LP5hhRgZnONDhw3Eby75pYCk22962JFQSuDmOy4Tu+SV599DeXmBPCoWfLsIt175Z2Swgcjjwt+evw8FxQW49/YHsWnLDvz9oVkqnh9y8Pm44spzcNnlZ+PTj+bi0otvNax4l0cm0jTUpa/K7XdciZqaepw380YxAjkvv/z6eUm5UKu+vKIc5513POrrGnEP5cSQxgEHThJQQeknSiKxME+WxfvvfIkP3/1ajVo05T71jGPkj7Fw/grM/PXJaNzdjLtnme50xgH3PnijmpmefPR1LFqwQuxtNey43bj2+vMxbMRA/OuVj/Dxh3P0vQSLJ04eLS8M+nAcO2M6zjrnBKxetVHrr19lCV596QN89OFcnHH2sZhx0qEy937i0ddVQBxcVYmrrj4Pbe0duOO2xzDrriuQm5OFxx/5F5YsWqPrrhhQKm+ur79ZiCOPmCaggt939x1PKtesrCzFdTf9FsGAH/fe86w+99rrzkdNdQOuuepunTtHH3sAzjv/ZCxcsBJ33fGk9t6pU8dI6mnr1mrcevPDOOCgCbj0srPw7dwl+OvdT2oeTJs2AVdedY6K+PSoYB7L/ZMySxyzC357Kk6YcQg+mj0HTz/9pmFUHToVl112Ftat24qrr7wH9953rUCUvYGKtWs248br/6l9jp/zwkt3a838auaNmruUfiKj4qEHX6J4LGcAACAASURBVMWHBG3EzDWKCdyHaLJ8+ZVny5z62qvu6WMv3vO3qzFh0igxS157bTaefmaW5s2ttzyMpcvWqsHxst+ficMOn4qnn34LBx88BcOGDcCDD7yCjz+aq73uzLOOw8yZ9G2Yo7347HNnYPZ7X+Hq3/8J3bE4TjjxcPzl3huwed0W3HbtnTj5zBMw86KzMO+r+fjjZbdKjre1M4GjjzsUdfXNWL9+K2Z//Liu489/fgxLlqyRZ9MfrvmV7uOZZ9/BKb843Pn3R7FwwSrtQWQl0NiaHhUfz/4WRx+zP667/nx88cUPuh/uwQQRyKh49pl3jJm2VcxwQUD188/N0ny+7vr7sWrlJs2NP/7hPAEP9Grg/nTlledgzpzF+MO192le0L/j5pt/K2Dlogtn4ZZbL8axxx6Af/zjJfzrX58qzz/nnONkcr1y5UbJZs2adYkAk6eeehsPPvgq3nzz7ygpycfttz+NTz/9TmfsLTdfiNNOPVL3y5955unbZBBORsVHH32P444/ADfd9BuBEvSo4Nn/7rv3K/698cYH5HnC5//AA9dh//3HCzh5552vcNJJh+KWWy7Ep5/Nx403PaR59OjDN2DixJG4994X8Nq/PlV9gXKXhxw8Ed/MWaoY0jIFVKtwAEvLlOD/TQOyI7fuSDgZhQtTx2INiPPDNBp7VCcUi1uSz91973USFhOXO+CUOXdN3mPbrVTTIRhHGU3nH8TmcOqG/EEj185aiynCr/uqyH48CFTY2pitASr+ciTU9Xd7G1f3vXOPOTbrb9zruA70UuPtjztIjAcigRITL9maif04nqmMVS2rQv9OKSYqmLAh2lGP6aPP/uTz+8Zrr/hQw+Gcy5x/ap4QY8QwPi0IZWtwrM2ZGg4ZuKzhGll2xWE/e1Ts9eR//u3/ESMwhEG5NW5hkuNQjEyRc2/vCqfUIsoUpVmIjhpjY3VUO34U9j3OHtDncaCus71oWUZSwBjhiFXRR7UyxV+7dVhGhjZbbR4Gp1URXRuTQe4NqGDZG0xATWeCFrHDCrG0LCMDtYddoI1SHUima0zUSBlWm4XPw5/Grvw7JtqWHcHPYCchNygVX2XEZeQeuAMyAOVtGZDAdASryOag0xwz67nBz2bgv0fWylDD+LP8HiOv0yOpJh0yNJ1Wx7G5RyNH5VXXB7/bdnLowHGeo7Zft3kvCw28FhZ+eBjZZ6PNzuNxroVotXlG7H5U550YFIbez88zElrmUEq7elWw4COi/j2ZEfxFcERyUEyY0ykcdeZZ5qBzwCYLjnH8NV5OsZwFAIFPewEV9KKwQAWL+fw9uzb5eew25/MrKy+VeSKLnW1tLVg4fx6adv13oILmbkygfR7KLYWQ6EmhjcWNeJy8RQcd5+063ZFeMoHYCWAAL7FDnEOa84NdfpSh6iYqvpeXC58/izqhSASBUAABdwo71q/ClrUr0NsdQy5lVkIhyZtYkIL3ZZlKPLjcXgNgcM7x3/iy4F8kKxvZOTkOWMh5acA0zhd2WVrmlA5E57rMv+/RfeTYS/sxlVIHWG31duzYtg2DBg3C8JGjZNzNzgizZllNN+ZV7IAUOJg07AIWCbKy8zBk8AgUFZXJFJuDpfnkmNMLZEhRB77DXGMwqH2lu70JC7//DhnZOThg+nQEM7IELrE8pY4ZyiTozs1eQLkpfs6O6m1YuOBbpBJdKC8ukAG1N+BDj8uL3U3NcCVodNsmbwN2o8qMHATjKKFmfF7oUcIJTKCivmG3CihPP/Ucho0YgeNnkFExALX1Dbo3M6bUQ2ZnLzXEg9i+vVrSUs1NLZLMiMVo5B1Dy+4mSQstXrQIf7r5T9KiT/V2o3b7Bnz45qtYu2wROqNRGXV3q8vNJ+PGYMBDmosYFcl4D1YsW6WiQv8BFcjPZjE5jcqyEvSmuiULxWIPOzbTSaCzuQNI9CIzkIGscCayMzJ032WD+yO/ogTusAexJBkRjWhpa0F1QyO+/mExFixegX75JRg+aCBi8Tb0pOOoKClAIOgSQDN+0nRklQxBZkkZulzd2LB2iwq0jbsb0N7WiiOPOEyslmXLluoa8/Pz1Em9ceNGFdmqqqqUwNXV1cEXCGFXfTPaol3ym7n0d5dgzcrl6E5QPmePSathypk5Ly8egjSRMMYPHYyxVQNQmZ+LkuwsFBfmIiM3FxmZOZJvIbbKYsCu+lpU1+xAwJNGaWku+vfvj6KC/vD4ciWDlPalZJJLrSayX3zeAMjiYDGaRsLcSxI93WiJdeKbhSsx656HEI0nqVsGl7sHEUqdFZWhODcTowf3w/U3/gGlQ4ah18M59t+BCoJsO6t3YufOnRgxwgIVFqTYi02RNp3HNsLnPsp+RbeLBVeXZFtWrFiFl19+BV9/8xW6uqIaKytDps4jyRC54Q95BYixsJvq6sDgknwcNHkMSnIzkB0JIDczG8X5BQj4aKDdKOmA2ro6bNlUjURXQvrvNESOBDKokaRjhUydQCQAeNPIzMnAkKEDBIo17q5DRjAEXzgL3rxS/O2J5/Dm7A+RnZOBww89AKNHD9c+OqB/JdLuXvSrrER5v0FYtmyVwJQjjjpCXfYNdc2SSKLfC9cdi5WuXpekt6IdnViweDHaO6Jim3Gfy80pRKongXVrVuKAA/ZHojuN1vYEWtpiSPIcjwSREea6yEKsvRnr181Fe+t6HHH4/sjOG4D2rmy0tIXQ3NoJpNvR1rYBXS2bMOOYw5F2FWDt5np4AtTdB3riKfztzjtRu2OzwHE2KFhvLe5LPLNbdrfIOJ5bVj5le4ZUYGT/MuRmBJAZ9CMYCCPW0SMpCXPm8VcSYZ8fBfkFqKjsj/LyCkSy2NXO7vwEOmMtiCdi6IqnUdPQjrc/+hqffr8EsTS5enwuKYR9HgzpXy7mXlFOBkZUDcKoEUORiLXpOkeN2Rf5AyegpTcCT5BrNVePtLmpSawOezbrXGB85fap4CUZHa9PUpFtbW2SFmPByKh9uiQ9RqCCTQQy066p0blFoJJNB4x9CITwDKFsJ1ws0vPsSaMzGkdLSxQ5uQVoqK3Bwi/fw5pViwVUuEBAvFfgAQH9UJBm9vSZCiIks1sjMcTVIh8J+md0x9HV24uqcRNwzCmnI5RXpGaEdI8BKtqbe/Hss89i6bIf4PaSDUNPrIQaXPgdBD3EYu1NoyvWgfauVrECxAh1vsuyQm2cqyR9L48KdRfvpYdsG3762MTqRqSnRK+YBfQl8QXCakAxQMWP43Gy33htPMumTJqAktJSNNTVKQ7hi7Jd8lRjTMYYTVk1y5Iu3Y+HcTcBiv8CVPCsNkAF0NK0W0wEAhUeH2M/Y/xqgQp7z6bIYBi5/3+ACrJbOY7s7k10xgQ+2Y7GaFurI31l5KtYpDLm3gF4aTju82PXyu0CKlhM5HPRXsAYUh5fjE8d5RBH+pTnvmHbMV42/2byDFPUZbx11IyDcfAR+6G5qVWMg34VJRgzYYTi8s8+nIPPZs81AMPxBwlg+X7OYhVX958+SfstAQ4CERdfMROVA8v15x++W4IjjzsYR+k9Hfjum4VaG/sfPFkxFE2t+Z5LrqH0U4Fkk7ZurtaTnbTfWJxwyhH6bAIVfP+EyaNRXlmCzz6ci/q63fjlzBN0H999vVA+ODST7ldZiq8++x7vv/W5yVudo4VF02NOOBiHHb2/DI8pr8S1Pu2gSQ74MhsL5i3V9Y8cOxTfz1mCdWs2YfEPK7Vu6VfEfI25wdU3XiimwvrVm7Fs8WqMnTASI0YPQbStQwDCjm21uOK638jrYuG8Zaitqcd+B06URBWZG7NueABHnzBdfhRkeCyYt0LSd6PHVgmM/O7rRXj1+fdwwe/PwNgJw7Fp/XZdB8Gc/Q6coLF4+N4X0NDQuKfblUbf+0/AGefOwKIfVuC1F95XDjN63HCc/esTFePecfPDjuSZC3+68zKtm+eeeAPV22pw5Q2/FTD87VfzsHz+ckw/6gCMnTQOcz//FrdedzfKBlbivkdmSfrp0IPPR//KEjzx1G0YWjUAn3w0F59/+p3YEMccN10AwqW/+wtefv1ejBs/XMXvL7+YLyYEGRVLFq/CDRyDow/GBb89SfP94w+/EQOFYM85550kRsVf73gCx804GCedcgRamtvw/XfLUFJSgLHjh4kNQumnV1/8ANdc/xsMGtQPixetxvIlazWOk/Ydg00btuOuv9BY2EjH2k7pgw/bF2efN0Nz6/OP5+kZ7HfAPhgwsBz/fuNTLFm0GtfecIHkdZ9+4i3lmDTbJkPigfte1JS68ppzUVScL48JGm4fevi+6D+gHO+9+wVefelDnH7GsfjFqea6aSrMZ3HIYVMkX/XUk29oXf32wtM01+d9t1QSSocePlWG4/TZuPee5zBgUBmuv+lCdZTT12L9um1ijt1004Uqhr///tdqpDvsiKmS1lm6dK3MtI86+gBccumZ+OrLH/DPf76keT5p8miHURHH+b++yeQuVCVwgN2p+43DlVfO1J5Dw2d20VOyq6pqAN5841M8/tgbfUDFA/e/qPPv8itmYu2aLbj26ntMXu0Cnn72dt3TeefepDG//IqzccKJBws0+X7eclD2inkYzxl7ltxx12XYd+o4LF+2Dl98Ph+Tp4zB/gfsA4Ig1193vxoNCeqcdtqRAjTef+9LlPcrwQknHIy6ukbceuuDmLDPSFx40elob+/A++9+KVm0k042+8df73oC2TR1v+bXqmO886/ZiquOP/lIycvN/3Yhrv7NtSgtK8I9j/0V/QdV4vOPvsIXn36LKQdMxjHHHYLv5y3DuWf/AdddfwEuvtQAK2++8RkGD6nA8cdP17q+/vr7cdVV52K/aWOxaNEaARW8jzFjhup777zzKXzy0Xc44qj9cP3156OpqQ2vvfYRlixaK1NrARXPvoPHH3tTeznPUVuvuPTSM3HuzOOxbVst3nrrc4FaZCDU6nuNj8Nf775ScmOvvfaxjOT572VlhViwYBUuuuh2gRannHIYamoa8O47X+m8PeOMo3TG3H//S3jllY/FqKD0E8GPhx9+HZdccjrOP/8k7NrViNde/0hgEEE2+kg99fTbeOThf+HJJ2+R1wSBitmz5+HII/fFn265UPf38suzsWDhalx7zUwceOA+WLBgNebNWyYJqPHjhyufmjXrCbz3/hwcfdQ03HrrRZp7L70yG4sWrMHYcUNx3R/PU9776qsfY3djK4479gBJkD3++Ft47PE3+uqTOqfZkMiCNwEx5tJ7eYbwMyxYYFhoezxkbWGc8Z5hPzEmMg3JBqRmo7FbzDQjrW7YSDYOtHU7W7Myza8G/JBHQ49RPdlbZl2sCsmXA6v28qgYeWiTU88wcQvvhWePJCUddsV/AypMncQU9k1937BItP39J6DC8c9gLcZILlEBw1wz/+P1Mt6x8Qnvh3OT92/rfBwPEz//2J/FPhgLgNj63B5lGQIp9Ik1sYkFKuy1C/BxG0CJXjnyK5S6jCOH9TNQ8X9Ebf7nm9hrBAY7pruGFraHMWEPS6uvS3DCgg9CG52FyQDbop9287NdUqIAClhwvCecJMomNhaksN3ddlOzXXw2OeOftTE4/+fPE3SIOVr82nQEFJguRl27o6Fq8nVzHdwk98g9uZwCv9lE+lgdzqatTnMre6XN3XSes2DP+zUAhdkgbdJpvSr4XQyiRDVPdOv3JvExKKhNYAUmONcrWlpfGcokTFZuS1ujA+xw42Ti38fIUDc4/SliRvOVtDDqLieT6mAUG8Lp3mOuTdYDAzRKLxD8sIVsARCOh4fdWNXcTekDq31nDYlI+Qf/3qF/OwcgwQl+f7cDUjDTZ/eqAAqwEEE6YQpH/PIMx9jVkfNwdA3Z+SyQJZ02nShOh9uPgYouB6gICEBiAZEFEcp1kQHAjiVK+3DaxeNdkkRYsXQJmhvq/yujgmZ/BKKon8wgsptFehbeXdRz9ysJNoeT4/8heQMaH5uyofw2aDLKa8nLE8jD9/MZ7JkbBjhj8TBAzWYWoJMxbFi5BC11OxHye0QtNybiZr5yzltAR/NaEgY0kAw7VGDKhZn5KDaQL4BIBsGOYJ8HiOnYNLrVPPj2ZktpPVuGlNOJwCKD1qsD1DU21GPzhvWap+MnTER+QaFo7KaLIK1CoXxL2HHLYig7ggSa0eQ7jLLSSgwaNMzoSPPQdforKFXC94iuS9AtSSCL2uc+eNGD5UsWydC4/6DB6GWwQCBIlQajJWzW64+BCsosLV+5GNs3rkN+VgYGVvRDdm4O3IEQmlva0ROLiXXA6ioTo6ysHHg93L94VUbvnCATnzeBiu07dqrYwS51enQce/wJqKgcgPqmZmTn5GtMuJ5okkqtfhavZFaXkSXpnfqGWtTX1Wju5GRly0x75fLluO4Pf8TQqqECbKo3r8P7b7yEdSuWoqujE72kU5Oi7fcgIyOIUNCLZDyGMSNHwuf2Y/73i5FIJlBSUoQB/Svgd6dRkJsNH4G5eAxZWRkI+PxIJ3vhdfn0f74v6AsgOzsLRaXFyCsuRCArDFfAi65EDE3NzaiprcPiFavx2dz5aIt2YFjlQFRVVqCprR5uH1CSlw2fL43svDxM3vcwVA6bgNx+lWhJRBGL9eiZV+/cge3btuKwQw4RSLtmzSoE2J2WiKOiogK7du0SUDF06FCtbz7vgqISrFqzHvW7W5UgXnn55ajevlXduHavtHuznesCqNNATjgoRsWogf1QnpeNYgIV+fTVKNTzCfgjSCR70dzchE1bN8kUNi87hEEDy1FeWoKszBKEIoXqPo8njVQX5XbCwbAKXuxq9gb8kqMjGCkT6a4OfPrtQtx132OIJckoIn6ZRDiUgYLCYvQrzMOQ8gJc+4crMWSfSUjC/1/NtLn+kkmajW9GfX0dRowYjsLCAlNFEpvi/xmoEMMhZbqQv/jiK7z11r+xctUKARXcl+wewn1EFG2/B8GwH/FkCtkZ2ejuiqIo4sf0yePQvyQP+VkB5GVloSg3X3OmcXejiqec64kY5bNa0N4aBTfHcCCCLLK4QhEZkIri43UhGmvT/C0vK0GQ/h6UC3L70BgHLrj2RtTsbkBxSR5OnnE0DjhgmoDKjk6yiZI4/PAj4Pb6Ub2zDrvq6nDk0UchP69IgGJbe5c6/blX5OXlaFwJzLV1dGL7zmpsr64WOMx9ety4fRDrjGLH9s0oLipEdn4RWltjaIvGEYt3I5IZ1lrPDmUjFm3D5o0/oKZ6KQ48aBLKKoahqzsbbe0BNDVH4UIUzU2bEGvbiuOPPhReXwnWb2mUhJ/A+q4k7v7LX7C7bjM6uzrUmKBuNYf9SfC5taVD3e3cA31uoLwgE2OHVGJIRRlywz4U5BUAvQRfDBNC0l7pXj2jQknVFcs3xRcgoy2J7p4Y2jta0NLWitr6ZixetQGfz1mAzfVt6HF70SOqKBkvHgyuKBVQUVlWiBFDBqKivASdXa0q5I8ZNwVFgyci6sqGO5QtIJNyejw3BcQ6QLfdnymtwz3OsCEorRQT+M75RTajiT/oCdOMvJxcFBQW6vnW1NYITMiUTKE5n3hus9GB4AIZht3xJFJJ+gN0o60tKrPtHVs2YtOKuVizcgna2xpphQM3eiW9xKSQEmH8XhrhStbCYQXQQ4L7YVesk+QfhLJzMOP0MzFk7D7ocdEQ2oPeHi96kxE07OrCY489jq3b1wPuGFKpmNl/eHbyLHO+qyeRlOdQEpTAcpixDiPXFLvNmWjjWHu+agxNimwSXafpxiampnDMc5OshjTCPMPDPK+Duk75XziNPkpcHdYDmzIYl1ZWlsvnhWAC9y811Ii9QqAijSTZR0zInQ7HAGWkWMDXmftfGBVOU5Cv14VmSj8RqMg2jAp6RLH5hN2GLHrYOF/ND5JZTf1noMLtNeBIskf7qRqJxKjQqGk9sejBbvx4Z5cYO2rUcbvR0c4OUTb/MObuVUGW3d6cS14/AR0PGtfVqmhB8IJ7g/X6UkGCvivdiT4dc9MNafS0Vexgl6SY2vyOgIlVHYb0SacfiUlTxyEUDonRu5MSNQP7Yc4X8/Hph3M1jjSSPuTI/eR3xvtqbGjGFx99i4Xzl2teUMZJQMUrLPwv0z0ccuT+AjnksyB5qxZ8+v43kijii3JLMtN+9h2ZdnNdcd3tM3k0jjp+OgqK8jQmHdFO/DBvKT789xd634QpYwWC2H8nQ3rpolV4+/VPHAaumU+m4crkPoc6109mCF8EZr7+9HvM+fIHPd8p08ZjxilHICsnUybdD9/3nGJ1Mjl9zImSPRqTX547AwMG9dO+Qfk3Ftx4fy888SbWrt4k0OTYEw9FYXG+EzMYSTi+f9aND6g4ePIZx2DivqOVa/HaV6/ciNHjqrBz2y78/fYnBFDRV2OfyaP0M7y+2uoGfPjOl1izYpORn2U87HTa0svi7PNOFqPiuSfeVL40ZvwwnH3+SWJU3PmnR/uav2656zIEQ0E8/+QbGvOqoQNx4OGTMX7iGDG4411xzP96Ph6+53Fs3l6NEeNH495H/yJGxRGH/VZ7/9CqCtx++xWYMnWcuYdYAvO+W4I7Zz2mwjuLuLfdfgVYBOe/M0dkMfrmm+6Vz9CIkcNx2umH4aDpE/WcZn/wjcby7F9R+qlaQAUZ4zPPOxn7Th0rRg29Nlau2ICx44fLA4QsitKyQr1n2IhBylUZ2xM8eP2lD6Wvz32ZzTqK3VMGtNv/oIk4+bQjZIDOtUDwZw69QZ57F7+/8hyBLp99Mg9PP/mmmpNuvPV3mDJlDD77dB4ee+Q1jB4zFL/69ckYNNjMAe7jc75ZhGeeflNgINcWu91p/E0PEr7INPnw/W/w5puf4NDD9sXvLjkTmzbuQEVFMXJys7RHLVuyFo8+8poM1LlWLrrklzjiqGl6/2uvfIjXX/sEJ/3iMBkWk7HBouH6dVtRVl4kj4o/XPM3HHzoFFx19a/kUfHoo/9SDErDbUo/dXUlcNFvb+0rgBKUN/UHDw47Yl+cffYJKC8vUn7YSRaw46HBZ/v3ew2j4oEHKP0EXHH5OWJbXHXlXzUHObcNo8KF8391s84AFqOvvPocAZ9kfFz4m9u050ipQj6QKd3H5VedgwMPnIhQyOTry5etxz/ufQG1uxokU8398ZLfn4Gjjz5Qnfncz3jfjzzyKpYtX6d97fRfHo0zzjhGTQjcd7Zvq8FLL76Nj2d/qRz7d5fMFDjB3IHr4ZsvvsM+k8ZoTp17/EzlJYOqBuLqW6/BxKkTBcQyBpg3dzHuuO0hrF+/RdLHt//1Opx+xvG6Ds4pMhYeeeh1LFy0CmPHVom5MnKkkQKmwTkBuP2mjcOLL7xv2BJpyMCaIAY//693P4NJk0bh2OMOxDNPv40nCY7JC8B6C5iGuWuv+RVmzDhY18/vXbtuKx544BX88MMKfdfMc46X/BPBPv77ihUbMWBAGTZt2oELL5ol+aijjpqmseV8CAb9Ws8ENh566HWN6V/+comkn8ioePTRN7Qur7lmpkCPrKyIfp5eIQQmnn/hfTz66Ft48ombBcZQ+um994xU30MPXScwgvc3a9aT2L5jF264/nx5WfBad+yoxdattZg2bRyeefZdPPDAq8qpH3n0Jkw/yLzvL7OexLvvfo0TT5yOS353OiorSzQvKc9Giau773nWUQkx7Xym3rSn0d8CBGLwsMbV0yOg3HqKEDjgnDUKI8Z7wgJDqic5DFJ50IhZYLw5jUE1Y6Y9srR7x0ICAQN+KVCwFsHPZBxoTL2N2bYYHo78GVntqz41vpt8EaiQRQnjDMcoXAwk5zoVRv1EXtO+1zZS22uTWoyjomLyrB+/+nJPJ54SE4VNDc53KObZi31imSMGtGdjhLk/KaWQGfE/vsFITpnmZqMqYrw3WIczcUlfTdJpgFZDsPxZjGygVcNgTdNIeDmR1M9AxX8Y7Z//6n/1CBCosBp0XPyWPmUT1L1BBJuU2EKhCXZNS6XtvLNJi6Ew8u/NErUgCH9vmQmmI9ygvYZiZanX3PCIyhJMMNVgob5kDqQZUDHhcfTcmLjJOM3UdZj48j2SfGJXnRNwcFPg37PIy65HLwEadqQ5XbpEYgm+GLDDp4Ipf2+uMS2NZnb1sOigrv6umH5PPwDK1jBxJYDA95rNmX4UAQWhpsPcbP4yI7WsBweV1mHCzcprQAcWuLnhcUwMFdUYgCtI6uhwDINoKu54NYiqGtezY5BNxNtqFloKHk0VGdAyuJGsAcdVagam8KvxZiLkMD+kR+41jBCL6No5YQIko1VMg2cm9cbTIqlnxS5P2UPSb4LAiCSgjNE2gYrDTju9j/3CceF38vutjJGSr44O6SRzrPhv1JqnBjSZCgJlHI1rvofGyOzkj7a3igbKBFaa8uxkb23Glg3r0dkexaCBQzCg/0B1U1JYitJPve40srLDkhqglIk/QLmXCFLsDEwZRo0xPTJSJ5a5ovFypJ94DQSQGPiyg5RrgcUwBp68F7sWOBelrxzwAakEos312LFxLdzJGPzUOve40NNtzdpN4myltUTJZFd5IKzCjDmUDQuB48fgkUAFi+zsMDXjuafYG2YHpor75mVRfE4C3hMZSbxWy+gxoBvQEW1H7Y7tqN21CyNHj8bAgUNE31QRjl2/LoKGZq2xaEVzUcv0oPxOTnYBhg0bjYxsmvSZvUbRMVEgrn1rcuVclwKE3iTq6mpRUFQMaC7zx420BLcrbVkq3pg9w8jfpBDviWHLtvVYvXgRfOhFWVEhSspK4Q2E0RlLIBbtkM45GRDZ2ZnIzcmDl8UglwfxRHsfUOHzs0DZgk2btyAcycDzL7yMqqphOOa441HZf6CAipLSfgIeySBiYswXi3u5uTkq6lL6ZNOmDWIYsIuYQNjm9RuxdcsWXHPV1Rg4cIB0wzevXYn33ngZW9atRiKWkKdBe7QLfp8LeXmZRTRj7AAAIABJREFUCAe9iHd1YvSI4ciM5GD+vIXYUdeg6x8ycADycjKQFQki4HXDle5BZiiAnOxM5GRmI+Sn/BEEXAR81IQPICMrS6brQSY1Ljdao1HsrK3F0lVr8cXc+Vi5YTNyszMxvLISQyrLsWPXdmTmRpBHY11PUu/fZ+J0DBk9BalgGDUt9Wht69Ac2FVboyD0lJN/IQbF6tWrkOqOaw6Vl5VJq57zdOTIkQ5TzEiwrV67AXUNLRrDKy+7HPW11epotmePBc0515XEOTJjWUE/Rg8eoM700twslOfnojg/F4UlpWK80Ai5K5bA1q1bsH7TBnkzZIT8qKgoQEV5ObIiRcjOLVNRt6s7iq1bNqN5dxPKy/uhML8IEXZ/U+ovbaT5KP3UFOvAB1/Mw/2PPIcugkEBFiGTkmPLyc7DwPJSVFUW4pLfX4hRUw9AyhX4rx4VvF/6vaxfv04+KqNHj0JRUeH/K6CC+yjXkWVU1Nc14IMPZuOtt97G9h1bkUhQFo7ghAGmLVOK3fj0Eoh1pwQy9HR1IpBOYtr4kRjavwileSEBFbkZWQj7A9JnV9cszydXAL3JXsRiSRXHYp0JREIRdfyTycWO6BwyWrIj6OyKIqUu+yBSbi86e92YPXch7njgYaRcLhkBnn7KiTj1tF+grqFeck285n4V5di9uxnFxf0EbA2uGooBAwbDS51+NzuuPWLiyKAunUZ2Lp9zAHUNTWhpa8fWbTvQFe/GpImTkIx3oaGhGvQ+Gjp8FJqaomJVxBNJRDJDOr9DgUwaMKB622osW/45ho2oRFm/QSgsHYmOTj9a2jqQ7mlHc+NWdLXvwLFHHQK3rwSbtjYhECKjJImeeA/u+NMtaCSYEesysmVOxsS5yv26uSWKeLLbxDSuNLJDHgwoztP8rSzOR2lJsRgKIX8QQa9Pvih80d+iqKQUubn58PsCYrN298TRHm1FQ2MdahsasGlbNZav24KlazahIdqNXpcPPeqKSyEc8GJQvxKk4lEMrCjByKrByM/NRktrk1h84ydORfmwKehw5cAbypG8lMvrQX1Dg4AKm2jyPhSXuGkm2qmx45yQtBIZFd3d6oAnlsy4hUBFbk6uvGnEaKrbJaNw7oW264wd+kwgyWIUoBbvQU+yF8lEEu3tLSrUbNu8Fo3Va7Fpw1ps2bgePjc9O5hAG1avL8RuevqmUO7J8TxjsszPS8aQIBPV68XUAw/FYccdDz/ZeR6eDm6kkh6kuiOo3dmKBx94BA1NOyT9lEx2gqbZFnRncivpRTaJxLqo5GKSRMe3iuCIPccU5zoQ495nrWQTCFj0de2bmNjGxtpF6CPm9iKUkSnpOrc3IAk6/jKdi+b8tuCjjLE9buTlZmP0mFHIy81TnCQNZ48XwXAQaRpf01zU8Rbjswn5A/ARnI0RlGFcZsyck2rMMf43RsQS8MON5sYGSaGw4Ew2Lf3HGOsxfjbAidFHViME5dhSBK13qohNibVAOCi2ldjDKXZimv10T8OBMdxk/MIYWHtLR6dicHmT+XwCKkzeEFBzAP/PdcVfZFQQzGlcVyNWJGNnGpHzXihHyViVsQrHSyxnjjsLIuzOFcvMp/iZL8W/6lIk+4m5hTXt3CONyRiOnfiUGeuIRiXJpPhQ8aJH10yZV8btLAbZogLHnnEpm4IIkppmEKMLLkkLMlKVrzg5U7q3z2uMY6z56DQNmVjcyIUpxnR8BK13G5lOVmJWTT+O/KdyJSe3YByvz+s18lEsZKt4kmLDCNndSa0rjhufv8xTGXe5jecf78uwyRkjG4CM42mKNEaCjGALzbQpX0XmJa+X92zWvPl+yzfk/OHY8HOZxzCW4IvX6WGTmcNG577E5gcz5sYnRbK2ScOol3chn58FGd0eSQzxr4yWuRkvPid1aGvsWCiSSY4YlJkZEfQmk8gOR/Dt19/Az+JYD3NQBZ/yXGpobsWuhkZ4ghGwdYtFVD46xi4BR37YG6BUnnnGzBEJZBgJFc7RkGFjU2bX40ZzWxNGDB+BUaNGSDY3nTLzXPlPMKgCOb/ANibxgxh3MSfinJTEcSIhpprkaE3yp7zESBEn5DfHZ8k4jDKJ3IPZYMM1wfnM+cr9nQxheRRSYi8U1t8J3HVyPs5X7v2xRFygKOcBr4P7JCcm9xwx53odaeC4wwz3+LWmpOEOKJ9lPKJSocuFAw+agEt+fya+nbsYD/7jBae5ysjU8HkR+OJYcg9hfm3Hk7kWC3yUiyPDj8+B84x/bo9GdXb2xZMew5jSnu40SnEMuA9wXjOHNLkQz+6wZDStrIv5+V69n36G/Dmyy/g+yvpyLrGBkkPPxieryqBiKvcDys4oBzfr1hQ72eRGab0s1SZkVOyoN0Sj5rv5snK/9s9cj5SgMabCZs9QsVlSMZSi8RtZZ12LF0E3x68DLk8PUuk4siMhBNhYQInE9iham1slkRtj45YbCPt9CEgC1SvmBe+NxXD6U7RGe+APBRFL9qCba97HNRiQbCfjMX4p9xDKxtmir9Yq14CjQsGfYS5MRqwaQJ3iuJkKhhtoW3W0pnt5dpDFbIBlYxJt8mvbxc5nyjnbnaQZumFgcy5znpCFaOMYKklwrXCPJAhx5JHTcMedBgDYM5Y9aoDQHuH45XGdyWjd59X7ORcClCVmRKqz1KwZ1mD66laqoxiAXv6pqrWYlj1JKfXl5KZ73nob2KZbzbduY+5upMud71KDIp+zkSq03yGWpzOvTdxhmAu2McDIeJu9V82DznXzGageJtld05yk+3Y8Zu3D4P4h6UAnxlVTjdNIYZ+1lYDSnutISJljbU8hv4/lwbXqyHnuDarws9Z+yXzIvEYe2qgaCOeCZNWddaHm0m6jbGJiKlP859/bGMvKuhsWmWkCNoAXAQhzzqtGKDbVHlmsvi93fmPiPFMTs99vAH/TJC2gRmwN07CjZl5+lzwnqJDA+IUyTUYiivLCfD/nJ4FwxZSWvfGTL1ejy38AYtRQI79Rc/8/Sz/99Kn9/Of/9SMwSOZRVlbC0J8VvFNGKEmDYGoJ8wDvNgZqPykscgAsxckE3gY0MBuOMRniZzKQYBe/BTds8V6H6482URMIWG19dYBzM7GsAKe7zHadK1FymA88VBjsctGLFeCwF0zHDk1/WVAyJmwMGALcGBzTHibP2jyca7fUfh5MennYoR/T5/Pg4+fLiEzJmkn0zOblyO0gLVmEgvx8RKMdKioxWFKA5HhI9CWvBIgo95A2rBHJDNhxdlBU09ln/p6HMYNySuDwAOP3sttLGu40gRYzgRqORq+XGyP/XomJQBHDJiENlIcuN3kFujTN5jMneODoDbPYZYNKsQikJWWyXlHQCFYxWWIgwQRW0jwcR15bXB4V1PGX/nIPi48pHHnGmX3Fe272lvpnDbY5BgzQLKOCh6pMcX0edUjy+fE9HAcG0LxPmm7H6CmhAM2YV5qDowerV6xAS2OjgIqBAwbKLJl9AUOGj0APGFCboCiD8jg5ufD4/DJEpfyTkh0L2PQY00kGnAoIWTRhAuBIP/HZUoZKQXwsruRobxYQ14ZhQ7gRizZi1/YtSHQ0w5vuQZpjJ/N0dqebNWUDMIu4i1Xj8io5Nz2I9BUJqKDEeU1zZxbZs7Iytc4ooWDmMwtelERg4myQfnUION07AgGpQbmX6bsFFlPJBFqbmrCBsj05uRg7drw+SwENOzKZojFRlI4/i3TdRiKEXYo+PyLhLPTvPwRl/fqrCMPOWb0oBfUfDl2z/yQRjbYLJGDxgvsDC0vGMJ57gd12nSAvbQKSZLobu5t3YfXSxWitr0NBdhb6D+iPQDgL3alexNipmehEMhlTF19eXgF8NJv2BdDR2ax1HY5QBz+IxqZmbNy0GXn5hXjuuRcxZOhQHHn0MRgwaAh2N7cIqOC8IAjHuc7kiPuD7ahcs2a1MTclmyUSQW52NrZt2ozv532PKy67XB4ZHlcKG1YtxRez38PuWhZUk4h1Ux4siqDfJQ3UcMiHRGcHRg4fjtzsfCz8YQmWb9yqZ1lZVixj7ayMEMJ+L3weF3KzAijIy0FBbr5MvBkYBX1BFTy4/9J4XYmE14+u7iTqGpswf8lSfPrNHCxbtxmd3XEMKC9BVXk5BvUrxaqNq1FUWoRMdal2g4DXmPHTMPmAo9Acj2NXawN27d4tFknNzp3wuLw4ccaJkoHZvn078rIzGEJrnrLwzOseNmyY5o/WZ9qFNes2Sv5JhY0LfovG+jqBPzbotXu8BSq4TxP/jvg8GN6/QoyK4qwIyvNyUFyYj/yCImRl5SIQiIidsnTZMtTsqpaUBYHT3JwwRo0YhqL8CmRllaiAnOjpQJQycQsWIDcrF8OqhsmPI0yzVhZqEt1IpLrRHOvEWx9+icef+5e0euFlktStZJ7f2b+kCGOGVuBX552NSdMPl0eFGqn3CnT3Dhoo07Vy1UpJ5YwbNwZlZaX/L4EKJgfG26Cnx4W1a9Zh7txv8dxzz4sZkuwxvhT2lwGiueZNckimSTicycNXUmtjBldi9NAK9CvJRF5WJopz8qXJzbOBBuQMgjl/KEnGJIxyTOxYph49gT4aahcUFiErPxu97l50dHYIYJPhnseP6uYobr//EcxfuU6F8AEVJZh55qk47Zeno273bhWVd+7cJrkzGlvW1TagqKREoPGY0eMRCGSgqzOOoiKyCwp15jKp5z7b0RnH7t2tcHn82Fm7C+vWb8SI4cPRr6wYra27xWoat88ENDS3o6OrB7GupIojPPMC/kx4er3oaKvHsqVfITvXh5y8IgwfMxVt0bRk1OKdLdhdvxWd7Ttx7NFHIBAsw7pN9QiFI3D3JsWomPWnG9HWvl0eOCaOsDFBr9ZhfX0TYt0JgTSUa8v0e1CYGUJFcQGGV5arKz47HEY4FEBWOIyMIIFBLwIhP/KLipGVRaDXI9CIzLFd9btQW7cLO2pqUbO7CdvrW7Bg+Vp0dKeRErWFx3QK4aAPA8tL4OrpwoB+xRgxZBDCIVOk8iKF8RMno//oqehCLnyhfOTnF4L0rF31dSqk2ZdN8GlQT/8dFsNsQwH/zHlCEMLEauzua5YZMj0qCGSQMUSggk0FLEqbuNKwEpig8TxNJlLo7abheQr1ddVobqpFVpYfHS31qK+twarly9G2uwGRoBdBH5P1JNz0LHHMdQkkaK9wDB6TqQTiqV6UVg7Caeech6J+lXCpiEKGXlqMip5ECJs31OOhBx9BtKMBLi+9MjoEVJhuQfp+0fzbLyBEBWi/MT9mLMQOeyah6vTbi+1gpQJU9HB+SV7B2Qhsg4g9c7mfMW4LkM3Fc8/r/xFQIU8uh5FrG0tM4Y1FVsrZlWD0yFFik/JZMW4JR0KS42TUx+SXP01Tenp7+FweFRrlvcVYNkXmhYkVTaJtCvkBl6cPqKDkoMsLARUsZnN+WjkCI7XERiIOi0teTDwPyVzyBQMIZhjA1jSfkFHhFEMs+KJuy6ByEUqadLaxuOhDiACU3w9KP5liIAtHbPgwDRmMp7jueRbvXleNgC+oZJ9nhWUISyaBGImaaUwHKT+TxVrGKypcODGRcgmnm9GCjaZ5h7GvbcwyvnaMFXgf3ONsg5Zttukr9PyEpW6LRswjWAi1Epz2/baBhM/ANnyYHIuxD3Md4w1m8o49YJcx7zQ+bzbOM8W7lAq6vGcrl2HvV/PayW8scMQ4sluFKFNA5WcZDztTIOKcNzGtKewwpmP+IXNTh1krhQwHzLj6hgslnSSfjVUb+yQ3RPhSI5spymqd0PtMTDIjZ2tZafw8M69MUxXnAdcCnzFzPTW6OYwYE/Cyv8VItfHamTvw/lnUlzSJ04DGe5MUCj0DbZMbz0Z6lnA+ML/rTWPx/PnIzsjkBNJ3C2z0+NDU1o7mtg4xdpPmpsX4YaGPQDOleQkyspfPADKMYiGQirlhH1DmNfkKm6qGDavCmDGjFFd6NdxkpZuCKp8nx1kAAiWCVJDt1hqItkcFdjBHlxyzI+Fq83MjK2yYTAJrWDAnMOPsRyb/7TGxvJP7Ge9Gc44JkOKegLTACT4j/hyL4QRYlVeowG4aIwzwZrqydQ1OUxHBEsYPzIFVL6CPEkEyhx1w4PQJuOji0wVU3H/fc87cMqwZzXF2EnNs1fRncnmvJJaNSa/me4DeUcZgWHuksRcyBVMZ8fp1jpoz0qV9i59rCp172N12ncg4mAVmB8jjuc/P5Fja4qhpKDOd0fx8mzerEUxgoAGl7Xjac9LWU1Tc9nLuUCbasM3lu8n5RnBa/lBGpluMRAfwkgySgMIfa9lzjTJm4xhrvtAnrZt1HRoSJtGdaEVJQTYiHhfciST8Lo8amghGdaMHMTLKeCaoPhBHJBJEZnYOEvFu1Ne1YHdLB0KRXHSyEYANZBpTI13IPYEvW5Bl3UWAjYdSjaG+859jzTOFQSnnH9eElcu2dRhzPu4BRU1x3UQlnF9qU5PEjvUuNV3vAtSc52DYckamiHsq/82qTfC53HrrxTj6qP1x511PYfbs7/oAZwHP3C8cb04jSZ4WEKVYmM9JZz/nvfU9taoFBiDgs5fGhT331bRrGLOak04nvJVb2vu+NV8IzgiwNLGY2E8EEfbym7R5vG0WFtNBppAm+bf7OC+Bc1lFeZ0p7j6ghNfDGp/qJ6p3cNydfVnNEab2Z1kFXN88a/qAFif+0c8JGOEeZeIxPlur3qGivZqMTQ3CGnhbENGAREZVg2tnzRd7gIrRR7SY+byXkTd/jqC2WZuGZSAAwkG49jb3Nv6z9p4MQENqvp6T6ncEZ2wDr2FM/PTF2MaCMPYMtiwOxYuO0bUAfeeZ83w03+WYbzugl4kzzBjpUTmSlPYM+59f7rBy/+dF9cVsqnn+zKj4H0P381/8Lx+BqoDPBBjcwBy5Aqs9x8PWsBMYjBgAYm9NNufkNVpzosnbbhpzYHNxGgq1OaRZzLEd4obmZFBIviwFymzGpqhiuqbNIlYgog2KRtkWyDD7kTZCJzji9/JgY9Bm6GomADGdOj1KNhlY8UDk5mlAGRMAKXDlhkuwwNngbbHM7TVBmK7P8R6wRWiOj2VAmE6jXvDnmdTmF+TrezqiLPYYg24lTtTBZbChur8ZPyPnZA42foYpFjNBMNdngy51HjlIN99jftYc4Crq02eh23SMMJDjdRowwGzECiDEmDDIuw1IJQkVMJJK9qATeMGA05F3ssCHfQa2iEiQxZiFeyRNw8ifXUHsqOGBxvKJmBX/Bajgd0tCyaHBEYBQwYFoM5kiNOD0kanQ6YybSZjIYlFyx/nXwwM9qK5kJqEMKtjd9MP336Nh1y4MGji0D6igF8CQ4cNVaM/LzdIzyMrIQmZWNhI9PejoiiHa2SEpCbIU+KIshQ5ZJmcMPl1m7jBgZbGCzyc/P19znwU0u2ZsgmWBCq8nhbqdm1C3cysCrhTSBHQopyDGhunuskEHn6nM0tVJwK4tmmmbQJxjz2dswIqggAoG0QQq+H4aamlupHtVLGd3i0liTbeBTc4tUCHwjYl8HxuK2X0Ksc5O6ejX7KrDPhMmobCoyHQeMmlksuN07PBZMck1HQYyR0EomIGiwnIMGDQUwRA7bh0RjN7/CVT0rXV0o7W1RQldOJLljIuRITNOx3bTNUAFGRW8x550Ep3d7di8ZjW2rl2NkNuDyv4VKCguV4rY0d6OrlhU0mTcGvLzChCJZMPvC0rvnTky1w49RAhUrN+wEcXFpXjm2RcwpGooDjv8SAwaUiUz7aLiMj0PrmEmpw0NLFyaJJJSQxs2rNezyYhkCSzgvrP4hx+w4IcFuPSS38sYtKe7A2uXLcSC775BNyVjkil0daexq343MoI+lJYWICsziFg0ipHDhyE/rxhrVq3D/BXrBGrkZEZQUpCL/JxMZEbYUexCQW4E+blZKMwrQElRobpt6U/BIiEBikAorK5oyha1x7vx5Xff4e2PPsHaTVvREU/C63dhaP9+GN6vDKUFuVi2ZhkKykuRTXPqFJlMXoyfdCCm7H8kor0pNHe1Ye2mjRrLttY2dEa7cOIJJ6KosBjRjg5khv2oranWXN22bZsKl/Q7IeNCczztxpr1G8Wo4Dy/6IILUL+rxmjE76XzzvnEeW4LFXx+EZ8XwyrLMZpARWYE2UE/yooKkJtfqA70cCgLsUQSq1avxvad27QnN7W0IhjyYNTwYRhUWYXMjEJ0xLrUYZYVCWDrpo1oqN+NqiFDUdavUlJXPjI5uP5daTR1deC5V9/Bq+98gvauJNIeJipMmilFkoOK4nyMq+qPs88+A/sfdQx63MEfeVTYOW5ncFdnAgsW/oCWlmZMnjwJ/fqV/38GKrq7ezHnm28xb973eOONtxCNtqqjzKxn88u8nE67ALXFKZ+SAaq4tzXUojQnglFDKzGwfx6K8/NQmluALM4VGFYhi4aRSEAeLuwgi4Qp4UNPAlPk4dyioa0nyG51A1SwEMrnFe/14PUPP8ez/3oH0UQa3qAP/Yrzcd45p+HUX56OlNuDgvwcNLfsxsrlSzVXW5paEYsn0NzejqqhIzT3PZ6AAEF6wAwZMsgw0FKQv8nmLTvQ2t4pkK+mug55+fno378MPncK1bXbUV5ZiUSSP5tAVyeln0JKNr3eCEK+DLELmpu2gbfE9Z9bWIHmloS6WJOJLvQmouiO7cbwEUMRivTDpi318Ad88Ht6EWuNYtatN6GroxadMWMia9mdvH+C19Qy7qK3g+rWaWQGfcjPCKEoOwNFWZkYWFmGstICremMYBhZoQz5pARCHuQW5iE7qwCpXiPxtb1mO6prarC7uUnsq2iqF4tWb8D6rdVIpJhMm64wt7tHbKvKkkJ4ehMYMrAf+hUXqIhW39iEiN+FcRMmYdDYqUj6i+AL5qEgvwQ9HqBe+1m4L7pV15fDqIi2t0vCjXEEz1/+WUXkjAwTI3o8AirIsGDhvK29XSwYJtsEMwRiO4C57diWl1WiF6lEL+pra/H5Z++jo2M3Tv7FcZJFamtqwdaNm7B84SL4XSlkhDnvkkZ60DEyFFChoo6Z8+yMdgXDOO7k0zFk9D5Ie/xiSKlj1s1ChwepRAirlm/Dww89gmSqA2l3l4AKAvTq+HaaPFhgYQxCNi0TTts5zDnOOMXuVaYI4MRqzuhZsOL/DqjgPXIMyQTwh8ICKjw+U2wnhcM2A9l413SnehBg/K5iWC+KC4swfuxY7a2UwlSnpYe29k6XHmMrtxtBfrYjVclYOyn5p5SACqPjbAocewMV6tTOzFDDDmMV7i1ieQqGNhIRxoeNf94DVNALxk8mcia7jxmnmefDmEmFAaejmF/L/YMFDBZd21vaBA6xCEuwor21RV30ZMuyEYb3zTmoZhyXT+8lo4JdziqAu41Ruy26qlJkiylOpz3jHyM/aQEXI9tlNNAZnzhMY2csDBhgh4dFfKO3bRkTamBxYh8j62qK/bbIYwsXagwKBE1hWN2wJm43MZkpONpczAJBfK8pPBqGsQU09gArpjDMF/dqWyUxa3ZP164t1Jg8aU9cz7UpmVE1SJkir43xeT0EMEzxmwUcYy5vGBbspKYclymqMbY0eYg5cy7/4/kCKp5/4k1s3rDNFJD75HUN2MICpWG375HiYhOWcjMnX+GHSlrEkSrRmDlSGfx+ywRXgU0MDC+8bi86OqLyazFNZeZ527ETmOF0qbIoy6K5189x5D264KdHYNqF7775BhnyT6PxrMmzQpFM1NQ3oL6pFd5gGC5/AHE2dXkohxVXHkQGMWX03GIROD4pYqyYMeDexxf3Pt5/W3uLvMvGjhujRg0CFbYQbQuMZhwImMZ1fwKIszKVX3K9MA/uy8PpbajCtxlXkYR4Tx6PGsHCGWGNlc37TGOUKeyzuGxYXF6xjXitBJFssxtzCXU1+01uzfdaINXkuV6pDbDpjQx7AhNck2TLed1GdUC1AOUiBGOMJO6BB+0j6adv5y7CP/7xvJOHMwdNaV6bLmkDVklSmY16DoBF0IS5Js917ZNePv8ONQhyv2EOZO7R+CFxHO3a4DjymmyezDVgGwL5fAQ8O93UpjZg6gycwGogdCRhOL/svtYHVjpqBeYz9qxFK8djgVH7rKxPqI15rYSnngHrMM4eJTBIY2/2MOXJBCWdtcP75Pirq93lBkV147EO+Pz0qGxBRWm+mnvc8RhcBBPYZEYvSaohMC91/H1YSyHDKKeoGD0JsuUa0NwaR3evR6baCUoiuz3opOQlGXVOLYXfa9g/Zm/geHD+2hoJ82M2bOXm56kGxbOV+4zT6G/MgQUkOfUOA4v3sVU1z5wGU1O/cmR0nP2OhV8xZVgzEjCQNr6mXAPca5y9+rY/XyI5srvuegofzP7WdOc74LOK6QIGjNeArVfx2sVccNg9ln2wd/HZ7rXyKxMYThNmx5/Bkf0xNSdTXLe1JivtYwBY7rVGCsyAf2Zf5Vo3IIipjWmfd/wRbNBmOuwNMGEZKaa+ZI2bnXFV44gxseb1WWBS8Yo8K1hodxgDfIbOuagYQGNtmp2NbJOJf6R44rD+LFPOogc6nx1AwLAQDTtwD3/G/J7fu3YvoGLUEc0O6GiZqEZq08ilOWcPaz57gRbarB0Q3LKhTBO0YaYazw7nzO3zPjFy1n1IQ18UvOc3VhJLoZLDrrW/19U7zBjLXrT0IANSmb2Jl9XHgHKuybILf+qb0ffN/0nbyvHNsKyRn4GK//DAfv6r/90jMMhjKEoG4TSdQhbttAVWbSzsfFNAapIwS8uzgSdHwRrT2YK4KUSZjUsBdIBaml1m0ydwYSn/ouWaa3BgCed7zNYl9FmUeociLQMeY4CtRMMpmnLD0Wah4MFK7uzRzOP18ICSZwUDSqcrg9fNhFsBvmO2wwCMF8mNhWwFBQROUZYHDseCmyw70mxwwM+RhA7/87pEG2SxTvRMrw+ZQLIWAAAgAElEQVRN7GIkJT9IE0BDyxQ9XaZCRMqNia4xNzbd7xxfdsIYgMgEOgqYYALybgbeTreTBVv4OdyEmbAqIZRus+kmM+wZBuzGnJsBFz+NGybvy9yLkQ2yHcx6to7cD4MmSiqxWMWN1ibM/L0OuZ6kzCuNSRGTjR4FqpTbSdFcu7dHZtq2GG47q/cGKnifki2S2WOPAmWfOvZciMVZSGBHiClk8kV6L8cnEaNGf6aACpOEduvnF8yfj7rqGgEVAwYMVOJP6aehI0ZIuqiwKE9dnCyQ0bcgxi7iWFzmrBpTARWkSxoWjaSgFE2Zw1GyMJo/fpm9MmCgliRNW20njeluI6MiCK+7B7Vb16KR/gXJuCRK+P3mcGOwbAAF22VgWTb8XOq3iznjGOVyjvDPTDQD4Yjow0zgOb+amqjnbqSYsnJy9DytNIApFpkgg/PA6EvuYUSZ7gTKCfWqMNHc2op169YhN68AY8aONcEf/3M2AnVpgdRzw6hQ4YOgWSCMnJxCDB4yHDm51D83QUg6xeC+D3HYq3uef51ER0ebip/ZWTlIpU3HiknqCBBZbQ0HqHCC/2S6B4lUFxpqdmD14oWIR9tVvOk/cAh8fuqis/u63fFN6UZebr46lZnIJHuMVA7p7+GMDDTsbsS69RtQVt5PQEXVsGGYfshhGDykCq3tUXkrSD5C6yol03b6oxCwaG5uNPqx2jPNnpcRDmPposWai7//3SUyGm5vqcX8uV9ixeIF8CgJTCPeA2zfWYtIwI/ysiIU5GWiK9qO4UOHoiC/GDt21ODrBcvN3uV1I0Md2BynCDIiQYQDLhTm50hyJT87B+XFRSgpKJJHhofdkz4/Ej29aO1IYM78RXj57XexubZWXgk0SQ4E3Bg1qFJd3oV52ViycjEKykqRFQijJxHVnBm/zzRMmDodOWVl2NlYi7i8VJLSmK+tqcMJx52A8rIKyaRQqqW1pUlzZ8eOHRg+fLj8KsrLyx0pFA/Wrt+MuoZmFW8uv/RSbFi72tHp3+PnY5NI/l9Sax4XIn4vqvqVGY8Kmjmne1BckI+8/AIUFBQjGMyQtBKNqmvqatDU2oyWaAyhiBeV/cpRXliJnOxi5BUWIJLpRyTgVuf2kkWLBbyUlpWjsKQEETKU2CXm92J3RxT3PvI0mjvT+Hru94CHq4DJkAGlygpyMWHkYJx5xik4+LgTkXSzk9h0edmzae+IgR2GX3/zjYC5adP2Q2VlP+efrUeF3vWTXzwTjfQTGRUEKmZ/+AneeustLFq0GNGONiMdsZes354CFRM/t4CKYCgDIb8frfW74OvtxsB+BRg8sAjlxYUoyc1DLk19KVPHbmfKOmUFkZuXK6+EzMxcydN4POz0DsDn8UtuiBr2BC874zHJopAmPm/pajz6/JvYWtvAkUIgFFCSfMIxh2Pq/vvBF8kQoyAe78TmjeuQnZmJ1uZ2jBk7Dlu2b0ddfROGDR2JIYOrVKBhBz+fP5PnouJS0Fp50+YdaGyOoqm5HQ31jRg9ahS8XibqaezaVS1N71BGLnY3tyPWkURGToY6Md2uEMK+bK2/aPsuuNwJZGRnITu/DI1NUbEhKTXk96QRDvYa+RtPHrbtbITP50LAm0J0dwPumvUXdERrtbewOUNnhdNFmZ+Xh7q6JnRSrkRyd71at/kZYRRmRlCQnYFwwIfS4hyUlxTJzDwrnIGgNwBv0IVIVgShcCY6OxLYvqMWu+pq0drWgjQZav4gdtTVY87CZWiKxpFKs7PVxBBud1IgZkl+DnxIYujACuRmsDMvjV0NTcjJ8GP8xImo2mcaXOFy+EJ5yM8vRdLVKzkueU44YKFAaHUveyXhxtiCZ/b/xd57RkmanWWCT3gfkZHeV2XZrq7qau+tupFDAiGEH7/MztlldsRgNPNjZw3LYXZ3BsQsi2AYDSBgBAIEkkCmhSRa6m51ta/q8t6lt5GZ4U1G7Hme997IbKmb3fmpPZ06OlWdlRnxxWfufd/3cdz3OPTiWu+Vflz3mNGTSiYFVNB6Y5FARTIhRZZsEVzOGGtCNfvc86sNnHz9JP72b76K8+dP4P77j+AnfuKHtXaXNspYmlvGS88/h8WZ68jEufYpsAJ1KqzEVjPGtwfnqltNHLnzPnzk7/03WFyvYm2zpFooHo1gcKgfPT39CHayePHYKfz2b/0OOsEaOoGqQrtbLbPo0V7WaKp2ZWYLB2Mc4cjWhLYXddauNohQxeMIJf7Z6z7zjrnrF4KdtbVYkm74n0xlEBaAxpDouGwWaae0E7TtsnBdZoNskJLmNd/f24u777oLKZKCaCUVhqztqEk01QfDwSMIurpTn4H/F2BBVa/v602ZQuuP1RVmVNSljrDjN2Utaw/+aZwE57OsbTrYVVQwDydKi7VswtiXLSPVqPZ1dq4aojiggk0/laCba+s6xwS2UskE1laYd1CV/zkJLwQJe3pyqtlYE1FtuXzOrJ84nONgjjW0HwTJOklMfQ4YeQXNDkWMU9YtLhPJ112yohXRxQZLYpOKkWlDEreaG3uXTHfHYlcugmP/83z7Ot7XYaqzXFCmqRLslTxAYc+tvYYxdqnOst3D8gzMMsufb2lq3CDUDyY1BJaa1+y4ZAMUNPWtFAHuTTXYjNmwXGuWU0yzByAZx0AOsvZtKGwEMrMa8Xao6s04cGE2UIdBxKYoF5jC4WjU7HT8oFKDGhFCYts9pD8JVA/QUscN8G2YbCQhggfGlPZ2U5ax4pUbnjnL4TM7Tt4PzGsh4SlFiyXatHCNSqa6mXsanPpr64g7VBnwOVBWGu1NK1W8+Py3kc9kdf55bql84jM6M78k+0eqU9tBgv8ccLJnawoIlM1Nqw0GWalPpVWjI42xPvR2MmaTRcvPDVmC3nnXHbLT5T4hQpnyJUi+owLEwBbel1xv+Xpcg1QXo61rnaH1k1QwLm+lYWAFgQ0bRBpIwmvO+4lgge65Laey5rPtQmR5XaUUo+KA1yKIrqKd4AKvN7/Pnp6fie9vQ0sj4lHVRQKbJScacBigClRZUtyfw9bL0iqKVskN+33uK1Tt8V4lWYCgOa83+2PvYU91iVQpTgkuq7hY1BwMvL2tGPfWq1uWo/nj77Rq8X2sZ6aLnCcbPuZa0q7LemXatPj6k/08PwsVVXZ/mtUVn1UbyDN/zPv229CW/8b725MwPWDmj5WvRVLTTnUWn1nWPPxZgrK8H9SrO8W92YaZsqVcLnUDfnmcAnfCBHOsLw+2g4jHw2Cc2PrqNA7sHsJwTwZhKvnQQZQYYziAdpDrI3cMoELFmXoTKlWSCATiAimWV6tYLlRRawVQrLdQb23JAqpBVZez0fJ23t42y+/LXSIeOhgcGdb1FvkzHNY59IoBs68LyTHA2xNp6C/FDwfSdM7weYU2J+qu9y6rykBdm8n4wbQG6g4w9MRU2QhrwO7zFWxdNttrX4N7ANnudVvLCfRZxgOPiX2QB5XNEtHlOTp3D1MbOeDEqYT84Jz3h81RzBpMZA5ZXhFAsDVJygvutw5o5u9qLXZKAR6D1A7u+fJAT3fH2pG5ILWzA5JYT/PYBGDzT5cNpXsyYaA638c7bmj24o7FjslUmKprHNnBk4b9nEZ2UW7eYLbNzqFCoMVOcofVUtwWzn6DmX32dcu7lt1ebAAYzyOfC/9McT3gMYn06wgz2usEmBmxQ7NJF3DP2R2Jk12C5A7LprezWeJxeDcLA65sHeC6asC+zSREJHUWZR4c3zHu6JLD/X1p++r2ffGWIEkXzOmeku5ffF0i67N3FBXffYLe+c739hnYrWwWC6f2bBQ+MBwwqDDhhqBN23xH9T8FBzr5GBc0J3m3Yn7bq9QGrEGFSNZqxsr0cmq/wexkD/nfpTenVApOzsuFQUGJDq3lfEboqFNxsJlTU+COw3xIuThZvgMLPKk63GZhkq5tL0CThJlNhqyIKH2Tt5EtlvxdSvwlJY9EkKE0X6z5iuS3XJQUChQOq5gwySN9QGlPZEoGnhsOLOWxx3OpAtnsiWyITUAkaQGVdfok22CAhTYHzwo9dNZBCi9yChgW1j6ngD/La+ibChZtHqhQUeRYF9wQvb+e2A1dKZ4BVbKd0p8edTZUn19eMi+lhoohbmA+mM+GawxFJcpDVi/P3VaHRWlTf7K4eN9P/rhDvckMiGnQxaJWTX/QNiwV2mL2NMxOzPlBy5uWHrcKpOaAuaWhCY+BwaK0BujtzTtvYB5DDS+/8AIWp2fFhp+Y3KVhEe2fbrn1sK7zwGBOx0O2MH1GKdmm/Yh5nYYV2Gogng1kfRMr7qBjj9GHm01QTz6vDbFUqahAtOFJwFk71ZFMxoDGJqYvnsZmYVUMIOYXWC1krIRo2GxJzGbKFfe8X9jkxOMq6H2jr3PjNjkyMekVTxsWKkvITCSzmT/T29un17Tnyp5LazY5oDC7L5533Qs8ZjfIkJSSHv11Dsluatj8xBNPqIkwtqKzE3MNQbOxZd7XvKc7W4iFokglMhgb34Xxid0IRmLml61ixg1gtQH7YSybdr5fReeaPudmPWeNjRU42wCHrb7233xJNrflSgGvv34MM9NXMNCTx9SuKeRzvZL0M2CdwBf/n8vm5Out3Jl62QEVMalSZmbncOXqNUzu3o1PfvJTuPXIbXjwoYfRNzCoJpVMe2Vm0BrDBfzyeSWDb2CwX83cieOvoVIuyRZpdHAYly9ewLeffRYf+8Wfw8hQL65fPIMvfu4vMX39CqIKNgNK1YYUFfzME6PD6M0m0KqWcMvBAwLBGE54aXpaYEZnK4h4NI4Eh7DxEJLxkBodXvvebA8G+/oEVowMDqIv34sQPWURxMp6Ed9+5QQ++1dfxMrGppQCfNb4/2wyilunxnF4/5Tu7fOXz0udwEa91qDNSQNHD9+Bhx95F4b27sHZ6Wu45bbbsbG2jnOnz6JcquIDH/igBvwcUPL5W11e0X21urKs4dLU7l1i5+pe6ARx+vRZMcXJgv/Zj/4sXn75ZSl5CN75L3/PaiBHEKxRRToaxYGJURzeswtjfTlE2i0k41H09PdhaGAAmWQGmxubWFpaVr7EJu2I2uZbPDo4hHQiJ0XN0NgoUpmU1vJqqYSTr70qu6PRkSEMj44jk+MzHUEnHsNMqYj/9d/9Oi5emsby6jo6YVooNGRFlYwmMZjP4u47DuCnf/of4eEn3o1QNGP3+nfesg5rK5ZreOaZZ7C+toZHHnoQ+/bstjuaa+oWBwx8Fg2Y3kmmoZpLj1AnjJWVAr7y5a/hk5/8JJaXlxTovLXFQYdjmGt/MaWfX08MpDef99XlZdRrFaQSUUztHsaukUE1sD3xKHKppA3NoxFkUxEFYPYNDKCvbxDJJNfdhALp+SyY7JnM8Do2qmUUimWcuXQFv/n7f4zXT19Ew9krpNMJjPT34IlHH8DjTz2OvYeOYGx0D0gIpjXb7MxNTI7vweUr17G+saxBBcF95sTs33+gay3HvWCjuI5Wh1ZDddQaISytrGJ6dhp3Hr0d8Sh9sBtYWlqQJROzNBgOWpKaJINoPIJELG3ZF7QrWl1BtV4WgLFv737l1PA55p6VSSYRj3NYEEUklsHMzIqUCYlgBws3r+DXf/Xfolxc0N7HplvMSqcCzeV6sFQogNfaGryOzmdfJomh3iwGcglkUgmBFYlYVJZJ/fk8krGEFH+qZRotFNY25TPOvZK1QpDXrljBi6+/gQvXZtHY4lrNgZA1erSWGx7oxchAHqFOE3unJh2btCWrsYHeHhy+7QgOHb0b2cEphJKDGBzehUqzioVFAypsjac60pi3VA4xv4JAowCKekPPOf+dYKzk64CACtZCVL9wb5xbnEaSapFURvY8tNQisMehBe2AauUqvvXM1/H001/EzPRlxGLAhz/8frz3fU9pT643AlheKePc6fM49s1vII46ckmygznspZGjsy2i5Qz3adYaaOAf/ON/jluPPoqb8+saxjOranOFFmCbGBodwpFb78I3vvEsPv3Hn0YnRCIFh6okSZgVo8gorgFlzaT9Nmj1KMkS8mt2SgXPvvRAAmsmsR69MszZUernunkDNvyQXelWW0HaXPtp4cihHFnfHY09TQXpa2xbJKyG5KCRe3tC9p3AxOQ4br/jqMCbjiPXaLd1oZre3kVDTtoN6h63YZQNZgIaTklNGowoe6lRryKdTaITcBZyOh67z3QMLmdOLPIOMD0zg2qljGTasmCSqbj1Bs4+k/WyrUcGKIiFS9Z1OKQ9rrCybPVUrkcDYgIV1WoZ2Z6srgkJJtxLqNoJx6JSUC+cnLManANcDZ5Dsrri0Fp1qBj6lm9nQIXztHZghdigXQbt9jDL295wHWeNutMbW3WOUy14qwu+Pnsnf+9IRR0IqlZlzcr6SPU4B+Gsv53VkTFqDfThz2owSe9958EtRrULkvVgA28DzwzmZ5P1FOtEx6IXIcUNpHS+yT51RDNvwbYT0PZDML4n73XeV5ZPYUCXt50yYIXn1AaBYtbL69zsYDV8dMM2PzTiZ+JrxnTeDZQwX3R6+dsATyCAhmRGHpM9nBu8+efIhlSmDPbgiX/m9D03bPT5HQLmRAYz8Fh7IJXftDBSILxZGPKzUoVFQlUkGEagvSW70LMnT6KvJ9+1aqJiPJXrweWrN5Qp1qQtKS3lZMdkFk+89uxrODCkCwufRaqAfB8ogpFjyFMhpMD4chGTkxO45567nPUTcxJsSM1zZ+xl51ag3teY1KwN2COyX+G9z9wHnn/eP+uFde0VUsM0t0zB0+nI3YD9K3MXjZVvtZZqIK+gEKi4JTBL7gocykVchoWY+rbm8l7jtZTix1ku87OxtxFoJKtgIwbyeeSaYvW6DVU15IMNY3kulNnisyMDBrBxzzN7JPtdzzo3UKDTtcHiWiOSG++vBveYdDfL0eYFVujawNgADL/HcR2zPY7vYe4GFkJuVo7+mLy9FgkTJDaZpZABmt31U7Zszk5KFjdmKy2lVreW2/a+1XuTkOgsjPheXnnEz6iZDNUxzqpb+Swut4bHqme/YcokIziaDZYfdgfaAYHXxY0VJONAtbiIowcnMZxLIUHaHof+zapsTKnBE700FECH96nLmajXSWAMoNmKYLMMzK+UgUgSG+UaNis11AlUOBtrO6eOHCkSG5Vq0EzD1AlGtCRJKJPLGvDqgCTvt+/XQymQZL/FrCF3n3oXCpeJZYRWmx14WyW/XmgALzsqu4a6Ti6D0d8TWtuk+mBOpVnFeftDD2AJhHLgg+WDGijLNc/CpDnLCCunjNdTCiOXh+TJtjwHnPHo/u+CII5c62Y/vqMVEcApUFgHGFBrQAX/w+oIU52pd3cWQzx+C7h2Lig7BumyD3NfygpzgA2XFu/SwLVDqhypwDw52ayJ/HxI660LsrbZkClf7NF0dlduf1OZsMOhRIN7Z42kOSCP35oZd2SOrtyh9dM2UHHrU6tdkN3vRdzDvdOJ1nZHXjWbLptfaf4i8q+RFHYqF5Vz4uoiK6mspvL3bvdkvekvdp/s/MweWFKfpjrCejg/K/V1sV1bA834ebn3efWI9iFHJNj58299DNvflbpRmb6WC/MOUPH/dsbe+ffvuTOwx7MpOJR3ITReWaGH1jWeflAtsGJHQLBfxD2LwDN9vP+mpJ2yZrIgIWNwWzA2GR3cQDyi2X2oTUfhPB9tk/OqDMmBfUaAAsAsuEnMECedFuOo63PnMjeYLeEQVYXnuE2ND7aaevc5eWySpGrztw3AT5m40HEQSna/l3FzUOkDvP0CzYWXCDXZIR6ZNZ9K+ukxRM5AE2NUGAqtBcxZ/Ngww21EDiCQZ6vkfwzEIpDRMF/PiAVtezmsL7r42hxK+4LFNi2Zq3blc96DzyTg1qhus6WcX58GHna+1BCx2HIyPw9Q8AUtPNCaO59RwQByhWlTTdGmHZDZPxlQwcKNOSFkD1pwn5DxHUAFWT1s4D1oQa9Zz5j0n4/gjOwkaOuytipwiB7m4YgxEWrVMl499iJWFxaxZ/8BTEzsQlubWAgHDx3S5xkayKlBIVDBITWLoWqFzN2igAp6J6so8KxSlx9i4etWOK0zNDmdQTaXU2NYqTGElvdRCEHZHZB5yWFEDbNXz2N15qq5EbgbyQ8guIHHwpY3YmwQa0x8YxtPJXQPeTkwz6NJ8pmZEUb/QL/8qllAc0i7vLKs46MlFQsp3iu8Ttwg/bPL+8j7nxIEMtaTWZLxIMl25fHRSurYsRcwNTWFu+++2xSVyh/xgdwEOwJiVfH4GMhGVlo8nMDAwCj27D2IeCoN2m5JrmSlu/3BH/YDtjCbmrquuwJvyajx/seq0Lbl0zsX3E6HDR3DZks4d+EE3njjFQXC7Z3cjbHhMbQCsADAalUMUQ45eK/QWoL3qDGXQkilM7h2/QYWF5fE+PmtT/wn3H7n3Xjk8ScsiDqVll+rFY0BzEzPiOXNc0zQjNeO4MXc/IyFp7OYam7hjVdfwasvHcO/+tjPybLp61/+Ap79xtexub6KoNgcYYV+LyyvIhpPYJyD8r4s6uUN7J/ajVy+RwqqSquNzVINF89fQTJB5nUA6URQvu28KHw/+s0mE3GkE0mpKVLxJBqBIG4ur+LsxSt44/xlrG6WZQuiEFRZTwD5ZAyH9xCo2IdipYTr0zfQ05NHTyqDWquugdWeyd1477vfj+H9B/DK+bO4/e57UVhbxyvHXhZrj7kDBCoYkre8sogL5y/gyJEjuHHtCvr6erFvzx6zxQjT6iOK06dPY2N9U6qVf/M//k/48z//rIF37tny15j3Jc+v7sXCGnKJGPaOj+DWqQlMDvQhQTuoeAy5wbzCxGP001/fwGqhgHK9joZCZQPIJNK6H/p7B6TUSed6BDyRuVuvFDFz/RqWF+aUFzA6PoFsT6/sWFrRKC4sLeKn/8UvYGGBDV8GLQ5G0ZDZTjwUQ19PGrcd3oOPfexf4t4HHkMgSAY7gdHvLg249qwXy/g674HCGh596CEc3LfPMA2Bv/XuYME3APqT/w/wmWNDAbz++im8/toJfOITnxCjn0N5U8tZ8JsV3baW+ObXmvCI1jxalXEoxD2rL5/GWH8vhnpSyMVCyMQYzp7VGjuQz2JwoBdDQwNSnGTTvUjEqN5KISDbjqbW/mK1hLXNIi7dnMenPvNZfOulV1Fp8E7juhNCTzYplv9TTz6On/oHP4n9hzlUzaDJzI9gC2+88ToeevAxzM0t4Vvf+ls9Q/fccw+uXbumz/TQQw+5hoiMqDauz8zi/PlZ9PRMYHltDTdnr+OOI7dJDUJm4ObGGmZnpzE00K+BR7lB/35TmHEYynuArdXqypqATAL8zKThM8w1iINIWs7EqKBIUNGWwuzsEmLBMFKxMG5cOIvf/I3/A5sbc6ppvLWBX1+pZlsrFrGyuuFUaoyBCKA3nUJ/Po3RvhT6enuQy6REMghyXeFgkEwwfgI22hxQyXIwoMETc4LW63WcunAFpy9cRaFE1WKIWcW2r8i7uiOgYqgvK2XTxMQY6rWm1C5Ud44MDSjA/dDhOzG86xYgkcfw2D6U6hWsrDB3Ju3AbLt/bEAYky3U6MgoSrQ92toSKMEBhIbGYs0Ba4WC1u1RB1TMLs3JaiSVymh9qpSrSERTUuKUNkr44uf/Et/4+ldRLq8CwaaGKX//7/84nnzqcaTSPWi3Y9goNbE4t4K/ffpLuHrmOHYN5xEJmYKP65eFRnekCOGoJZaL4Bf/1f+GUGwUlWZY9VJls4TV2TXMzk9jYWkWo6O7cP36DXz72DEEI6xzWthq1tB2wLhXIvG+89YmbaaAhCxMlpaPUpu6fVyhkI6B6Qff3fXLDV3533xd/rt+RsNus0tkPoWGsLRnorWEAyq4r3oGbhf4UB1jNR1rWu7rBKlj8QjuvPMopvZMoSUGvg0SrBE3lr/YoGSwO6tGZVToM9vgjwoj7uvhYAxLS0tSpqYzcSDg8qdckLYNk3YcG0OFHVDBDJlUOqljose5Z+Hzs3PoJpa5q204p+AQknUIFTsFBv2mMsjnelSHF9bWBMDmenKqqTlMzuQyyMnm0myn1s4ta9hFgM0G7rwuNhpQdp3sOtwwxQ1Utm1aTB1rFiqmRjNLXMeK1Zm2mtKCN8kwN1WAndcdygO39kqR4Ni78uR3/QrvG7FL3yJY3Vtg+CBfEWMcw5zrlY5LvukuiNqTxNwQlMNhASsuL4Bv4q1pbBi3HeDO4+bn9ZYmNqiyYFKvsDW7K7t/PPPcX3MRmrxi3ltcOSa7v+fteeAx2LnUsTnVkT/33tdcw2fmQChDhENvO/fKqnA9lz8eG8KaBZWGj27wrT1OOR72TFFxI4sinyOiUOmqwrllgcqgbeU2WM4ah78c5rN/jJD8tLSCcydPIptOi1mvXJNWE6lMFmcvXEY4nkKDgzCBHxEpIaiqqCngOokWh7dNKm6iaLlrw3MjFZUyJ2gLRS982tgWMT4+jnvvu0f1LwEPrq+8/23N2GYgEzCzobzLr3CKIarXuafLb15WzeyzzaqNtmh8X/b0PAdUuPFZkmLfPYesrBXqTnBW19x6Ovn8N2h1RFtjG3bynJvqxobvHrTw9xh/pr5lNszqZ9UHcb0zNRPfh9eg3qRCKuqUArTLMoUa92oDpKhQr8gK0asUfT6HVDsONLHZwra1l4XBJ1TbmJrIgEKeW2OPOw99+e1bnqAN/DmXsH+THZH6aGNLe6tk9lJUMJhtnPPd9xa9jrGt8+j6bgF0cctx8c+4+ia5Rdgz7RnZHnTTPKYLGMalKPM20Fqj3RBZLZEjw1geg60ZAgSoMvCvrQvQQDTURGHpBh5/8C7VeKGtOsJ0c6BKN8h+lmsL+3bCFY70wIykaALNagelShvrxS0BFS1EsV6pocI+nYpwl3/Aa897l3uMyJxunuFzPXh/8TkfGR9DOpMVyJTJrnAAACAASURBVLKzPvV7nO/7tO5xUN4dZhvoo5mDs5XikfLZ13ojsMZAMg/YyMpR2ZpmHb4NQHD9tuE0f9bsv8xOy5NdNUx2hFNvZaTnwmXHWCaVvY6/fnpmXY6nHxht23Xx562P9YN2s4+yGY9/nnQeHEDin0PZfSsLwuzIfX6NX/N8bopmC26P0efz9YZbnFWzOKIlf9fmc7xuXlViBAT7ns2oujkfTjHgwRMppjwI7qwSPbDhP5fmXG7upnvXnVOzEnR5Mo4I7fg8OPP1Pr+V4PD3rbm63+4FEYud9Rw/q0izLnfG9gGXN+UsG/3viCzsgAy5WPjCiGddz6I/59tAoj8I2tT5580+r7dINPLndwJJcoJxIJyBSQaU2F7bLR4c8Oqs3r/jPu+egL/rL07Zqkv6jqLi/9Mpe+eHvofOAIEKDf+1SJrFg2fv+0LQhqTGSOEC6pURkpu5jAMtjgq6seaLX2KecyGU7NyG8iapNAmYQA8X6MvVwmc0qFhqmUS5J5dDpVJ1wIWxHCSBdSHaeh8Oi9gcuPcUc8p532qxdCg8Czi+L4eSXFAs+M75xfH7LOIcLsFBH19QYUnORso3e2p2HIKtPx3zQsFHsrth0BJVD6aKMLsday64efI4WHix2FEhr/95JhWbYLN8EhOKzNcYMyPIBt9mrQi9Zkg5WRSuyPTSPQ0NnGyW58nLpysVyl6NkbIz7MhfL6lU1ESySDarLt+0+U2K11+ARpjNkBUjPPdkjLDAN/kpG2gLe+XxKdi1bWHhtCR570/8mEOUCabEFGLsgQoOnlTgMq/CsQnYSETDYbHHJZmWYqUpRhL9scX8JBOvuCm/U9pNsFnnz21uFHD8pZfkce2BCvrGsgwnUEEmX74nrvs0FksIqOAHq9UY6FwU45tDY7FKHSjgC5GwQDtKoWtiJ5G9w1wFNhbVRlWKCgJZZLMQpCgVC2LPF5ZmgFpRmyULZy9XVSFMRUXIWDpdlpNXQISCslFQhohr8j1oyPNVrJjEnyxWZqNwCLG4uKjrn8/nBU7Qn9uYGqZKEgDj7Ab0fk62yfA1a9yD2NJwwwrgU6dOYW5uDh/4wAc0dPSyVfNeFedJP8fzQXZxhHZikQRy2T7lVOR6B9AmWPZ3ARW6f7YEKPDzeYm7WMoS+rw9UEH7pFa7hqWVWbzw/DdQLW1ifHgYe3btRjiRRL1ak0pJdmLhsO4VWsgEQgEN3vjqvAdo+1RY3xDL//f/4NO448678cBDD8vjPBiJyhKKoYLLi8t6pvv7GUTbr9fmOSULlRknfJA4vCdD7/grL+H1l1/Ef//f/VNsri3ia1/8HK5euoAAw0GjDJWPY7Ncwer6Jqc2GB3ow/hQL2qldUxNTgioIGtvZmFV3vJLq+u4ePocUtEgMvEAkiS5hY1BSaaybObCZGnHtc5uVGqYXljFheszuDa/iI1STTkitMURS3VrC72pBA7vm8CRA/sUqLuytqrzn01nUKlVUa9XMTYwhCeeeBKTtxzCmZvXMbJ7LxZml3Du9Gnkc3n80Id/GLFkEnMLC9gsrovh99CDD+KrT39ZOQz9fX26D5mpwiDUM2fOolDYwB133IFP/f4f4N//u3+PMp89x0Lz2ynvQVkW0Au32UQ2Gcf+iVHcunsCk0MDyESCSCfj6BvOI5vKotMOYnllHQsra6gy+L0NPRPNWlOhvRy202olQMl5LI5Wu4RYqIPRwQHEI9agDY2MIp3pQYQhgIkkvvj8t/Gx/+WX0WqwUYwgkoyjsVVHLBJGLBBDby6J/XuH8Sv/+y/j6O33ot2OahjydkBFYbOIp59+WmGxjz/yMA4dOGAdvfapunkMu0GYB7Rl9wGyV8nOiuPzn/8Szp45jz/8wz+UEonDdm+P4Aes9Gr2DYzfL7jucNjBQbNlGQUw3NcrECGXDCMZ7iAWDor1mozHMTgwgKH+XoyODij/JJfOIR3PKq8iwPWKyqtmS+HOr546i88//XW8evKssiZazhJGa1FPWlkJD953N370p34Md973EAIdDhTquHDxJG5OX8EP/uAPy8KIwboXL15UzsPk5CRefPFFhbQ/9dRTejaD4Y6CwS9fWcLmZhvLhTXcnL6G2w7fagxzNZ91nD17CiNDgxqaLBfryGZ6bXCezGhf5ZqyvLyKcrWMdCqJ/fv3S3UgUJP3WiaDKIGKGIe8SczNL4sZnI1Hcf7ky/jd3/kNrK7OGFjjGKpqrDsdZTeU6w0sLK+ZpZ+GQG30ZtMCtsb6Ujqv+Z6s7CK5FhC45J7adBkJQiBkvxEXg5yA5vnrN3CWqpMys6CCqDKImnJ01kZka4WDGOzLoy+bVKg2ASeCuQTuiuUixkdHsHfPHgyP7MItd9yLnpFJ5PrHUK41xM711k/eEsZ8km1wPTw8rDWee+za6pr2RrJ5fd21vr6uvW10dFT76PzCgoLRuUeyxhITMBTFwtwcPv+Xf4FXX34B1QqJAcxp4JClhZ/5mX+Ge+65G4lEDrFEHu1ODOurRRx/+Rie/sKfIhHuoC/LjAaXm0BVLAc/wTa2gm307RrEv/j5f4N2qB/1trExa5tVLM8XcO3KJaysziOVyuPcufM4ffYMwjE26qbWarusMQ82dFncJKGEbUDKdY3APj8zrzW/9Iy6DtT/bhdY0H66nT9l+5nVywQ8+KcUFcoOM394AhXMJuG+ZyQhew2/JojFzzyGCO0/bMDBrZiqnFtvvQXjY8Pu9xy7zw18jJ1K6ypTffJ6sAbzIckEKuSlHIzLzpBs71Saa5ljpO8AKvyxGJDC2jigTCvat/AZezugwter1uADISoqQkEBFetrBeQyWd2zHLit854tFdGTzzmrsJZUcLL9dErnlTPzOi9U7dgaF7IgZeW5WVKeX0P98N4GSQbg+tdRzeusbrjXcAilehdBrQU8MaylSM5hLe+z1fh5ZGUqtXXV7gsHKiiEdEc2i1dbmBLF2J9+kMP7h78r4oTrc3hP+PO8cz/gueNgVd9zNR3/5vMqpCSgBYyz9vSsWc/ANetVDoKr1qc45Yd6Qa7pzuPcs2X5PjwnUoawLhcYbHkVss6kXZlPjiWA5Ww5RRqq1bXfcP1TkCutRNwe79mu1otuM3N9Zhr7TD+0tufqzbZZ3Z8TuW7bM53XWRkLzpqF97QGg26AaUBgB52WkdXkFc9AWb4fAVcBFaekcOMwlSAxSUixeAoXrlxFKJZEJxRBtWU9tPIhaKHj7JIJLHOftsGoBdT6dUK2Li58lvsS1ROs8e677x5bx0WoM/tYPzQlYMMvXZ9wxGpk15+bx7wDTl3P4JXIUqXsCI73oJm3POP9QeUiiWMkh5FAxBpN4IQbUHIdJxGBim2S8wh2kDTlh4/ejkV2ZcoWJ4AY1Bqmta5F0H1LPZGY76YtQChilky8btzbpMoXyGfzAV4zUzoYMOjJFsp4caAQbaS7pAxnE82D4PNKoIHPnmyfZAfH/L417W8+nNxADVOXbNuvucwap4zzXv8GSlPtYvZqvh/kvc0ZCW2D2TvzYA1osHNoAJ/PxXGsdRfsLOtpr9x3uSnehs6D5fa5zUlCbHcHsPCaSfnurJJJXuR9r/tBId9mhQ326J0G8tk4lmauYHwoL2VrlH18q6HamQq8SIR7TMBUYdwfwhai3qpx7aN1bBDL6zWUqh2sblZQou1rG6gye4iFnluzpAJyuS72bNl11f3LWUm7jbGJCbPqc6RQHqvcKRRsbsNr7a18bvlsOus5AW7aC63G4tojxaOzg/MqF8sZMesuXutuDe0G5j5rybsLeBC6GwQdDrvQdPZIRtgzYH5bocWD473E/Y5fPitC6pEdPYuB33bvmAjBW5mb1ZOut9Q2NuPy6jJZd1MNItWytxbazp7wYBbPk6z2tI8bYCNiqbMg8vbfPGdcC7wjBddG22vMblBgIkEYKo5kdW3h9fx5y/3gHIoqSHsPv0eJLCnSrwutdrZUetYd2OnnTvoZ2QA6FaHLYTXysgGC/NzfqajgmukJAF61458ry9IzxRi/54nFXsHjZxgiYnYB/oBmmMry4J7P+ZiAPwM5zLadFpHWlgXDzm3E9WQCwtwMz2F6tvZ5crUcWZy9lP+7+ze/buzMpTC7NCONf9eXqy39OTPAYzvw3Cvu3wEqvvvUvfOd7/EzsN+x8c3/NaONt4tuahDuimDn/2sMfWNgeBsZ/rfkXK44UjPmmnRJ9bhQSqJlEjkW93wfDvVoTyM7IVdIc6FtkMUQN/9JghRcDMjq7bLpJS224+Tia8WZyatNimxFAP9dMs62FRV+kWfByY+jYsIqCGORezTXh+04lpsvGAwNb+nniXrz9RXkzXNEQMBtrtxgGy0OmfwgN/CmUCcuhmzGeL492mzHa5syNw4ftM3D856BbI6MgbOlTd5QFe/RuF0EKydDYWUm/fPXpV6366TgsmhUoaF6LXf95N/MUGZ3LahSyWTM4oefkUUxF1GCIOubGxoQaGNyC3+jSVaEKUk40CRgIduntlk/cROinQkVFWanYPcQrTfkcU/7A3mv230nRqnLqGDBw/PCa+1BAxYj5UpF/szcwEoVDonbyqigbzOPrbC2gjdeecUBFfulqKDtE/9/gGHaW1vI5xKkHumaxuV5zAA52viU1WTE6WvrJP5WIBlgxtuEx0BGMv+b7C0OpYyVUzMQicMFfo5aBVcvn8fc7DVs0V6k3RKTn4NXP7xQo69Rv/ke7gQqjGVJFro1v3w/D3J4+XS11rQmi/ZkAkzCAioE+PX0iD1Myx1vXeCBCg53zLvZhSs6CbgHUGilweKX13Zubl7WPEeP3qZhnmpI1zSS9clryS8BFe0GBTKIBhnCm8PE5BQGR8aIDGqYYV/fragIBHlPsbGwQFNK2L3tBpmfbw9UsFgHmu06KrVNvPzS85ifuY6+bBp7du1CMpfXM8vgQTZZfI4Z7tyb70EkFtFwweToUbxx8hQ2iyVle/zJZz6Lu+6+F+966vuQzmZlLyPvcGVyNDE0OCQgiPeyD3efX5hHhfkw9N4ORhhlgPOnTuDS+dN44L478cbrL+P8qddR3iiI+c2sAAIVq+sbApyo4hkZ6MNIf05Axa7xMeT7+1ScE2wYGpnA3fc+gGtXrmD22iUkgy1lLASiXO7k0SAAkIArhzVcLpbWi7gyPY+r0/OYXS5gs0xP+47uQ1p6sAAkUHHrXgMqbszcFHhDK5xsOqdhVatZx0Auj4cefBj3Pf4YatEIzl6Zlr/89LUbKrD/4T/6JxgYGlYmBMPLz545g4nxcTz37DfxwAP3o0nlVAAY3zWlUPJr165jaWkFE+MTePbZ5/Arv/IrWF5cQkdsNCvY/CDQr03yaI5HcHDXOG7dPYndBCqi9N+NYHRiAAN9g9jaCmJxuYDX3jiN85evoVJvoiedQyaRRDxCdncWA/1D6Mn3Id3D0PY1XLlyFslIBAf27hLLvX9gCNFECgjHBFT829/6bfzJ5/5atlt8PiKJOGrNKqJsSMK03Epiz+5B/If/61ex/+BRdNoRrS1d6m23XiDADRQ2S/jK019GcX0DTzzyCA7dclBseg9UyH7xO748UFFvcFgRx2eoWvjm8/jmN79paoq2MSg9Q1aNiQZuBqTzWeL/+fyzueZQmfct16m+XBb7d09gIJ9SEDXTpLiO8/wn4wn09mQwMtiH8ZFB5LMZJCIJWfMEwlFZYFyfmcfXnnsRX3v2GG4urqJJ9ZMsG/mZCHrE0JNNY2J4ELcfOYQPfeSH8Pi734tQMCVg8Pnnv4ZkOozHHn1SgEAAYVy+fFnNoq03QZw8eVI+1MPDQxjfNYpgOIbrN1axvrGFxeUV3JwlUHEQiVhCtkL8YOfPnUJPT1oZQfOrVOHlFUKaSqZRrdY15FhdXsNmuaicIwMqVmT5yOfC1tMAkrEoQtE45uYXkaIiIxLC8Re/ic98+vewtjJjwK9Tf7GB46AkkUqKabi8UjByApV27S305dLoz2cwmI1geGgAA/19sk+KR8notWEU9zvum3TcMfZwDNVmA/NLSzh9+RrmltfRoDVYMIJKzZSRGkpwf2AWQ38euWQcvT20WTLG+PXpaVmWjQ0No7+3T6qmux96FHc88AgSuT5Ualta+7jPeyCct6ANi+JYWVmVEo2NNI+RgA4HVwQh1GQSFN2wMGSzfiphYWFJQdH8GashGzh/5iy++MUv4uKFM2g2SwgFuQ+xViTg0sDHPvbzyrNZWNxALNGDPbtvQSySwPrqEv7qLz+Ds2+8hj5my8SjCLIWbJGl3yCEh1agjYlDU/hnH/3XCMX7UW0TSOugUqxjc7mM82dPoVBYRG9+EM89921cvnIF4TgbUgMqCIRaZhQZdlR2mme5mKphU3pWSgS2Ocy3eqvb/Lr6wA9auqoBVyv5obNX3qi2cMMFb/1k/sth2TpxORCrnMoJ1/wbU5LLBAetljvDtZF7pTGm6wgGtnDo0H4cOLBfz53PpPIDc9aBPoCUtWKzaXYhsshw9iRBRGUnx9ybRDJCnNxUt4456pcmG96QaMHaxIAKrikpWT/F9dyZVY9ZXdne7qxJHPsxHIk766dNbKwVRFJiXg1fe2N9vQtU8LPSVpK1DEFF1rvsL1bPzGuIys9OGynef3wfgn9BWujppHEN9Pk/ds26db0byHqPPdkwuGwIeeq3ba/kWsS9lXsj62N7Lsi6tvXVBmf2vqybeE55z2uQyFyIBJURxuzVQIXH786BAARn52F5DQnLrguyBjfWsZjobhApgplTanBNlAVJjCpOY6J7iy32DnxG+T6y+XS5GgTu2fvxWedxkkBFZbAnWCn81Wy+DbhwXt/sy1iPM4+uzeBdkjUG+lEuVgSSkLxjFie08bFQVqnfRT5q6DzoNclIlrc7baD47zbo4/F5S6goczQCAQUj857i/cd/88+ctXAWCGt5fB3lRXD9JcFJtbIClrct12SlQhZup63ejPkzXhGuWptrJTq4dOYcigRdaVe11UapWta9RKDi6vSMSDedcExqZlkQkwXP96+yFwlIVRFgf0PwiyuTC/W247XBpCepsTciOHD//ffpZ2mBzGfHsgm3M1L4dyp4c7mc1iWGVkt5nGQeRK1r02fkQeuRRY6rmCWrV/OLmOfWEw05NeTj2WQ+jRH5+GWZYCFZJxIsJJhPOygfsO4zTATiORKchu6A7g/vKsC8NvV8YQMc+PME+9jzx+IMAm8ob4g1v88p4bPFtVAEQ6eI4u9xWErQhp+RfTfBL+5HlhNhg3DuVbyf+XcNWZ26iooKf78YeGEgmKxifOYl916CHAp3thrUs+F9iDZBOfbEfG0+D7aWmLUQAR0fAM611dbcoJ4LfvE682dlj+X7fipk2DPICtAFdROUdqx3saV3sLM9YCMyoEDSqM6b31e4rljYdAv1agWJCHMo2hjuz6EnFUF5fQWNakWOCfzcS4uLGsQyL6xSLMpwkLUyFT/xWBT53l7U6lvYLLdQrLbQ7ESwslEGJ0QVWu7Wm6i3zPaHjaHlJphtmb7nmPYeJOX3h8fHHGHTnyN3LVxA9M7aX/iNXppghoEAfOZ5Hu0eddY5TmXFNYZkRgOeDIzl37kWFNbXZZe2Tdi0e4ZfHvzg+yk0nkoW7fH2bHD98oAX35fn22z6LEeG97HWXwck+f3WZjJ2nbgH6f6SXRTJwSS4GPjC51U5lPW6A9IY/s751bY6ziukdW8ap6pr3aTBvWpAB465v/t5gp/nCMRpWU6RZmI7yIuy+BPIbr1/q2lZMHpfR7D0drKyRHfzCk/a9YCP6mFnc6nr44BPnWintOMH8KCDqewMGOD9c+brO62fVnRO+YzwOfBKEn+PSCnjLLHUx3OvdL2UzeyolvQWeja7Yo3F45DC1Vmgm3rEKXh8FpcDSOkK4ucvHpTxFluW//oWX2+BOWjPeisw4q1fwb7bBSqsPzSg254x+zf7sXeAir/rJL7zb9+TZ+DWVFqDXjVTCoeqaYhnG4H3xOVmR/sehjOxsHRWEi6wiUM6j9zzWSHr2A8+JT2MsJg2T0IuFB4B16BfeRDOS84L1IWi21PHRsOYfVChxYdRbCiHsJvNEtFZKjBMYswfFpPHeSIqZEeyLtukaD9EloACrB3yLN841xAYM4zyOhv2iMEmxj03GBvmcpH3f/dyLpNYGqpMhrYGRGp4aYfUtqLTefNbk2IbCf9OQIXvK9aLskBMimhNrbElpGZoGhBjS6n9u3kk2gDK1jP6czaMnRmPd+VpLKa4uFP2rM9OtNxbf7mF3DfVFthsg2I25QpM0zDbMVvUWLVQLVdMGixvWAMlZDXCf6tVBFAQfOA559Sag4R3/9iPODkmmcwxDbetUbaf5eeXdRDZ8a2mNibbHN+sqFAGR7XWZdwzH4DHywFWPGHWRoXCKk6++ipWF5awZ99+jE/usuY+EML+gwe1kfXlUyqA2BSSTc+BBptdAhVeUcHz6vMyeG/Y/WRMNTIOBbZFolJU8O/KWKhX1fCg1cL1qxcxff0iWvUSAp0WYqGwjpsFDo/TgwICy9pO6SAJtg9is6IpxPtEHpJbak780FGBcm0I4PNsN/4bgQo2nWxq+H/L87Bhkl1PWmbY/adiz8kSCZn4nyM4wmeYn5usqrNnz+p13//+9ykTRAwGtmgSw9hnYWFVqRUpqkEkSIAtif6BEUxO7UWIzCinwHgroIK/FI2aHFusPYJqzv6JbI/u73zHimtsOeZ1tlBrVHD1ygWceO0YsokIxkaG0T86ps9XLpXFfuFzybWrrzePMFUFboBCFPO114/L2oHNJ4GKBx96BI889rgG8JvlMpZXV83zOhTR8I3XUpYTbqhO1jHPa61OsCaAeCiEi6fewNz0VbSbZZx64zWsLi9Jbp1KxBCnhVssgdXCBkrVGhLpLPp7shgb7EGzWsTu8XH09OY1LGGOBUOB733oURw9ejvO8LVmriPNxz/kLFDI/mnzWtCqJo5GvYXFQgFXZxcwu7SGuaU1FDYrWkfISg1HKRNvoScRx4HJERw+uB+Xr1wWe5DnI5nIoFqvor1VRz6Rwt133YsHn3oCubFRvHjyAvp6+rC+WsDi/BI+9EMfRr6vH+vFDWUOFNZW5Wn/7ee+hSOHb9U5X1icR//gCPoHhnH16jUBFXffdTdeeeVVfPzXPo7nn3uOXeObrrAv+HnM9PONhQOYGhnCbXt348DkKAbZeDSrGBjqwZ6pPYhHU7g5s4CTZy9gemERxXIVsQCHwqMY7BtANpVT1kK2J48o8zsaqxjoz6BaKironh7oQ8MjiMQS6IQTuLq0gl/85V/B6UtXFQjJ9ZXPRn3LFF+pSBKZZBQH9o3iP/7Ob2JkbA8QsAbZ43Ie5DTWDARMffkrX8ZmYR1PPv4YbqUdHeXcfF0yhFy4or+vrMCFAGACFbMzCzh37hJ+7Vf/A6anb6rxNzu2bd9pP2z27G3P8uJrcf3hAIhgBQv7NK//1CQOTo0jkwwDBD3IVCeDM0irqCgyqRjy2bSACiot2LA320EUylW8cvI8vvg3z2JhvYyWy5NhboUxnAiQRNGby2HX2AgO7p3C+3/wvXjPB38AkUgWZ8+cQ62xjv6BrHIvJsb3aE+n5dy5c+dw4MABDci5BnFgxWF4rVnB0OgElpYq2Cx2sLiygtmFGzh6+KCpisCBFjA7e0PDcIIVKxvMeLC1kCo6guRcO5aXVrBR3EAul8W+vfv0+nwf7uEpDkQJ1pDcEOaav6L8jnQ8hK9+4U/x1a98AeuFxW5ekx/C8vdpG0WH7dmFJXBYo8HFVgs96QSG+3vQn4lgaKAPw4P9XUUFgS9+SdHBoZugC1qIBVCsVjE9N49r88tYLBSVTdFoscYIaEgWDJhFCOsVvmY2QaVPVhlZsVgaF65eQSKX1nXggI5ryr5DR/DBH/lRDE5MoFYPY2OTgI15R/PLhiesAwyo4DPsFQEEKjgkymay6pW4/vPccf+hYo3r7eLiClJJZifFsLQwi+MnXsPX/+arWFleRL1WQiBERqExOZU50d7CL/3S/6yBR4FB2GubiEVSuOXgrRjoy2N9bQnffu4ZzN+4TAQFHdqEgOoZDsZa6AQ7GNw9jn/6P/wC4rlRNFhjkNW7Fcb6UhXHX30RleqGLAk/97nPK3cjEOGYkczfBrY0xN8ORzRWoDWDBO48UKHhlAMqTBmw3ZX6AZc/h3446oEKARTOHoRDFQ7D09mcERdUFzuAU29rIIlZ3xhJQiMhkkTY2Lv8OA6Po/G4apHNjXW0WmXceushWe9xAM1Vxysvqqyx5DJmtk9eCcTPRNsb2Ra1mP9CELCAWJx1QMCAbcf684x5vzbzmSOZ4Ob0tAY8rA/og8/al4NQDmh8/e8JT7y/ZIMTt1qIlpUEJmj7lE4yJ4VWf1RUlBRmz1qF+GcildCxsL7n0LJ4aVnnhEQgAbEcHnv7Ow35jP2pAbfL55K9lWPCGxhkNrOWcWF1Ngk7PJ+8JlRksu5k7cxzJuYucyScDYlnRxpoZQNHD3BpAKwAYWP+yvJCntbGKpWy2TFUeUzKaHBAhBFXLBfQPPINGJGf/w7rmp1rPQc+3tLGFLqm2uH78fU41PZkF97PAlyoqiCTv0WA2qxFZNUTsZqOoDS/VJ8TyGOBF3IMf6pMWLvEE85WxSxB+V6sg3ituBZQhWH1MxViRmDzpBlTp1iGnz0fVJQzI4GDaQPW1Ys6MIf3rAApqePNipVDeQ/Kq1R39r1e8aJnjjkUbpiue5mfV0NC1vQxZXFFg0GcP3Vawe65TFrnngOyaDKGYqmqMG2OYDuhKILqMW1dIMBBzSOdKwmYURHFnpo1Fs+pFExuIM5+lZ9Rtlqthur3hx5+UICHQrmDZjnn+1DnnqIBPPdTngvW9bxX+CLsl6hysAG/ebKLPc38jbopfmwdc8fqLIW5x7EWKBfLscTE6AAAIABJREFUqmNFcnB2YsoPCUVAK7d4Mq7hplc5bN9/ZqXkj9U/08rECJqSVeAmLQxplyxAoi0SDEltFjze1H/zXHAt1KrnehXPsudza9lBZtHDA+H580RDvq/ZpRkQJeVTxdRCfA09uxw0h4M6JoW6O9uybbvMNwfs+hVddn8CyqJd0IK9Lu8X3vcCP9wchfZVZsNmtlH8P58h3su0KfQB2d3rKusmI1T6YGb1mcoINRKoSDrMivKkULdGsUbwKgrPcuc1932l1jMSTrZqUl0zr2qrWkKgbYp3XnsSsObnF6WA2zUxjlJxA4HmFlJk21dK6OvLY2xyEtev3cT8YgGlagvVVgB1ql0IIlaqsj+r1g0o9K4X+kyyy3b21FSX6EGy9W5scgLprFO1uvvX1lJzlfBffsbi1wkO8X3GjxFJbZak8a8TNXqQi/VrN4PRu4c4kNjmMY71zv3UWZt7NYT6cZfHo2G3y07h70hV4DIdPQjqe2/efz67RRbbThnCe17PoCMfeJcShd27z7wNQDHU2s6DVA0OqOPn5v4hcFxAgIE8nmFvlmCmivDMfg8cyK7PvZ4ADUeq8H2F2VeZEkM2Yo6Yyz5E/bUjagp8cEHUXRWA+4xcL7oZC86qkK8vwNu9p4EKNmczcN/mYfy8XuHI/fj83w5074Fbn1rp5mraNTZHi22AibWRz9nyyiuud/Z3u6fsenNv9rWAP6Y3nQtXx9meYPWW5nBShlgWjV7DA3KuTv6OkYT9538lUOFriO98LbNg9Nkm23nAOxWMOsp3rJ/e8jK8883v4TNAoMKkpSENADjY5kLqgQd+NJNhGZJIiSobBaohrGi0BdOjiloQKN31CK+kUS0V+/LFd0UBCzYOOIjkarMg69w1CgJCxEKy4+IG7xUHUhC44sUXXJSOsnDjA8uhnFkXWbCs2SUZu4ivwYaDPt62odti5xcSociukeGGpGLZ21m5RcKAEhsaeEsEP/SVXIxhPWLe2ebnUXPlTzjk1jc1xtighzkZWMzYcAVaIKBim5szCw7zwbRj5efRgNl5cSqwk8ctma35Q2tQ7lBnC0c2NoNH7P31koTPgRsmgdwOGmTYGhd9j4iLuRJllgStnAzgYYOgpqvF4EmT+/K8EpQgiEJVCYsEWpjwZ6i44PcJVEi+F6SNBoEKQ7ptaG7h3GLzuJAgIejuc9Gjn8dk5y6mn7NgZza4GzpnBCrI5OP9s7m5jhOvvIKVuYU3ARVs7g/cckifpb83rcaX/tnxREoetMyoMEUFfcl5jQyo6EoqFRhlUk7mQFBNwfuMQIWK4kYFzXpFn2FjZQWnjr+CTrOkjApaRkUjVBnQFiHxJmaYWK+w5k2MPofo87OwGKWljpc/8nrwHEiVIYZ/QAwSDph47Pyam5tVcc3vcTDHQGYPRnWbWsci4ftxkK+N2xUCaqxkrcDi0Qr1lZUVHDt2TOz4vXunXMHmfLBlGWWy0M3yGuj5wk9Ei5psrg97DhxEMkN2rwFwbwVUkE1GWykPjPB88lzpGhDopJWW+/KgkeoBrTksJjpotGpYXprD889+HRE00J/vwfDEpFQlbFwIVPB+y6TTGBzoF1DBekJsrUYLrx8/gRwDFNHBf/n0n+G++x/EY0+8C/n+ftkzGfHMAEU+8yxsZWtAZU0yqfuSaxvfi8ykWCCIq+fP4MLp47h66TSWl+fRpB9qkCHMFqJLRUVhY1MS6ngyjVwqjvHBXmCrjt3jY4gnE+ZL2trCzYVlRDI9+NBHfhTDA/049/qr2FyaRxQNbHXIODOGLM8zbURoQ7ZUWMONxSUsrG5gbnFNORe8r/K5nGw0Wu2mch+mhvtx+JYDuHDpvLGmO5SBJ8EQyXarhp5YHEeP3Ia7Hn4Qdzz6CL78zEvYt/eA/N+vX72OBx58WKqO6dkZRONk91Y0sLxy6YLCIvl+9FIeGduFfO8Azl+4oCbptiNHxLz+tV/9NXz5i19Cq2HsM7u2xnDR0I/yeRb8aGOUgcBTu3DLnglMDY9gq1VBJBrA/j17Mdg/hLn5BcwvrqLaaGCjXMbq8ipCnSDy2bwsQnrzfRgcHkXf4CDS+QRC4bYGn4WVRRSLG+jrH0QoEkcnnMRnvvw0fvvTf4y1YkV2bhy8BCJBNLYaiPEepcVZKoY77jiAj3/8/8TQMEFRBk1v16rWBPjQPwMqvvTlL2GjUMCTjz+OI4cOac3kkEG5Ts4fmedAgPkOoILe19/65rfZMuEXf+Ffo1jc1OCCAeaCsV2jZ3uf7ad+/eK6wXOpIPlKRXs/jywWCWHfxAhuP7RPtmMpWnu022rqKXbjVkSRIm2FqNRJJlLa1xudEAqVBl587SSeOfY6NqtMCXBrScCCpQVUhGO6/lMT45gcG8YDj96ND/zwDyKV6MexYy/jtqMHkUrHMTM9h9uP3mOhfu227J+kfurt1XFzDdI9weFyMIT5uRKKZQiomFu8iTtvv4UYC8KBuBaGYnEds3OXMTiUx2aFoG8amWxWNYiRAAJYWbaBLH3w9+zZo3NCOwyeU+4xytuJRmU1tb5ZRC6dkOXan/+X/4xjzz+DzfVla7w4hHENMfdhDR7CEYELXO9kIYE2cskERgZ60J+OYKA/L1CBg1kqrGg9wmtFZRqfdzb6Wp/aHYXCM5x7Ya2EUq0jW6mllYLyHrZILnDB6Yl0UmtDJhFHPpPB0sISMtleXJuZQaYvh1QipWtI8kOmN4/H3vMUHn/3e1BrxLC+vqm8JZE23CDZWNZxZXdwOOb3YQIVHGLSHk6D+3BYjF/+LhUVPIcrS2uy/pifm8GxF57D6dPHUSisoLXFGoFKQMt94LrPZphKvJ//hZ/D2Pg4NkplLMwt4tSpc3qP22+/HaMjg7JSuXD6FOrlEs6dOIEQySoKkadGv4NYJol/+N/+c4ztOYImFb0cQmzFcePyEs6cPq7A7kw2j09/+k+wvl5Ah/eSy6igooIn/M37i9FDSELh4FEDMMe+tqbZsrx2rln8nie+UB3BL6/Q9SQV7kO0fuL+S+97Iw1xP9oBVDj2oVh0HGyrMDegAm4ox4kx61u+Pp9LAj8rK7OqiR555BEBff768E96w5M9aNeR9YYHNzuIeJ9vARUrWCusIZGIIBILqNbhl7et8efIhoUcbncwPT0togoBvp1AhT3PHdWxb7Kv5CAvZraUzAYjcEtFhUhUwaABFcUi0tmUhq6BMGsdrj9xxGO0EAxh6dQNW48IXDiyko6JNZUGPr5WNna6iDXOk9wDC94P3AMwGhDJysYGxkScWTdbCKgFPfuhrkABvZ8Fpmq93TFssyBrZ6nkSEJmAbVtB6S7x9V8GnxKxe0CZBmO7voqX8Nr+M6Bu2eO6te937dZz2hQ6noEP4zxPZ3seroe/3pxhZYPDgwaeE01hDJ8eN9a/ghBEqlxaJMT7KAti1fLA6A968bmpuWbyKLXgqsJYGltdHubqbi3jEjlsqjkKe6yJ6Qcke2IBSuzReS6qqGRz20LWPCzf/ZkC6mcOwM51FM68MX3tLLy4DCczxjBFx/qDqpaSFazgXKr3tS6eer1E6goNJnh6AZuNLaaoGHvwtIqWiQ9BSMGWCiHoa38IfZGBAYsOiCs/ByqtQQ0Om92PcICw9wAilap0Qgee+xR9Y/xGK0PzXGAL27AlJGLPDuY/RifR8uV4BC7KUCSdZut3QaE8IvrfDKVNIazC/nlNSK5gXuUFHwu10MKS7cGNOtUeiRRa1hNy/VPNkckyPnwV7f2qd90vSiPh/0aQQHZqnAPI7ilEsvCrEmaI2dJwJeAIGOds3fXINoxsJXHqCwMy64gSYT3h3oWkg4FXFm4sWocBNVTs4/lvalg8fV1y/dj3k4qIRKAJ/p5Bwi77wwY8Mxz/6zzHiIxznIcLcvG9x08Ln+PqVZTJo4p1vTaLkNF9jTuelpehilI+PsiFBFw93WebHnN19/stOxZ0PxBKiQCLqZWMpDOgD0eh65dd41jjgHB5y10GmWkoyGU1lbQ4bUjcEqySTyJYtmuOckELfbV8ZjZUDriGPf8ldV1FMsNbJYa2KSFaoj7agglZlSGWRt5cp1dKw2HOdwNcL21PsnwfquDJ6d22fMtFarlnWjusiP7yGYQXpXhcEdakDvFnAc1uO5qViJVq3f+MCcA7VfdMHV77mzovq129uuI9mXeQz4HQcCCAWI7yaCadfF4nWKZr8V7w0ABG4bzmBLxpFRP1jL662KDelsDbO2wfBWzITLyrctHcsCOZmz+M+rzUGa7nTvUzSVx1nhdCyJXk2ifdjMmrmPaO1wIO8H97rrkADKzLbS8H67fnrDr936SUf1sSmuM1IE2Q9J96dQUZtdmSi4/p7I90+6Bbmi3s43S+Vf+Ywenv7adUXHk3QXLUxLQb2p7n7EkW1LVTLbX8R7i+RLRS9k+todaVscOcFMzPvscAo3dOTVwytaRriW9s930ChHfk/qAdQ+CdAtA37u+DVLhiSzf+fOmPvrO7zqQR7Zhzlq/u1YZSOWv9ztAxXefu3e+8z1+BsYl5bXFxTMpvOzXL+4eHSVIwcWK7Cg2q5JTalO2QboHKzybxYAGC7LzGzmLBzL7xdYLBMWE4aZhG4A1e95uSghrKKimxgc3cyjCJp6LrDZ9WjGwgCbTzZYiJ5HjwmMDcDLfudazsNFwlqqAuBV/Gnw5VQN/hgucDdEtjMoj9JREGqJtzYnP0JDEVYwJV5A4ew0umFZEGNKvhdl9Ni7aBjZsqchkgc2ClGGuYsE4OZe8B8lo2upoEMDzwHPLn/cIu4AisujcxsP3UeGp4GRjc6gpdb6C/rPZRs2MEduwPevPswassLVBuRUSJq3WZheEGhIy5vzgzYoMFmRbKmYpfSVD28K0KWs08IJ/f/ePfsSaPxemzQGWZ/ORKczX4WDMXxdv0xNxhZ15b/pgNAadGlBBFp4BFYNIZxgo10SptCmgYnl2/k1ARTAcxS2HDmkwnc+z0Q3Kr56MMQ51mefBxrjZ6iDmGnM1Su58apNyWSps4skm5TXtWj/Vy2g2KmJmnnnjBFbnpxEPb7FtcJJVY7rzvhcqvyPXJRIyX2UPFkqd5FhDYRXwdo/y/XiN+dyKQRiNKQiaTHALXG/Kz51DI4IU/H+frD5M9WCF7baqRuwQx2Lqsh9Y5JHNw+fMWYCRgX3ixAkVVo8++rAYw05RrsEHN30eI+2XGEqKNp+lKGKJNHbt2YeB4RH999sBFQrsozVbNKpr4If/9v6WU+G/uvdtF6jgbWPS63J5Hd9+9hvYKMyhn+z48QkNP9j8cMik7JNoFKMjw4gmLLyU91WpXMGJN05ieHRMTdGn/uDTuPue+/DEk0+hp7cXzQ4EYhQ43GozRydvVmWU5Bc3xVzmOtekpzHPWwdYX17G2eOv4uKZEygWllBrVOXnTwlIMs4MAEqAYyhsFNUEMxMhE49hbCiPUKeFfbt3yetXeTnNmpqEczfn8Mi73oP3v+99SIXDOPv6q9hYuCmmFIdFrSatYzgsCYjRuLS+ghsLi1hYXcfCUgHVujUODNzO9+cVFJwIAbsFVOyXZVON7EUxXRKoNioIbDWQj8Vw2+HbML5/Lx7/wPfj8twmotGE7NVuXL+B++67H8lMBjdnZxGLs2mPYNeuXTh35rQ8x6d27zLWajiKSCyJS5cuY252Hg888CAWFhbx8Y//Ov76C19Acb3Qvc6eVSQJtkICgWC7ib50AlPDAzi8Zxf2TY4jHgkpo2SofxD7dk/J63x1tYAOZdMRG1Y1qmb1QJA4nTbVRH5gAJ0o1YJNxGgjt1mQ4oUWXMFoHLPLRfzG7/4Bnj95kk+wGKdUE5CFXVdAYQipWBp9uSQ+8IEn8S9/9mcwODyJAAflQTJPbYDpB0XGSAbWNor40pe+hPW1NSkqDh+6RYw7Ng4Nxxr0RbZnYpuignlQAfzpZz6LQqGI//s3PiHAgc2D1lqneuR7mrTcBmK+uOZr8fscONAyxNZyrmlbGBvoxaP33i7Aoi+dli2ZgLcqWasdJJJRRJXVEEU8QYZtCOVmB7PL6/jWi6/h2RdfR6XO91IFoSE0G24PVPTl85iamMDo0AAOHZ3CR37qI8hlR/DqK8fx6KMPiXF7/Pgp3HfvQ3o/njMOFfj8e+UZPwuzNeLpGGgZc/HSAiqVIBaWlzG/PIN77roV9WoT0WBCzNZ6o4RLl05iaKQX9S0C7CllKhA4YU/EQp9ARWGjgHy+B1NTUyJjUBnA99oJVGyWqyhXaujLZZCOA7/7iY/j7KlXUdxY1aCS50oWL3EjTZCFlchkcXNmVvsJ6xHuHVQ6jAz0Yqw/hXxPBv2y54sL9CIownXKW0PwXMvioN3BerkkwCKczCEQTqNSb+H4iVNYmJ9Hg4oaMl7pm5xJY7i/V3ZS0VAYaysFxKJJrDOYNBWXuiPUDoDMeoQDGN0zge//0Iewe++dshTjkNnWaAO9pPCJJBSUzfrN1xWsBVmfEPRlk8X7SkBFIIDB4SGUNjZx/LUTuHj+Ei5dviBFRalcQKNZQatRVe1mTD7vTUzLsaCA8J/4qZ9Es93EwvwiXn7pFeVhUB3Qk88iFACi4ahA6JeefRYrMzfBmIlgiE1wR+SDW++8D7fd8yh23XIQ8UwW1VIHZ964htnZa+jp5TA/jt/7vU/J9o+m9O1OQwAp9y0/gPd/GjFGOKmCtBu1up5TTwSxoZUxkfV3DmrkH0/moCYSxhp0gIUNnR2A6IAKhmlruO6Gcm5GoWPxw7OuCliTmSC9p/QMciDK54MDYyn9tC9XsLy8iL179+p80ubBgpw9UGENMIeYrIX8AIA5J6ZcDsnai+HqyVRUqgoO/WyYo8Co7nmywTTryY5lVHQVFfGuooLrL4+fDGQ/cFUtyuFMJK7j53rkgQqx87mvbqzrnkplCHzExU7nUJcDS67jzOkoXV2yLLxOEKl0ykhLVWe/yOGi8kFskEmSgHlhe/W02ax5e4+d4c92XW3AavUxvbt9Fp8pJ7o0YUcXtkGwY8MTJHb2I96GxIJdLVxT7FvHdOex+aBsAfOOJKZcOGfl0z1vziKJ64xXX6gGdwMiG0S5TDqn/uU9ZwN/DgYtPN3sbTgYjyLC32/be505c0YZMxpi086WylwSXnp7ceXKZVNn894LmeUNPxMVM7zGVJnymO39bPDGGl+scCLebnCrASstp+oWaM01x6vISLrhII3PJpnoVHtI9eI+o+8T+fkF6lYquqZxqZQt+a9ECxuXC2NAA0EP5hrRZpYWKcZUDzqejcJRCQxttZFOJHDi5VexubamNVSADol3VIi3O5hfXkUnQNQ+ilqTnzWgc+iir7XvEKgJBqMCc2Qb4ti4vg7gedCgWuR5+/cnn3zCHT97ABuG+zxHDt27e7pTHfjht7IaqQSJksBFsoK3IvKsYyPeUeXAutVqKnNLoGXaxsa6PoPqD1prIaB9j72EagceR8QAAB+STkDB1yeWpch7wBQXJDQS1CGwwXuAeAyfG+9hbwHiVSmjCKz4ftk/b/w56zlpmURQgWof9gA27Od78R5Rv+mAD79eUiVoA0rrF0ggKxU3VWO3mjVZTRmj2l6bzwyHzJ4M4uul7XuH4KrZY/P92Sd44oxtCyTRmN1yNE4Awmow2WLx/gpSWdDSPWzPgj3//tzRwYLrql/bjQyJrlLI1378Ptcp9i48H96Jgb/Pn+HaRGtb5X24WYVmGOzDa0VCZqhvbiDQqEkdWqvQuo0qoZSUlcx85DWlwntrq45QBKrfqfahinJjs4I6s7ACMbQQQbHWQICAQauJzWJZa65mDH4IvyO/iRu9t+Tmc8xZwNSeKdUqZoPVUM3E88bPsxNU9323f/bF2nfXTlmKDjDQuiKgwGY7Pl+0Cz45iz0PEmlvd9kBBnCYO4SRNg348c+qgYOW+bHTYktKOdkCMtyeik4DiG1fo9WQzcd0PzTsfhD+5AhL+jen8NAar0G71Qye96B1yQWv+3uSszO5hDjLPD9/sz7D1SBOCeqVIrbeWA6Qz8Xgs+ezGTQTcqCXgaoWfO/zXfz51z3M3FERoAxQ5xyOx8C61c81dtobOadym+W5XAdz4iDgYvkt5s1gMzye15NP57o94G3vXXfWWZbD4ddB+0w2y/KKCltPvUW7rXVa/7lP6e8eZLH1XjkeOxQXBnjSGi8o8gfrW09q8IRfr7zcSSbtHuyOv7ytxdPbKC3eCqTwL2cKDwPhBfxrduc9n2zPeweoeKur8M73vqfPwH7n9ek3fzH0nc3QTtmxZ8NwYSLrTZJGj/S7M9Bl7nvGhhZnUy74AYNYgS7Ih008NzbPLJNKgYhp2BQaHKKIre/CBrk5sPnh8fHfFDbdaKDeasg3VMitGhAWOAQi2HiatJpfJstkkcamzIobvoaGvA4t9QFn2ry8/IvB2Fsm1bbNx3nL+qA4g8+7Cg0h91x4QwRdLBTMS/68H6WX8HMQwaBQyZmdMoEvR6YQj4sLKwEK71VOpg7/nQsnN3dDks22i9fQB35Jku58yY3J1enmfnhptAp7/Z6FdHuAyQ+2uKHyuhuo4MK+5S3rfCi7+RhQQcrwW22IQcpvaypEmNVAwEIDNDInO1v4vh81RYUV0iwODX33hYEf9viMikat5hpEC8T0uRo+WJdNqTW4G2KxjI2OKki11WygWinjtZdexsrCIvbuO4DR8V0IsHkLBnHo8CEdX18+q/9OysLHgIpypSqZOgdLZOjJGsy99zbCbtYcZIeTNSHmPwNFFU5Y0iBmfn4a05fOI0L/VDew5NDSy1vtPrBz6+2QohEr9nyx5YfxYmM4CybvPcx/kyqDx59MI5PLobe/T0UnO+srly4LwOnN5+QhnMv26DXE3HCDErF0HIPX5qn02bXBkT5rKGTNqgtnI3A0OzeH06dO4p577tRQjwwjKwCs+VMQV7OOGoenDniLxZIYHZvE5K49iMRSxhh9i4wKgl0eqOD55f8JxsiOjF7R8pBUOeYqMqeK4sSrYxZUvOc4nDx37jhOnXxJLG56wI8Mj0ltRZZvpcKw6w5GRoaQyefF2CLDaHl1DcePn8buvfuV4/BHf/hHuOeee/D4u55ET1+vVDepTAbLqytYWV6Sdy+ZsAxd5/1WLm5gfWUJs9evoN2oiS0/e/MmCivLqFdKaDcbKFdLAic5lCAAzKE3n3EW+7weVHhQdj0+NIBwZwt7p3ZrKMDnis9SIBLDyfOXkRscxod+6Edw/30Polmv4Y2XnsfizDQSHMoz/J0eqq0OKtU6FgoruLm4iPmlNSwur+t7nqE4ONSPoYFepMJB9GdTuGX/Ppw5ewYdDu3l+U11GpUEWxqwHjp4EH2D/XjPBz+ImxucZyXQaG7h+uULeN+7n5S6px0MY62woGHSrl2TOHXiODLZNHZPThrbiI0/lSZXrmH6xgze+77348bNWfz2f/wd/NXnv4D5m9O+2u6uxXZPsjHhQKqJOAes/XnsGx/B/slJDPf1KZCXg4Zd4+OywqGdAfesdIrZSE3Eo8xVyCASpXVaXAAlg34VCB1si6Vfox3SWgFNDnLbwOf/5lv4s7/+ClY3i2a3Ag4lYgIgmgQqwiE1KgN9PfjZj/4Mvv9978Hw6LisyOR56+9Y30G40dbaZhF//Vdfxsb6Bh5/7EFlK/CHGSRt4KSz+XMMfduTAgKzllfW8Nyzz+Nzn/sCXnjhmJoJ20uNne2bXjH4XDFvYL0xvzjQ4BrKAaAV38ZxSsci+OEPvgcP3307tiqbyCYtlLpWK2nPzCST5g0fiTFdDrVGE+ulGq4vrOCZY6/i+dfeQLNjjHDaLPB4ZOkXCOoc5XvymJqcxEBfL/YeGMU//ic/hf7+UVy+fAO333EXU3Vx6qRZPaXTpmbToHAHM0x2NY0GStWiMiNu3iygVA5IUbGwPIu777hdqioFd24R6KhgeuYyEKiht2dQmSMhkgSiKXSapqRcXlvFmryLM9i3bx+q5aqUBXxGOXgLR4LKstnYKKFR30JvOoNUtI3/9Ju/iovnT6BaXpNlXalY1nCNA2N5I9eqsm27MTOHWt287tkCMlthbLgfk0MZ5HuS6OUawtpF93fYQhHbFjKqPSicRL0TQirXi7FdUwincghGE9qnfvd3fw9XLl6yPZhD33AAPdkU+nvzSGdo+1RFvUGFZhOxZArlrTY2Chsa9ihrKR5DKpvC8NgYxif348DBW3D06FH09fVbkKuzBgrHGL6+jmQ6rc/GQVNhwxpIqh1Ya/G5YOaKH9C/8O3n8dKLL0jhRpZ9vUY7Kw6qaYjlw6et2dJQgLVUpyPFyxPvegKPPfGo1JKvv34cN65fx+EjRzAyMmxD9U4QQ319WJiZwQvPfB3pWBiREO88NvtbCMViyAyN4J5HH8dDT7wHiwtlnDp1Bc1mBZlsHPXaFj71qT+yeiRklmrMqGA+jrdB8A00nyeqIUm42CwWuzWlTRQcSBHcDvkV2O/qStZoysYSwrodbO3va9axZHeT8ewDWrf3NwNyuKdyn7a5uAV6UlzYIZNYgw1T+orZTpZsLK7Bfr1eRr43iztuP6L7mHs17y8CVBymElgg8Gp1lQ3YtL6StkAAb3VZCiYqnci2TTiWooYNbiBs9TWPw5TLBCrK5ZIIIwQWkomYbF34O3x2SUSR1YtjQUshF7WMCqpBixsbyKTS2jt4bglUkCCh908mNGj0Sg0NE2JxFC4umUKX6zPPD9c5ZT9FnWc8M32MAWs4gjNZcB7tImqIbGOBoCJoOWsZ2YqwLq+aX7nISk1jtvtBhK9hzWaHxBxHxXCBr77O5bW0XL1tqzCfObETvDFvd/sSO1QDT6vzPYNUDGxZcxog4XsA9Q4RDpjoc26WMeqX5IXubXNsmMzzyj817C9uYO/ePcp4uHn1mgb7HNT47DoC+s2a1TRcd5SJFqeXOmkjAAAgAElEQVS9kd33ff39WJhbcMCHKWS8zYmOo22gBJnurGfIUDdVhSEFPA7uY9tqwLCAXsu0s/6L/84/PRGLgDIH6iLvuHBxHjdfT0QxZ6+kvkbgGgE+Y6aK6d5uI07VpGxng2iy3yIJKBDAG6++jhrdAxzDn4SHlshYLRQ2y2hxpQlGlFUh0g+JJMwsVAA7911TGMn6kXW/iGE+R9HcByxgV9xi/Umggo8ylRl+7+OwkM+LLJQdE9znGJjdjAH5vM685/1wldfaiE5UwNvP8d957xrhicNzku28YtWA9q4Sx4FNVj+w7gyJ5OfVFAQKeM/xmniio4b8UuqYkoR9cJOhzFLV0Ekh1nVMUH/OalGDQhvo8n00FG40XbAySUR2Hnn/UMlKIhm/x/cgGOBBXFlMuQw/rnHeEojHK+snrQdBFDmsdyq4nXZrUilI0eBmEdz7lNFAcmZBvbpZRZqqn8fM91ZmBoFd5WfakFMOAzzvjmCn59jNRnQvd8PC7ZrqXLoBvVlI2xrl5zBeCSPHBmc54/t/XmepXhgcz96Xn1cET2fx26TLRAN9VKR12igszCuHiPVAiyBNLK5nvlwqIR5htl0YjXYN0YSBFDyGsfExzM0tgbf3erGBWKoHTYIPgTDawYDIq1ybme/oXSx8eDTPFbc+nRdXDPNaTu3ZrX1hp3rRwsctB9Jfoy7w4Opn2ZE56yURQZ0DwY4JvVnrOXWaX1f53ySp8Tj93tv1+XfXi+sBe2qeS64ZAo/ddeR9rewRV1Pzdbm/0Cqa593uH5IAHTjbHcLbINzfM7ZXGzAikhuoZHHqXrfoe1WA5gMOYPdroIHjBoi4wsmUJG5PFrlEczz7XQ8+7CTUysaSGSJOrePrHQEOqguD3VpFe4YDvbuEZBcS7QkcAvdpOewG53pPB/boPiTxVgCfXVuvOtbvuzLQyM2WUcHPcnZHRgUVFfy+z5nw4JUnQut6ggQuF0guQoH1Hdo3OIPhvNFZsWnmor7CWdPuALvkjuL2JFP4uJmeVOKm/LIJhO0jlm/0NsjD2377v/7nrT72FpFOPcbz6eaPcnl4x/rJVU3v/PH/mzNwMBZ3DY4FwO2UtvkNkh/Wsx3IcKSnZJdl7zZ1LdgqDg3RfhPDyFkoCbl1DHK+Njd8W2yMeeI3Jf8nCyiGJUvS5hdUL+Fzsmj/npx3GsPdJH9aTMho0gDe+786ufoOGb1UC2IgbqPgKoCIvEqeTEYIwYltJJyouaRiRIObBsRoU3QLJBsE7aeugeVr2SCYnvVsDo1FpwKnURcLn74aBCv4fTLETO5trDbPpuPC7ZF87xNqqC6RVS7QtjmaEsSaFvNttEEPGzvv18gPbECRNXYsZgmOKIiTRRoLXDYNbLgkh/avYwu2mIHK+bCAdLEiFYJdp/hO8loeG8EJnjuFXJIF3GnhvT/+428CPzyLRcWfK+K1edP/kg28/m6yQm87xc/kGassKmhNVK6UlIkxOjIiRgjfmxkar774ElYXl7B3/0GMjhlQwYbj0OFbUG/WMNBLix9aP6UFVvAzsxBmw8w6gz6zfqP36hMbmrWxvrHeZa7wXCYU/BxWqG2puoGLF0+jsrqAPrJfOEQMAk2w8XJenbJ3sOvMAYIAjPC29drOgpb3qg+AV0PqADF/fVPJLBKZFHp6+8S0pG/+9atXsb6yilw2hYHBfuRyvQhF6YcZtbbIhRD6xobPmSkrnMUZC2KGEjrWhgcVqXQ4deqkRqb3P3C/7lnCV2RO+8KKkbD0N+W15xfD7fI9g9i77yAS6byGOG8JVLBhDNFixsA2sprZiMpqjsOULlCxM4jbDW/axm6hhUetUcTSygz+9pmvIJ2MoTebxeTEbsRjKTE6qbbh0L+vP4fB0QmTpdJLfnYer504hV17bsFKYRN/8ed/hgfuvw+PPvYEevr6FEJPlc1mqShbIx5f7wBVPMxIqKPdqKC0toTnnvkaLp09g0qpJJYTm1+F/WngUUatUtQAleeU946k5c4qhjd/PByRl38sGMTU5LgLY2xZo5/N4vLVm7IhuufBR/CBH/gwDh0+gulrl3CaNlDLi0iEOqiT+dtsyVN5sbCKuZU1zC+tYlGKigYoqSeoMDSYx+TIMLKxCPJpBkLvwtnz5xBJJLC0WjDfY9oJoINcJoU9U7uRz2Xw2LueRGz4IGZWyzh55qx8cH/swz9gg4V4GleunEdfb06huG8cfw29+bwULAQUE5mMnueZm3O4duUa3vf9H8T07AI++7nP44//8I9w5fzFrq/pmzdcFv0cRPHIWxjoyWBqdAgTg0PYMzGBXCqhIVk4AOTSGfmtc7w41N+HRAyy/8pke2SvRaCCgAWH7gHKoNFAEy2UN4sorpdQ3wIuz8/jk3/yFzhx5qKaLV4vXiteM4GXbYb2RcSmJCDzy7/8S7KempwcV1HtQeBuY+w+DNfMtc0S/voLT2NjfROPPX4/jt5GoIKJBLTZo0e55SNxT9WghwsSi9VABC+88JLW7o9+9KOYm5v7f9h70yA7r/M88Ln71vfevr3vaKwEQIIEwUUUV1ELJWuzZItabI8tJ5OZuOwfjqtcU3b5R2bKVWNl4iSOkpkpx3YixR5JsR3JskiK4gJS4gIuIPZ9RzfQ+3r3fep53nNuN2gqlb9KsV0wKKBx+97vO9857/s+W0cxIVaTU39x/xAQ74BIn8fA85fvn8MFAtb8fg6PWOTXy0Xce9cd+Ge/9b/KemxtaV7qsGC7jHKhiGCDbFNTAhKoYabK8loJ12aXcfCNw3j16AlZQTFzhYxmngXeR5eB3GTmEazq7e1BX28Kn//cJzA4NIJoNIUdt92ORiuMmZvzOlMmt4yp6dvctPq1QPZupVZEsVLHzEwR5UpIQAUVFQfuPIBmm1YGnBmFUCpWBZpduXoK99+9H2u07WGgdlcPGgVa3oWwsLqE5bVlrY9dO3eiXKxgjQon2mFwrcSCiMQjWFxYAZpB9Ka7EGpV8P98/Y9w/fIZNBt5XdP1tTzy6wUNHrjnUfbfN9Ajq5B6C1JjMNAzFg5jfGQI28dz6M0kkeYQloGjAsVNEdVqVxFOUJYfQTzTh2277sDOPXciQJu4QglHThzHiz96DsePHUWtxOBQqhGARCKM/p40Muks4okkllfWxLpvMF8rnsDMog1+WcdwOMhmm78rGyEcRDbbraHM2Ng4du26Tb+oHAtGYlgvMHcjjXq9JWYyw7Kptsik0trbuN6K6+s4fvwojh09giuXLyGfX1ZGCNeZwnTlM26sVDWSBlkYGOV+8Szlefehxx/Dgbv34/KVKzh79qz2EioExM5shgTyJsJBvPHqTzA3dVXZNVHar4SYVQG0E3EMbt2BL3zlH2N+qYLLl2fAcobqFaqRvvnN/8+aUoGCZJ6WVCdtABWusZbPsfnY069drFdnjWX2WBz+bWSP2UCGgybLN+Ch9l7WUKp7qnxOyjrjNFhw6uLNw3SrOQ0MoP0hrx3DgAkmGyhk79MGywmBW6l0FqmuKIYGc9i2bYuRGnjKtYMiZCjTqcYJktn+0IqLZyffqwEVASwuzymXhAqNVCqOGC3G3pWfxU8qoIIe8g6oIBBPoIIDGP4i+M7BJf9eIaTyvjfwRTaIUaqjwigWSmL2phJJ/WKdU1hflw0aAWcOzUlESTKjImEWMVzTy+fnnco0jqisLAyIoJIrELQcDqkctKdaEKW3RNKdclY3qnF4XVkhEVRUmKj1FBp2a9jCga4NPviaNVq3kujgrIOo/OR9lA0LTynXk/Bzc8+1QF5TaHiQ2Pvqq76W8mTDxsWrH7SPO0kpB768Nh1ilGNYEijhecHaSf2WQmZrAmON9GKB2ktLy1JIqJdgPgLBjWgQA8NDOHfilDJ7eE5wXxgdG9Ga5zA0NzCIS2fOIpFIYa2QR99gn4gf/QMDWjfnTp5GOp3VnsLro+un4GaywY3MxOGSkbiCNsh13vVSOeiZYUaT2fYSXPBWV7Ibc97kcgKg0ou5IW5wqF7JWVT5/kZD+kgEJReKq3pZkzHeTwNPuP+r9qIKoFKRmiLQauPVl17G0MCgrN547bjP8ZmvNVs6u+scaNHIjwWrhsfs6wKqWzqDQv4de2BmCrr7521CPG/B2NO25h579FGB4tpedH4RbCBAQzAi6jLlYqq1pSTQALTWsQsMUV3vrE74Hlh3cn2mGARP+1q9Z+4TERGSBKaXaP8U135l6oWomNR+TxZLnRlA3Bv4XepdLZvFFDf6TjdwN6KhFNu04OFgl8RGDTGtT/Y2Vvw3BtpxXVso++bcRHnw1+21CMD64HcfSm39ckx7g1QcfD7d63hLJAXwVu1Z4PNJYhl/HnsK1j56jtoEMow1rR7LoYy856zdeRZ5iyxjVhtR0w+LxbS3TcRmGm6QaUxtt/4dn0pZAk7dusHsNlmhWN/KtSCpgAQh1oE1gf8enJCykWCUzhwOpG2fEIGR5ERaeHINuHwc2d416wihjkCziomBPoTqFWWwyHECYa3nm3NzItyQbMPVWqquS2VIMJHnDUlGPC9L5SaWV0sIRknuiaNUa6inpuWbZa6YTbF32qAjhLe9Zj9PsqhFbgUxPDrUeba9qlLZqIRVnErdj3N9/qjY8uap1llTvkY0+x9JFDrkTQ3kpVClIpRKGlPweQKpgHmeF7pvNpPxdlQiebo/573xSp7N9noGRpp1Nofepi4zZYJBkP6+Wl/f2cPbnC04qyoHoFLNpCwlp5bz68nXvP6Md0vNKaLsNb0asAPAuBmTADTNHDasCPxn4UU00qhd5Y6aRHZ8Vk9sZEDYkN6DyL4m32ytxX9jahdTK/F3s2jiGjQVH59RPdfOhmFznoV/Tc0R222c3mz99PEVWxci6ZpbiVefeDtsD055gErAic49A2X17zypRHWn7VvvBhn8XNBfA+6F9j1mV2UWkRbYbe/V6j4/r/Hnsu6X7/dcZohmSe6/O33tJgIbX6ij1tA81REo3H7T6YWkLPS5FfY5xd18H6i4dVzw/v/62b8C212joKbPDS35APLBFILvHw43dxcLqGWeijwcWNxwYLHBgnEydzcoZ1HPpsmG0Mba5INnmyKHs4bo2sZizHqPLPOg8g8tn3aT/Zq/LJ9JeWqqwG2ruDBQwpoMXygJJHAekR5ltiwHY8ircHeou2cq0L+eBxUPf99YC+QVu8FsiqyRNGk2axIfzmN+mRt+fZS6ev9Mymr9BioJuPMyZbG0urrcGQZTnmrsErIufOBQXUCCsYh4yLLoN3mksWFC6Ep3OU9BAjYurMwVSXaQkplp9gD6UhaIXVMPgCj3gf7B7qCVx6gDPnitLWzPZIP63GIlWdHA68tCkg07Cz8CEywKCW4ZYEE2aR0f//KXO/Zem9eBoezGolDOiAMqVAS6Q51Fmm/sPFBhOQ0xlCpFFff0Mo/yYGrUUCpQUUGgYqEDVNDTPBgJ4bY9t+n9kNnLXIqudFZABa9zpVLTsMkDFV6uKxWOY+wQbFhcWpTtE794b2QnEomgXC0iX1yVF/fS9UvojUQ12IolE2iqaa7JGoi1A5k/dphS3RNVASf5rBs+eFaMV0/oOrm1KwZgu62hE20aYqkEcr29Ct3mUHD6+nXMTE3LWmRgsF9ARZTTWnJ6XRXFRtQDMW1XzPimVoqPsFkTqPHYJFm+PnUNV69cxP679mNsfFzvm//cWFJtDd1Y9BHYZKEUCvE+dWH79tvQ0z9CdO+nAhW0f+J95c8jm5MNMhm2Co7/qUAFbYCtUeD6q1QLqNbzeO75p1Ct5NGTTmNsdBw9uX49w6bAqSp4XSHfoRDikSiuXruOYyfOYnh8K2ZmF/HM00/j4Yc+qEDtnv4+xMi+d0FjwXAES8urWFpaxNjokHznL5w6ipdfeBYnj76DtdUVsaQYWsd9jc8qvV7pdU8pNq2iPHPHN+MCiMEMhgB2TE4gReuksVENN9n0k8GcymRw/cYcbswvIZbK4mOf+BTuuGu/lAj7b9+L7kQY89PXEGjUUC2XUSjmsbC2qvDd6ZvzWFopoN5soVguqanNpFPYOTmGnlQSfZkuTIyP4eSZ04h3pTAzv4h0VwZVPl+BgAEVk1sw0NeDnbftxn1P/AIqgQQuX5nChbPH8aGHPoB0thv1QARnzp5AXy6rMO3Db72BgYF+DPb3o1QuoruvD9V6HXM353Hx3AV84lOfxuzCsgCPP/njf403fvJq56z4BwFjLMhCgsYESIwP9mDXli0YJBDS1yurhsL6mgbrmXQXUokEMkl69meRTqf0HNBmhUzcRIIgWEogRKlVwVJ+TYzRerkhi62fHDmKb3//GcwvMwNnwyPbgArb6zjAI0D54AMP4Pd///eR6UpicnLSWJQcLDp22OaKgc/fSr7YASoee+wDuOOOXWJLh4NsygtmfaDm3jyYbb/lXhHFt7/z18j19OC3fuu3NFzgF89MMW7dc+qZbZ59xn2FA36ziOFnt5wp7h/j4xNiJy4tLiCViOJXf+kr+JVf/hIGenswNzON8soMqoUC6mTg0mJDoagtFCtlLK6WcH1uGT9+6x28dvQkOC7P9fSKnTo3v6D9lXsM96Te3l6MjYwItErEgUcfvR+TW7dj9+59GNuyHeVKE6ureZw6cxr33XtAdiB+z918/aQIo5VBvYWLF+dQKocwv7SEG3NTuOeu/bIA49nTbodRKdVlN3TsxGt48N47UWHzyUDtdD9q6xziRbCwsoLl9SWtFVNUEMykPRFBnBSizAhKRDE7M49YJIrB/hzyy9P4v//kj7A0N41KaU1nOMkLZF9y7yTAUSgWkOvLymIhlclJhcJ9ngHaVD3MXbuAdDKGZDiMRJTwLvd/Do3bCMciGJmYwNadt+H2u+4VwJsvN2QR9/3v/x3++m+/g8X5BQGkYQ1AGkgKgKIlEm0Au/U6M7MLOt/Ipl1cXsPCyrpqGc9o94pXDVgiNiiUhV+Ag6g4BgYGlUvz8GMfFSBLRRIbMAbU5wtFWfKlEmmxiAPtJn707NP48csHsbK2aOrKWgntFkEKhrPbgNhqEiNi0DLQmlp0rEdIQqk1GOCbxL59d2D/XXdhZnZW5+yO7dv1/rlWeF+CBLcbdZw8chgz09cQZdhyqIlWoAnw/U/uwGd+8ZdwY2YNhfUaIjGu/xhmZhbwzW/8pSltBVQ0UasUTZniVKRWg1qt44EKnt16Ljc91/KMDpilh8dbCArwOrKepD2Rfx3f7HvwktkiHAR74ogNIlzws/td/t0kMtBKgmAm2d0cVIWoYnUWpo7AY7lVUYSjMakpRkYGsGvXNjHDNUjR+mJtakBFm6AY67MmFRUclphKg4UdgQqyZQlUUEkVoXrSARWeZML3662feLZO32A2VkEKEakgEjHVnsyhE9uXILn3qXdABcFiDm5YDxfW8tqbkjGz9amUi07NQC/3qF7Pv3aYLOloFCvnFzTIlQUKA7W5vkWkYiKMDY7ciLoTSu69yD2DUqQjWVA4qx43MDK2PIk5FjJN5YbyDWh16ay0+Op+4KFBVouDqIgNHKUcMesQriHWsfx+eZo7O1H1Ik7dYXa8Vpsba5fDLxKGWFNxDzf1gNatC/W0mtApRjYxsvlGWH9TPmO9EwEzrW5dbyo8CewFBVA10Z3LSuVIwKhea8gOanh0ENnuLn2O+cUlLMwvK/+Kqpz+kQGRfFaWVlAuV7V/0f6SSTzMqPEZZ7JNIgEraP7yuuau7+S+4Z8l2XS4a+KHSP65YV9qzGF7Fn1dYAOwqIHuHNwytJiWfWkOo20wzesr4EMENAOtrK808IxfBMCoHoxw7TdbOHbkHeX4RMMxrK6tqZYi8NsMBHFjbkHgBDNiGrzXYlTXzSqVwCRrBddnqp7XMN682X0d4Rnxfl/hG3r4oQcRS7AH5LlPpXpN7m4i7jSaKFZqzo7WwuGpWuRJSPWoriF7OOaT6TmvISjwuiUljOyFaKXo1CcRetaTbEaFBSwXi8Aen+tYnISPomp5rj8CqezpRKwDLYFiKJbLqm+lApY1Di216CNvRD5eARK+pIIoWzg8X9+eN9qccUhsCiWx4uWJb6xoKbtJtOAsQgQ2gqe2D/N68nywntHmCexbk8xxc+oyr8wgqCHAjlZBtEZ0THbfX/ge1A/9zFHAB7yb0od9jHp3X4PxfrvnntfOs8N90LFmFQ4Y9M+3HyAb+EaGutmh8Us99aYMMdmZCexx2QghEjut3/dOAjav4T5tVjqatcQt7JwYqywG3aCZj02wXUWtuIqtwwMoLs5Kvck9gLZltWYA8wuLiCdjGOzLIhlnjgtfxJRBfX0DyPYNorCax82bC7jJ3Lc6Yf0wKvWWcO61dVpOUQHVBOEPKZ9lxaebJosdASlcs9wcQwFMbLGMCtlMt9rKJOJ9tLkGVXZRIzxSpeOyFzhH8rMj3wdrNiNQ2NaBB4r4b31fpb2XtbOrx0X68QC1wCz2V1z7Gxbk/Fm0tPSqIVqk8ey3DB4jhOoZlruFqUX8rKBjNehIpLIQcuCxshB+ypdXSYjI4c4fqTR89pCxcHWNeM/551IpOTsjrmNzS3CB0a5/8Op5v3/6eovrxCzgOHOw+ZpmTO53s2YyMq7PDxFo5taunl26LdT8bMS2VgODzD5d9Y4URGZJJuBcz7UBn/Zln8nPHfnzTv9oI6Niz0cXnVLJVEYeBvKzQwNOHXnxp17dW//CVEvOGs/ZRdFVwdR/Le3j6qUIqNbqZvvoziZPNhbw5ezTNcdxQJjv2Qy0MlDBqztsRmFnjgc4O1fB5dzptTxg5Ug87/X5bKfcCEZ/H6j477z573/bz84VoPWTZ1v6B0/BVxGGbFW0MfnizpQDHLYbesfvF4vKbdj81Cxu+cUmgq9rAMZGsCeLC2PhG+OIm70xoK0oMR8+G6SIeeGQSm6msn4hw999L38X018bjb2mmt+gefd7kMUzFXwhbEWyodzeW9WHBvFzeQaqAp3bbfnd0iJIrBXKZCVhtE3HiiFDizmIp/WD3rtjpLMQ0+uABZepErhZ871yqM8hsRhQHO5rEGzvicWcipS6hbvpQGRz4sKpvGyUB7w1zFaYqIircWO1xlGZFwy94+HF4WeEwIp/3+YzbpusscHYHBo7wdYwmQZkhPLz+ZB03kPvRdoJwnO2ARysmLy8Jg9DNUgBNhZ1qSn450986Uu6Jr6A8weliiondt8MVAihV6AvBxOVDsjB92qqkTBSXUkh7dFoCH29vQjy4GzUUMwX8PahQ1ieX+wAFRwYcZC/a/dOtAMtDVxZzGa6c2q4aPtUrdYV6uiBCv8M+KaT64RWOGvra8hmsrpmXBumqOD7LKFaL+Hc+RM48cZrCBcKYqwPjQ4jmU1rGGBMZrKIPOOCvvmU7Vph5odz/FlSyoTMH9pLL8XWU/gZ5bYVlMt1NMnETyakguAgcO7mDK5fuYqe7jSGhtls5uThy6aEBSO/xGbyDB8GHFLm7oKv5KsdDIod7FkC/uevrCzjwoUz8m09cOBeY6EYD1UNOwth2m9VGCou5Q+bmTi2bNkuEIAhzz9NUcGBkUJo223Mz89rbxgYHFAj898CKsBIDA1zCVQUZZ3y2usvYWrqMnozXRgaHMbQ4KjeY76wpiEa0MSOnbt1fVkoX756DafPXUb3wAhuzizgxeeewyMPfRAfeOBB9A70Kz+CYeyqv4Ms0oCVpUUsz99AfnEOh378ItaWONxhAGhBBRXZl82aWfmwcN+5c5vC7egLTEUGP6f3WlYTTkZds4U9O7Yr0JhABd9rIpXEwtIC+odHcO7iFVyZmkG50cbO2+5QRkmj0cb/+Yd/iIHuNH701Hdx9cJZ1Mp5VIoFLK2vC6i4OjWDYrGugGkGJLJoZhO8Z8ckhnqyAtRGhoZw7ORxZU3MLBAoSon1yxDldCqJyS3jGB0cQDSRxOd+9Z+iGe3C1OwCTh8/gg8cuAtDw2OotEM4deqIlBfj42M4+s47yOWyGBsdtaBVsTkbmL05j3Onz+KTn/ksFpfXFVb+9X/zJ/j2N/5SLKj3ZJ9wAE1FBevSVhPJaAg7JsaxbXQMw7kM0l1JDZPpL13K5+Wp38Oclq6oclqGh4aQyXaL9d/VlRGLvtqoY7VSxPTstBRH1VINU3NL+P7Bl/HCK4dQJnPMNQjcD2x4ZKFuHKaSBfmLn/88fv3Xv6qfNUTbLhbUmwaavjngc8f1s1LYACoefex+7N27U/tBlFZaNTbYIQ16WDxrUOYUFbUGcPDgj5UV86d/+qd2rgQCGiwQtPDPqA3t3JmkAEaz/uCf8fliODW/nwqpdDqjgdT09DQKxSIO3HMAv/7Vf6TskIG+XqC0gKmLF7G+MI8ABwUOKGLzv7C0jmtzi3j5jbfxxtETCEfjmNwyqXV18sxZrK7TZi0ghjSBitHhYQ0VouEWPvz4g/i5T34a5UoDsUQKiVS3hqynTp/Gww89pDPVnxWbmxo1rkF6HQMXLsyiWKR90zKmZ67jwF13odGihQVrC4ZgNlEoruLK1ZPIpduY2LEN1UAUuewICgvlDlCxkl/SMJaDcFo/FYuVDaCC4E40grn5OXSl4lhamMazT/8t5m9cRmFtCaUCQ1c5YGjp2WdzybWVL6wj05NGVzaHvfv2o2dgCP0DgxgbHcbEyDDOnzyGp77/d7JrS7ARqjfRPzCM+x54ENv37MXAyAjaAfrktrBWrGDqxhyOHD2Ob3/rmzhz6qjWP8MyuV+0m9ZYp9Nx5LIp9PT0Yn5xGdVKA5nubkxN39T51gqQ8cj9lzWU1YC+/moGXeCnADFj8WvY2wKy2T4cuOdefOyJJzAyMqo/W8vnte+kE91Si/z9338Xr7/2CkrlVVQqealFyQq2uoCZYda0Wv3lahveRClINwgkZuFhhA4OyfkMb52clG8+FRXduR4UaV1Rb6LVqCJFr+zCGo69c5WwB9UAACAASURBVBiLc7OItMlADiCUTOPxn/s0tmzfg+tT86zEEIkxpySKa9duyvpJikEHVNQrRTf8M4acL4a8f7UIF8672ggGBlhY3WRNrRNcClQkO9kDFZs9s7mWPRmB943KO9Y4HpD0Daz/HmtyLZjYUVLN+95Zjvj6lvdSKhkqxaIxqb1y3Rns2rkd4+OjshziZMmCTx1Q0eDa4dlqigoOnMzYwIAK5sEQ4OU+GZa9k9WrrDH9l91Lszm9cfOGVKWsVzph2jEHVDSa6gu8HYcpKhrKqOD75pCbVl8JgsiOrMBwc9qpMSid+y5Bf6+oiElRG8bcqRm9P5F7giRXcMDMvcOsIGWPJNay2XVYXoZTLTgGrwaOslK1CQI/HwesfE0SrsguVn2vQb99aQgjglTbAlr9sMfZXOl+yP6F2UNh7be8LlQMmO2IAU2efevk4M632xivrNNl58cBqasFveqCoIdIVbTLFWmMjGC7L3x9I6IQADQL10DQfLrZY8hOSEBFUFlYyVREQMXU9RvKxqMtIOuVya0TaDSqqvUWFhdx+swFCzEPhzE4Miggd2V5Vddn5sasPcvRKPbu2Sv2vuy0CIq4YRt/LvP5/PCVe4wfNPksQQ+ii3jWbKrO5Wf2QdGys3I2XH7t8/OzR7A8GGPy8tfq6prOOgLyZoNlNkRyEXAZHQrRrtcQYxZQuaxA+WNHjqBcMBs/3p8d23dgcXkF1UYDZy9dkl0ZrwHtc1iMyAKVn5GscpIAFWZuWSBSd3E+64by/H5vHcJnUjU4Wnj44YcExHHfq1ZLiMkiqyQbNK7rBgPdNSQMivBCm1lmoYHB7OrzgqhpyBsT6Mv7y3OFD/s6VXSsW9RTBNGkil59YlT1uDJ3GI5cLGu9sSaNJ+MKojYv/Ja5HDjmPJ83rjv+b/aJUk7RhreQV9/HdcF1TxWUPfNuvTuQyCwqjYHfIUsRMEqSQEHQ1/zYlc3A54egNO9bzWycZLkUtr6ItY/mCupvCbxaD+GJglT9qBYiGFo222PtPQ489DWGDX9twM19iGQQDl15//3ezD7ECaJ0lvkhrf97A7UNhBfhknOUDut9QwmgDJoWrcQIQphNE0Fc5UM5i2epFDQktbOB15GvyV6FdRrPe1lNOhttrnsO6/ka7AuNgEkwuoRQq4yx3m4UlxZkPbm6WsDA0BgKpQoWV1ZEdBgZ7kO9SpKeZXnwenAvzfX0Y25uCc02laurROYEUlQbkAUU1yZVelQZtZgtxvkOzyuy0AlsO2UMgURlK4WCGBsb65BCK6xLnEWZKS9sruHnN2aBGdVn8+CWVyionnZMeX8fBWZRacJuUHMhe964h3iQgc+QJz4qFFmEPANF/KB/MxGX64zZVLZnO/sfnYdmLcafx/XF9eCZ97wfnE0YMObeh88VeNeo0JNlfXi6kSUso1Jr21mGqUd0tnEkF3m1kO81PLF3c33igXQBaC4nhf/tQRA+SyILExgiYMk9kjWgcwuxa2wzOV1HWUTSAcKIq1IDETzU3M6pvRyYJ0DJZUTx7zjH47XkOaBBvrsO/v2bcg44/Vxf5wrd/sSSZcFq3mY2fQJduNe5jKR3Xc7O//xvuTJ5Oz6zkovITt7PJEXQ7BBrLKNWz7JC0wmocrd1BBtv+e7+t1dFyM7eOc/wofa2Xz6bw9uVedDd1B9G7PL3w5/lm/tH/+G8m4nUN7xu7ysqftoyeP/Pf1avwI5N1kDaBF2SPDc62SGJtWIeqZI6MQvCIY96kCj1dgwHSXZdKDaH+t6qxgMI3OQEEmwKEeIP8QAJN37JZR1TwDd8vrH1vn9kM/mNWRu4/A9ZlNpBL/kZLQYY8OwCekT6d4cDNzXvca3iy8nUxAB5F9OPr8NDhp7Puh482FwR6jcGASZkQmqDMV9I7/mpoa1ks9b0Cf0UK5cHgGVfGDBjwUWG8hPAcR6rAmXYdDn/TrFQDEX3w2U2PywSNNh2XrGeaWAFmxVN3NfJULQD2BBeARwcRMcYmEpE2lhG5mfrC3qz0OLnUtPmB2YOUNLBIYZMQ/0zARiyYljU8ucRMCBAYVkVTXzsi092QCX+O75/z0qT9DsQVNHJIkdhpG64oZC4WkXvk9ecjYtJZSMaevHnkInvgQoW/bRwOfTKq1hdWpbl0Oj4pKTaDDzbsn0CkWgIwwMDYpZTrk5FRanCwPcK1ulP3qLtkYWXcy345po/n4x8PgM+bJDvg82sSZGLKJbIls/j1ReeQX5qGr2ZjAbdmd4M4nHK4sn+Y7FtXqwELXRtHXDhn0dfUHtQggCHL0D0M2UxErXhKllJzYZCkAk48PNfPHsO6XQSIyND6O7u0YCY68sDFWSWeqsYy1oho9s8gLmuAhEbyppE1AEB8mit4dq1S5ibncXdB+5FT2+fWWH4Z67Rkh1OuVKU9Jw6Yoa5dnf3YeeefWIWm80ZmwsOpaz44T3k2mFRThbK7Nys1tfg0KCeI14nY9e48oYdoKooEgI5MLL/0WxzuLGu4NSXX3oOPZmE8iTGxibVeK6vc5DGAOIatm7doQEqf+a1qWmcuzyFWFdWQ8FXXnoJH37sERy4536ku7Ni4gc53KNNRdn2nkYpj1cPPoeXX/ghZqavIpWI2ZAyX9awnY0ri1TaCvD69vVkMTKYFYDBe282LMYsU3BwOCTW+taxUfRlMxgdGhTQx8aBbNWJ7dtx9doNHD5xGq1gFMFIQs3rI498GL/5m7+JbZMTqJXW8NLzP8TJI2+gVFgTaHJzfhk3ZheRL1T1/bRD4HrhgPD2ndsEVPRnMxgc6Meps2fA8PZ8qaJBS2GdNmch9HZnMDw0gL5cTsPOL/zjfwrEM5ieW8Lpk8fw+MMfRN/gCMqNAA4ffgO9uazUBcePHkF3No3JLVu0f9XoN5xK4cLZizh/5hw+/4UvolJr4sr1KfzFn/4HfOM//Lmz3PDi2Y1T1v6kxURtG+gA6ErEsHNyAnu2jEm1QZ9d+vWvLS8rK4Xs8miI62gIYyOj6M31qrkjOKkhWwBYXF9FMxxEo9pEfr2M05eu4ztPPYXTl65Y+Kb2zY29x55RstyiYmj/zj/7bXzkIx9GKhHXQFXNaXDjjNtcJ/AzrJVKePoHz2N+fhGPP/5B7N69FdxGw8G4BkOxmIGRm5nb/HcXLl7DzZuz+KOvfQ3nz5/veOoS9PKKCg2lHPDurTH4d7QV4uel9YFnFWq/5dBpuN9UFcur6BsYxBee/KKyWYYGBzDenwVPpdlrV7Fw4wYa1aKG0GROLy6u4OLUNA6+cggnz59HqiuNfXv3Khvm1LkLOHfpivZqKioGBwcF5LDRjkXa2LVrEl/96q+jK53DwMiYhj/FchVnz5zF1q2Tum9qDKVr9i0Nh8GM/q4LqDh/fgalclD2BdOz13Dgrv2IRE31GWzHUCzQ/mwFq+vTuHLhHXz0kz+HQpPZMN2orzN7IIa55WWs5ZcFQuzcuRPrq3kpBQhYxKNx590cxPT0Nbz8k+e1pyQiLfRk4qiVCygVaP0UlyKGOQ6sMQj+0Iasu7cLvQND+OCjj+PBRx7H3MKSnnmCdtvGJ3Dsnbdxc/o6GtWqbJUefuRRZHN9aAQislsiY5F5Gdembuq+HzlyFM889V3Mz10Tk1bB0mKfhtCd4fkSRl9vVs3h6lpeChxmyMzOzltGRoT5KkY28eeMBuLs/cImqdeQQYGKbJjMR5qqPbPSCWJ0bBwfuP9+7Nt/N7LZHGrVAL7/d3+Pt946hGJhFaXKWoelzUbW2K/GhvVsUGPQkZxi544Yew7IsGeHg/4ghoaHxM7mYIN2Nfxvrs9yvYl6taYhLDN5aPu0trKMY4cPY2XhhrKE7rrnfjz4oY9gfnENxXINoSDJIbS6iuPQobfxgx88qwFIncMoDnQaVTQcg9aD81brWkYJzz2/DL3FQ8fSpe3BGGNNW5gu2cmsMy28mf/GK5501nIg0G5LfcfndEMBbM+vz37jeWcMWqoqaJ/AoHp6hNvQhN/rQ0blxc46OWb1CAkcvT057N+/Dz09WQFblQrtRlto1cnKZjAmQSRj1SucW8zABpZXFgW88d9xv+TxbACtfdl7tNpbSuVWWxlWtH5KJuMdoCIai2hozYGjB1MNVGGGBIdEfJ8RZR8wV4sghUJJxa5tyl6ICinu+6x5GKhOUJGMdt6/5YtL2m9ZU4gUZDPOjdDnDWzBDQtskM+1bISpDRslY2nbs6GhQTCAWNT8+HkPWIOyHhWBRXUh61AbxPvajGqLjWtk2QpeNW5EKl5/G0j4Gp3fb6ptUx+Zgpr7tVklyY/dWZH4PokHF9nu7L1MocDBr32fCEYilzUFYprNBoe1tK6xzx9h39OoaN0nE2FkejK4duGKVDccCtIik0pI5gVl+3pERlteWkUoGMXswgLGt24ROMuaqljggJvM4gBW1tcEJgp8I0HNZ0DU+JnNPsiAf7NM8kMYT7ryKhLaFWkY5vz9vSURr5UUBQLeae9XFnilYaCsv2DWPg6I8BYl3ra3M1zk+lPRaFmDBG34PPCZfPngSxgZHEK5ZMAa7wf96BPZLM5fvqx8KyVdqA+2volDbP57y9EysxA+9ySEECCTpz1Dd2VzZLkSXEckc7FveuSRhzWo577HuplZFcwJ4GsFCZIxD0N9G7NmAiiV1hHnmqyU9HyG4lFU+Tw7dVqMDOZyRcCfGO3sZWjTW63KDpM9AS2Jjx45bgN+kvNSXWLSZ7sz+jckKrGvM6GJDQYLxZLLFyF73gBb9mfaB4J+ZkBPeevRtM6l/jEmta9N/HlgQ3unpnH9FtcOB9gcaqrnWs/LOk3Pp3d7CBgBg7MI7rM6Z7gmSBijxSNV6m7f8etI/a6zz/UgvbdY8o4M7D2ohuS65s+zmYZXLDlyJQfu8iKy33xGpPfR157swEifOeBVaAIYw6ZYpDJJ9REH4S4nQwRPAeJUr8acTVVUoARrIn4f91HW5uLrOIBCswSuY4JYpZJqw1q9jEQkgFCzgrH+HIpL80hEI7h+bQ4DQ4MoVGuqL4rFdfT3ZtHXkzaVZpifiYP+NkbHJrC8vI5Ko42FpbxyvuZX1lFrtlGqNrQ2RSKjIoHzCqGj9kyxn6xV7DlmfRkgMIc2tm7bZvucU7xI2eMUAwYiEbDYsEy062kApZ+BiAzkACF/nnhHAl4TsfcdaKRplrNls3kSgWw3fOeipcKoZYAy9yfNY7zFl7OB4j2W84RTytn32b5r78vsK62XN9szD5r4WZifRf2DuaGrc410Sbs0yypRj+Pmc3bGkvxheQ4C0Zy6gs4i9p5NJeCZ9n59+rzSzkyoE85sqlFPirCenD/Hs/7NVsirgjTz6oSLm+rJz870Pgnecf7mVFD6d5od2HkrSzqXi2Qfz+wOvaLDAyLvVlR4dZcHN/ianZkM662fAgD5nNp3X28Cux6okDOL8nNMFav6SipGWqJuABOqeTirdMCEiBGOeCZgSYC11X++TvLrzwMg/h+4beOWtyVS8Sa7dVlWRez6ahb6ri9TVBj5R33i+0DFz+o4/v33/dOuAK2fDIG2gE0PVAildX5uLJr550L75RtqzZf3xOPmxwecTB6Tr8fdw+/yJySl8ywCKyw924WHjv7bZTF45oIvWr1kU8WDvGFd6r2z2lGxShZew4p+a7bJYjFpHRFQbWp6/y58Rs2PobGbvfdVpPEQ9BLCqsk9jSFfVMEiGWjVEGzPDrEG3AKAWQBJqspNzIV4e2aawqQc48oYRCxOTAruw3jMA9AaXPP8tSGsyVlNVWEBhvblrwvfu2eP6M8pW2MBTuaHk9vRholMbb62VBRsYHQOW9AaCyfJRcVs9L6Lxl7hZ+T3aCMUmLHhJWshy+aNydev1CzUlbY6kszSoKNJb1RTWDzxxS/eClQ4my0xQaomCWRTx0EJizEOetVAuOLShm2W18HPyd/phcwimZcr193tZO7A+soqDr36KtaWVjpABRUV4XgU23duU0E9NNCHEhUVmSwSyZSKRkrYCVSQuEQJtBUClqni81pW11bkBSqViztYWNDzPpBlXCqTRVzFxeNHcPnIUfSluxCg4ibBAX0EaVrSJNNOpcNi2yzV2AD4AYgvHPwwievOGt4NKbtYHLQNiXchke5SQVColDTAIUBz4dw5ZLuS8hnu6e1FKpO1QYcbMnDI6plNPJg5LOAqUHMhmyyzrvDDFT/c4iG8srKASxcvItfTh9179oihruKBz1HLrA1oJ8E1xCFXJBxHMpnBrr13KiOAQI1AtXcBFRxI8DPzPSwtLelnMwycN8wCtU2SbcxV94wI4rMCgY0ymz6yqIulFTzz9PeRiDaRzeQwNjqBXK5HA1b+KlcK2DK+FUODg4jEYlhYXsGFq9PIVxtYWF7DKwdfwkcefQT7D9yLTC6HGOXzLETDYQ0B11dXcezt1/E2PdJvTqFSLuh9EaiIRRNS60ja7Owy2NHGokGMDWe1X3BtkbnIwSWbMIEWkRDtYTExNITB3h5MjA6bxVBXEtenpzA6uQ0LSyt49dBhVJoMsw9IifCxj3wMv/xL/xP23bkPyUQcC/M3cOb4YRw5fEgsY1rAzM4vY2W1ZM0Rn12qntDG3h1bMdbfh950SkOti5cvIZpM6nqwPmrUq2qsBnpzGOjvQyQc0DPzwEc/gUCiG+cuXcP66jI+9/OfQk/fMFbLDZw+eRTdmS7s3LEDh99+C1naSk3QJoxemmENmK5evo5Tx0/i53/hCxokvnn4Hfzr/+uPcejHr3SKxnefX74wpKqCAyXth7zmsQgmh3qxa/tWqSYYfkv7g1q5DLJyKWlnE05VxejwEPp7+xTwzLVMZjaiITQZtpgvY32tjLdPnsV/ffY5zC4tm4etKwb5jPuBlK3TsIY5/8f//s+xd+9uDbWHR4Y1SOA+65+ZzZ+DS3e5UMCPnjmIhYVFPPzwfdi9e5vUY9Ewfcx51pq9oLyoXTNAu4+DL72itfcHf/AHHVY6QQoCDtwfbpG109IsTv9pWkNZICdfiwx1Pl++4SWTjCw8qiFpL0HA4LHHH8enP/1ZjE+MIxGPIpfOIEu7qEpZKiIqggi2zU1dx8nTZ/C9Z57BxatX0d/fjw/edy9GBgdwZWoax0+fk1IjEgoLqMh0ce9jKHcEA305/OpXv4rJrdswPDaOgJi+LVyfmkI4GFYmwWbp9MbZx2aX2UdBARXFUgAz8/O4fuMK9u/bh2jM8gRCgS6Uiw0Ui2solBZw5cIx3H73XQh3daMr0Yt6sY5IMKoMFwIVtPHiel1dXpOyrsrBFM/+ehVXL53F9773Nzhx+ihqlTzikQAmRgZlr0GrLuZ8cMDDwS4HZ1Tt8AxMJYNId/dictdefP7JryDXN4CF+TntcSOjW7F1YlxAIEODyVAlT4tgTZkhpC67iOuT+/TC/BKeeeopHDz4LErlFQQINrRbSESjSCUTGvBmMkn09eVUk9HGkGfetWvTsuLwQ2HfIG5exzzba20LhLTaw3nau7UXky2I+fXSOo4Dz3377sQjjzyKy5eu4cWDL6NULKBYWpMFFJVtrC+8h7QadUnp3fnicsWcAN4J4R1oIWuboEDArZNbZBNBkJFDG9rnjY+NodG2rAC9JofnbOybLczevIFjx97C8NgEPveLX0YDIaysrKu+4FA6GjHA5ZVX38Czz74I2gfJ7ifAYOkqaMXk7YA845JnrgZnlZKGj95bWc+/8zC2z2pnE1Umqpeo4WD+h8sLUG3kwu55D0RECFhgtM55Dfzta6P+c1Y9sjywsHVrUANosh58V0C3NdNBKZSSCYZS05ougsHBXtx94Hap4lrtEMpl7o0crLIQtLwdyLjDlBusa1dWF8WophpOGUsM4HZKMmMHWnPuSULcXwhU5PPrSKUStwIVUrqaosKzYc1mgQxcy0MoFstYX1nRgIc1oKmrmw7Mt72UKiu+H9Z9/Jw8t1cuLRvpJsrPasHTUh5LYcGBKe28DBjiMyCFuFiZ7mLrf5tNH/dCX+d2iDluQGR2rFabcIjQCSx2uRN+r2INYHZYpjC1PsCy1ThA55cUHQo3NsY0fxeLk+/B2RvJXz9KZqcRi8T2diGveg03vOC1kjrSMc35uhpkNQl60ErVWP7cAzQ8FljC0GYI4CPYmklFEYmFcOncRYSDZgFEkJ9ErWwug56+Xu2LtHkJhxKYXVxEd09O+wTPVdr80FaK16hYriCdTQuk4C+lHHDt00ovnlBNaN77BsLwZ9m5ZatfQxmF1xthjkAVh648Q2QjpGurItbAPToBhEkeYa4hiVXeYskC5u2aG7uaP4NntgAC9mpuAMq9s82iv9VEfm0dJ44dQyqRkiKDQfQMClZ/GQpidnFJNlBcz9wHFeLqbZ0c2UfZJlTdsw52FigEUbQm3ZBNfSrJEQ4ofPiRh40NX6+J2MGzlkNjKcx47/j+9PkIqBDAoLUTwWojvJVrFWVRaC03W0jGkgLaC+sEDlNizie6aHXZwkB/L3K5Xl3/V37yKi6cv4juXA4Tk5PqtzmMpfqV153OAlyHBANMrW9kOp1XzgKYe6UClasVDSqVzyBnAHNQsL3CyI3KHHADdg8S6u/DpnLogHSuv7LAaq4z1kaWw2WEPLMU8/70fG8EBzxrm/9tmS1UYVgeBfs0rgev6OPa499z7/LZeN6VgeuUP9cPxE3Vag4Jsn9z2TV8zqUEcP75HXKJG7wrSJsEAOdA4TMRTGXXUv+9kffhLWFsbuJzIvkepNBww1096+zbHaCq3pQDzSZJYgYu2TWuI5uKoV5cxbaxQdTza8pxpLI+ke4WGensuQsYGepHNk2lK9CslVAtFQVMVqp1jG+ZxHq+omyWtXwF1VZQdqghks3YbzGrQYoeqGfUYJvDZ85b+NxXTCWh+0FlG1rYMjmpflqB7wI4bRbkr50Nu22mw+veyeHkdaA9NPMTNedgXWGMfk/g5Jpdz+e1Xvl9VJfQ0pgkPbOu9vkBtFDcyAEQscgHUxsrtwMm857zPXEPkgJD1ntGMNUQnfutU9Z5dQ33cwXUu/WuNcucpPf6cqAInw+etfxdg3in/tG1c8RTr/jww24Bba6XsaG1k5nI4WADQPfXh+/Pg4R+zduczIAuOX9QbeTWlA8d32xHqz58k8OJJ5n4+ZFjNRsI7cAk74LCjV3X0uefekWCz9tqtXBqk/XTHZ9gH2pgkAEmNrTnNVHt8dNkE/4yvMf15pmk/UJ7mM8ZcdfKKRQMRHY28Sqs7Mzle/CgBE92fy21n7v5jNUSXD/2w2WL7eatm9+OwTgOkHK5uVKgOECOP8fPNN/9MTQCEcHT9oz3gYr3frTe/9Of4SuwnZvEJljPgq7MP9IYjIZ2cpPloNp+J8uHw+mGBrLeU5CFi4qIZsP9mQ3gGy3nHefCZowNsYHeSrXhmGN+IG/BXiYR0+CF8in5vLpihxuqJO+GqHpmEpsbbqzmz2gPsN+Ytak56Z0KEwX6NVQcdGe7dcixeOHrcdM3yyYXkOMKFWsyCZjYJs/rkM1mNHAkS4b/xsK2bZCsGsUNVH3YDt8zCxoWyrQ04GuSdUnQRKzfCL1OjeFASw5vzWAWGGQLmXKCAyvPxvHDe8qpuYmaF6LJJFmYcR+r1Kudxo6sNRbPyXjSVB3M+yAjkcw/11I1dYiEFcLMAp2Sb34pcE4eu5Z5YUi6NXZ8Lfo/kxFQLOU1pCOIQZBCYEaghY89eauigoWGZ/aWKywmOQyodgLUWWDwQnJN8HX5s8XyccNC/p7NplGuMvAugO5sRoMb/uyVxWW8+dprWFu+FaiIxGPYuXuHGtL+/l6ts3SGwaMEPFic1xSKymEDFRVaO50sFWuoCFRk0ukNZQsDdqVuMCZPrUmgpoBmfhXn3nwLwWZd9jKBKItekzezceD95tqOx5NOdm1r0A5POxD55ZUVnsmhwYkDefjvY7EUuvjZ2Yi3WigWCsqooKKiJ5cRUMGmJJVJy8vZB1GRXUqQhMMA/iw9QwoaZB5JGEGFrZqigp/bD125rmqVEqamrmM9X8TuPXvR22d2Nyz8CFSwASOjzxhkfGb5fMYxsW0XevsG9BzxCTGFjykq/HDLNwccvvIzM4SXSFS1RvYnC0NTgG0GKjTAFjmOxT+DpwuoN8p44fmnUVybU57I0NAIhoct86FQ5DO2ipGBEYyPjStDhKqU81emMTW/hJX1Al598SV89EOP4c79B5Dt7UGITCv6aBcKmLo+hdkb13H87Tdx5eJZNbjcw+oCS/h5gwoz5F6kwReBSv6fGoegwCoOXHhtmcXhWSoEDximPTLQh9GBfkyOWZg2B3TnL1/AyORWFEpV/OS1tzC/vI5YMo35pWXcc9dd+MIvPIn9992vjICp6avIpGK4eOYE3jr0E0xfn8Li0rrCtAnOMVSeP4vbJdUIE4P96M2mkU13abDcCtH3f1nDTrJwqZChVRqZrGyMeR1zwyNoJ7JIdfeLifzgA/cj29uPhfUK5mamFNC3detWvHnodT2nzL+QryoZ9fEErl6+hhPHTuDTn/0cllbW8Tff/S6+/q/+BAs3Z51C7FZFBe+xxcPZL2MNOWYvbaDCwHB/D3bv2qG9gPYftEbQydFqGpM/GkUuk0Uum5EFBbFXAgSBeATFJplqdeTzNRw+dQ5vnDyFm3PzKNLOYNN5YOC9Dde4/3/840/gf/kn/wS5XDdi4RCGh4f07sIR7/l6q3+qByqe/9HLmJtdwIMPHsAdt+/UuolFkgpAFFPGKe14vnJ/4zDkhRd/jB899wKee+65jkUcwS6uIbEm3Z7hh9Bs2vjFs0vy6ZCFSXrGsFjetDaMhmVlx6wdAlk7duzCl77yFdx2226EafsSDCIRiaOLVlnVitRn/IzxZg0XL13EH/6Lf4F3jh1VYPonPvI4cukunD5/QbZZJ0+exPrqmlQEXOe0LEglGEIev1C+MAAAIABJREFUxm17d2P37r244867MDqxRWuXgGS9WkcmkxarT+eSmktf1AfRDNhQ//yFWZQKAcwsLuDytQu48/bbkUrHzGc2wAFaXQq3UmUF1eKS7JQakQSS0TTatRbCgTDmVxaxViBQkZDFBz3XuS8y54hs1sOv/wQ/+uH3MD19FfUmB60VeX+PDQ6q6W+36NUd1sCO4ehra+vo7s7J0zidCiEaTyGZ7cMHHv4QPvDgI7LD4DAhEs8K8FtZnJN/O0FyVV8EKNweJ0UMWfcrqzh+4gS+861v4/z5U8rh4HCe5x3Bn0xXSoBFT1+3WPS0Yqk321haXnPKCjKbaZnmrGHckNMD4hqaOFWl2VWY9RN/5wCS2Q+W+2FBnhzY8O97+vpRrlawtp63ukqNuQXBsmbRL3qPO1a0zhWuZdfI+TBtG/JbzWUe/LTciUlZQ1UWwWSuTZ4x/N/xeEq1gikqjAXIfZZ13KXrl7HnjjsxOrFDyjfeD6lXg2wkuRcE8PKPX8WLL/7EhrYa9nOPrgjUlLRf6gcywM3Pnz+XDHM/5PYWnL7ZlpJUta1jauocMKa1rBoU9GvWjt7TWudcgArNgmuWbYghFYcbatnQ3Opkgnfyeee1YzPtlDAEMKxkt2vAgQnB4Hg0iVTSwIpEKiIw9I479qDV5PC3glq1hXaDHuJUvFJxy33HwBDWR6vrKxrU5nIZ1QYc5HobCg/cGlBhJBezfppBsbAu0HOz9RPreIIEHL7LE9yBqH4tsQbnQJoZQVGGkHMwmUwJJGctzL2Wg3cOS8j2TnUlTNnAjIpLS2YF5MA0Do85MGAQbJiKaBHf7ZpyPzGClgtKdz2JV/YKcHI2tD6TzbMsZZvp2PBm/2LDCNr0mTrbrr+RsWywKGsr5yclYMYRtLi2aBfKGteUuGUNSm2fM7UzrYx4XhmIAvVcnsHKGt8ITFYrqh5yOReWj2G+48qnoxpeYaQGRPkBDDNZ0qk4Qq06gm2GMrdV+7IuJSO7kF/XZxseGUKiuxuzUzewslLA2PhWnDp9FtEEyRjMW2tKlUyQmdeM73vrju1iWKv+o5WWrDRs/fP68Oxl38N62QhYjqnq9wAPXjifde79vFYc3pqixT4Ha10DV83WhHuCai6eTfT7bxLoKqK312xeZdfrFOFUEwSdxQeJBRxm0v6pkM/jtVdeVUaFXk8ErrDeb4lKew7gSbrToEg2/I6R7M55Pfs8W4J67mtNqsptP+B+IXWGck4MYGDvxOft4UceUX0llUipoIwK/m+eK8wRiMQZMG/rl4qLbFcC7WYdE2PDUvKSKKb+q1jCjembqFfIEI+jkC+KPMNcsFqzAWbM9fX14sCBe3TN3nzzLZw5fVZ5BFsmt6q6euutt5FIxkUSo1I92eWC4OUnbzWEKbZsfTZadQ3HaRHGLwImiVTabL2ccsj3pz5cl3sv17yFL5O0s6Y+iteIg2btsY58x2eXdTfXOX82v4e2dFSzKjS7UtF1IvBi2S28hiVks90dVUWtbrZR7CuoYODzJNDLAx4EHAQc2h5ueY8bVrSybCHgKa99A1R4W7mm+eyRzKPP5tnPbn7i90wLnDa7Ve4L+lnuNWQN664Tr5nsvlz4Nu9Rfn1doBF/ebDX72G+RtBeoPdLG8qmOUJQ4VLNI9cVQ6ucR4L/u0znA6ohmkimc5ibnxeQPTY0gEathFQ8JDV0MBhBIp1BrCuD+elZLK0WUKw0sV6uSqHN36uU+LjZDK2fSLQSyU3XI4JKoejU0XYuUV0VicexY9dOncusn/mcqXZVNo/ZWOtXu6VnTnbkJBy5fc7v3wZ0Wg4Qrzu//xZQic2s1EX0UnDuEE4ZzT2K+zL7Vf0bZ9vHtcH/lkUfSZMCvxqmeNFMheQod6+kFnDOFS47gWtGgDNJQbSCohuBc8fw58p7jQ074JY7lzRDcgpTm7NYjy5Cg8tM5f0VgML5hKuNBUj7wb17Lf48DfidfRI/t7de8rM0U7iZC4ifM/n1ZXudA5LYjYrsalbi/stnORg5y0AAX7PzPRvoYrXnhsXRRt3i1SH+GdisqLjj4yu6B7KjYp3qABuvNtGspEMOfq+r+w//zAb8VgN40MGGdgZQ+ffr1XSaA2kGYvfBA84dJMKpFHlduA/Ydr8pONwHaftr5lVhnZ7GQA5TcXqlir1v++z/8IvnqqkwTLn3PlDx33fv3/+un6ErMOGT6t3B4DdKblJe/mXsMGNEsFHhBiUUn4xYt0HyQbVhox3YkkvJB48oum0EfoPV71Q3SKJrqKGXsvHhZIAND/DN/rEWNGVMah70Fmq1EfbtDy3zU7ZN0BR4hrz6psGH5Uka74evboCoUNtNXneS4TsLJPM59BYFxq4gi0jD25Y1yNZEmYLBX0e7JtbYm5Wt8eD4xebBfjfGnf8+Mo6M9WrybZ/VwfcuBFrsPXod2mHkPyu/XwCCa1QU7MnMARZ99F1tcADPwRL088REoGc5vaK5Odas6JLkPWDyXfbHJns1iTqLKxYLbJA42OJ95HvU+pDPah0N+jQTIGJ4Jos8l1dhh3kDTzz5RXd/LVSTRabCCes1ASICfegDqcFaHZVyWdfPmBN8zYb+jGwsn8PR3Z0VUMGJUk9vjwEVQWB1YRmHXntVyoodO2/D8OgE2hw6xGLYvXe33l9ff07vn0NsMqQIllSqNaytr6PVpJ0ZwRuqdpyiwh0k64VVyaa1BjjgD0cUxheLhVHSa5TRapSxcvMa5i5eRLPCgMG2vGr54dh8clDLAoz3ksW0ihH3rPjr6sEBP7Rgo2VDUrMEk5ycxX48YQW5Y6DQZ/f0qVO4fOGChssjY8MCKrqyWWM1OQ9fZb94qwuxUmIIs1kjE47NfpwydCtqvKqE19ZUQ8xZWMPlK1cwOjqGbdt2aADHwo+DXzVqKtRqYqwHAvbc9A2MY+fO3Wp2FDnoKAc+xHLjeWZxQwZmWZYoKkqdr623wiBQYU+UPVscTBjLhWulJtnzkcNv4tKZd9Cd7UJfbw9GRsfFussX17G6voTe7hy2bt2OVFcGCEdx/uo0LlybxlqxjFeefwEf//Dj2LvvTmRyWQ2KeQ+oJDn43I9w6fw55FeWJNGXRZuurUZNJv/XZWDxHNEAT4MNAhHRgHzphwd6kct0YXl5UbYXfBbyZGdHY+jNZjAy0I+tW7aIOUfW/smzpzE0Pi6v2LfeOYETZy8i29OPQrmKXCaDz3zqM3j0wx+RYoXPJwcUaNVx/MghvPnaK5iZuom5mwu6jjUCr21Tg20bH8HEUL/CtMm4XaA9TbWOxRXauJQRi0TUMCfjMSRiEUQjAWVPBJMpHD11EcmuPuy/+x488MAHMDA6onBiNonxVBwDQ0N48/XX0ZftxuTWSYGm8ZQBBtevTuHw4SP4whe+iLPnL+Hffv3f4fv/9XuoFkudPdEX2XZVTTmj5sP9gbB2nmXM4QlSIRbFru2TuPfuu2UVw5wKDtmTkbCGuSE0Zc/ENc6GSoOGRguBSAB1Zl+E4rgxu4rjFy5gPr+u8GI2/bw/skNz+T22/wBbJkbx27/9O3jg/gd1TiViYQwN9cobmE2bBaNaQe+bCa6j1VIZLzz3Cm5Oz+ID9+/H/rtuc8M2grK08+Czw8bTlGP8hMzOef65F/Hnf/GfcPPmTYHbHPrNzMyI+Szm3iZ7RQ9mShXmAFDuHWx2rSEwoEfFbrOJ3t4+jIwMa/8jMPalL30Zd99zLwLxlNkrROICGTicIpjBPTkTC4N78J//x/+EP/5X/xJjI8P45S9/AaX8Ko6ePK1njcDX5YuXFKzerNX1/ckEz2EXXthoYGh4BHtvvx0ffPCD2q97e3r03FgDssGAoz0AQW+xdBHBhUszyBdbmJlfwuUrF3HH7buR6U6r6Q0F4ygWqyID0AquWs4reyXFjJJokgbL2ksXlqmoWEEyEcOunbdhaWFRYeBT167iJz9+CW+89hKWF2/oDKOPv8B55pPEEwoWp1qH+2R3Nqv9YWV5WaAP965kKoxYPIlwLIFszwDuue9+bN++Qx7ewWhKCq/Z2Zvo6+9HNJpAQLkGUduD2XS2oLyl2Zs38cILz+H73/uuMnb4PkJs5MNh9Pf2KFg+k0ohm8uiXK9qOJAvFgVUcE8S61GeOI7RZ0wKa9Bd80S/dZ0vYjpyaErShdVVYu86hRBfT4x6t3eTUykSAQNV+Sw55aU8fgVUmK2IDfdtoG1NoZFKNJDxBBmngGVdks4kpcKiqmdoYEB2WjwfJsYn0Nc/IJIB91VT5vkgzDpakTCGR8fRaHJQ2pBtCO9XRH0xF3wATz/zI7x+6A2re1jLEKioV9F2oDxrXdV3XPcMjydYlF/vWEl4go1UEJ6hKdDUgQ062yxboh20oQXXMptOT0LgXiYLl2JR+6X5sPtcKp5t1jg7u3ZEI2ZF6a+96kZtLOZprPvIXDAXtE1SAusLqm1S6QR6+rI4cPd+9Pb0a53yvGR+UpNK1QYHfNw/TInAz7uytqRhUk8ui0jIQkO9JYmRcbxtl511rHNvzsxgPb8mZjh96/mLNpsWpu3WibM4EXNaIkjL1mD48erystlPhqMaSFIty8ExGe9UaPJ6pzNdSHYlkIgzFyyGhYsz2pusLoo5RYKFj1v6mQ04bAi24bXth2Ja3w6kMwtKY0AK/HJBuuxZvAWdkarsHOL/57r31qm8H2ZPsQE28RmSYqlqjGgNc1xOCwfWVBmwDvMKDtZXzFzwbHGvo+br2hBMpkMapHn2t1jdjYZqY2Ne2z1hLU51oYarGjgZ4K3XaVSBZhWJcBBdyQhQK2NubkHriCAR/22lUjQLPg1LiyhXWYuM4MbNeaxyX5qbw8TEFtyYmUVXOq0cHNo6joyNIppgnc5BfV31SChg6lzPDheD11nz8jqzD1FovDJjbPjPdeOV87Lq8gxrx3S1LA7mNVQss61WU73Iwa7qUefvbn0MWflJDXo7wE7HRqohoILnC/fvk8dPahAvBYr6UiPqcC7L2omgLJWHZrHr7E0aLudESC3VGVQLBbTvcnjMGpr9hR+smuKdbHSqOht45JGHtOb5+FGdRhVquVBU/c0zhAoFKe5ZVzTqSMUjOmdp90nFbatZ1YIUcFBjfV7EpfNXEQwyZNtyLPicEUDi9eD14hrToIuD/TItJ239KN9EfaoN7JlPwfdG0DCZSOlzqM8n+Fgpo6evx9QjytgLokYiYNzlsXRsBunhb88Aexd+P9ew1jnnAQ6cNcupmCyDzMHALEp5b/mseEIkg8f9F/d43xPxPm+2W/PqJV5HnztgrHLLh/Bnhw9ttueQuY22fsToJ0AWi2qNeotb7cubyGR8hnWfHRjnySIafLqsBLOq9meGKXG8TbOfCZiK1gbQJNfIxowWhe69iGTSaMhBgFkaBAEF/mqIbQNu3yfy3kWDDaITqK2vIFCvqvfgfUtmerBI9WiNSoEABnozaDUqiEeDqoWoqBgYGkZPb7/qK9rG5st1FCp11ANhVJotC9RumpJDFm8up1OgvavNeTDI4rjZkM0iVT1jVMu6YTzt0gTA8vWcrZIpnqx2sD1zIxPJW3WLWOv2RAIMnsBIQCvDWqxqz7nmJrKRtmG97dtBy3RUxqjNOdi2+vWv9++s4Hg/pXhxe44sefiaZv7miKkbA2/eT0+o7IDc3trSk24Ectt+Yd/j6qNN6gN/fWxuZmtGqh635tjHSenoFD1G6DWVmsgODpTl5/UqDwMOjXzBr82KAQ8gduyKNEvZIBPz5/j9m7/7HAuBSi5DT8+OAzKs3zUFY+fLWdJqtrHp3/hawsi9bZx8lmo9+/KKCv/5PeByKwBkdld6vwI3rbfxQ3x+r7/G1ovZGa9nTlZd9hm4VngNScaSVby7LwrS3jTfExjurIel7NsECvE1/c/V9RaJwLmjOBWEr7H0GqqlaDdl79ln/3olyy0kLX9RXO1nszWbBb4PVGxaZ+//5/8YV2DLLbvHuz6T+iNjMHYGh7ReqdU7vvz+MLej1pobfzja5kYLoJrzFXQTWscO7zRqISsS/CbhCzhJ6Tik8JuLY9z4IUynAHASWpOrWbPrh/s6itzGYuCCNQfa2Mn4qBq7wrORvOWO9671KLB8OSm3bhhTQZu5pNj087TgLxuimwrBh3/z8CarkZueDbspUXU+zAq3dl7DThKm73OINhsbHQS0I3Dhxj5umge3pKcqJg08cmJR19Ra0SlwQc1dU++NzQKVMULhnZpGiL0Dkf31EoOS8vcA2YAuWdB25Y4sUh2pU9zwmiujghtshJ+TCgugUMzr/otN6ayfPvnkl6Us8I0WGwkO2hUSVrEi2bP3BVQokN2ulS/+2NQnyUYlIBYIil1HJhEZqZSns0EgWLG2uILXX3kFxXwe23bswtDIqBriSCyOPXv2qpDuG8zq/Wa6DKigZJ1MoJW1NaDFhoBsIcuo4HXkOuJ7KleLCiilrz7XB+1eyGiKx0IoVjkYKwK1Ei6dOoLq2gra9PyUdRmzLM2CQPZKjhnBBkDMC4aGOaDPI/2637JpoVczrYXsmWQxwfuvQUs0ogwG/hnvHwdkJ44dx4Xz5zE6NIDhUcuoSBOoIFvS2aexWSBzS8PKpnmbys5Nao2o7CP4XFGBoHB0B7KZL6cBk1evXtV7uv3229XIsCBnUUm2vuXE0HbGQDQukky6D/v2HUAkFLdBsapGSvAJfnSwPPezQgrnY3Pi7czEnOHyk6LCAaFuCOwLD7Mkq6sJmrp+BYdeehY93VHZooyOjCOV7sV6uYC1ItmbwI5tuzREDEVTuHR9RrkE+XIVrz/3HD72+KPYfccd6OrO6qfM3pjB3/6X/4KT7xxGg2xBN6wxZpnZd+jPHENKRZGXE6swtCFdBA30ZeLYuWVUA7Sp6Rtm+xC04rUrkcDQQD+2b90qNcCW8XEcOfkO+obo5Z/CqXOXcPDVN9DTN8RUD1nx3L3/bvzyr/wK+geGtFdnczmBgbXKKn74g+/ixJtvobJeQKlYQalRR0XZMm1sHR/B+EAvejMpDTsXFlewWqzq92qT/tVJdJFhVGbeQ5fsIkbHh9EOhzE1tYBLl2cRS3bjnvvvx0ee+DDiKSpPysgNDqB3aADvvPEW+jLduG33bVjSECuhdUY1wWuvvY4nn/wynn/uBXzta/8SZ06dVqgZr5FG1L4AVFGp0vi9D2CG+AWbYjFm0l144N778LnPfFYhzqdPnlTYeReH42igK0Ew3UvWyVSOIZ4Mi/nYDiVw9eYSjl+6hHa0jUgshWtXb+Dy5Ss2MBQrkqAkfdTruOfuffjd3/197Ni223yBY0EMjmQRDppFWIft6opXv+GulKt46cVDmL4+i/sO7MPdd+3WHhEMhFFt0nKDTb8NJuS13A7i4qUr+MZ//AYOHjyIXbtuw9DQIL73ve+J9UwQWYW0awq45jy7zBf4JA94JvPmQSMvKBtJ2jaRrc49jv/mU5/6FB599DG0wmRWxpDr7tVAlECFwAOBkcaoXpxfwh/8/u+JofuFX/wM3n7rdVy+ch2JONfTIq5eviL1IvdjDr7oe66jsQ2FcVIVQobxrp07FeZ9730HcOedd2o4bfuCryG0o6BFUBARXLx6E6v5OmbnV3R99t1xm4Bn3ideQ3qMc3jGc6NcLYklSrUDrdnkJx0KY2lpGStrKxps7dl1GxZn57CyMI///I0/x9tvv4ZKeVWqCVMIbABP2g8DUNA2gTwq9Fg13bxxA9lM2uwKIkF9Lu4L0UhCgMT2bTswNDSMXP+AMh441hwZm0AoTOA+IcBYdpVkRVbrKOQLmLp2Dd/85l/g8NuHBBJzE0wyFL07q/MuFY9LDUUrnFKNqsYy5hcXpfCiNzktoDjEplLQf4lFpyGteQfz/fI8lpJTNYTZP7lHzxQ8qgmtqdbWzTXXqAmcV5Cknlv7GcaMNCaxakPXEJoFiw3UmAXlrVr0ei7slYq8VCaB8bFR5VOMDA2hO9Ot83qgv1/WEXxjVIf5gGv+PA4UewZHkUx2aZjDgGbee6kbWJe26B8fwnf+5q9x7MRxUzxwwEbwi2oK1idOTcEzj+87Ho/os/FnecsQP6jWGnCMTNuh7JxXvhgtUrh/iVHuFKjO/tTIKZYxwqHn6sqqVE0cKivcUeCJlXZUtKhWCBl7WYMEu8BOIUDSi2VY6H1x6B4xFYfeEQf4sYgsXGindted+zTQbniQgoCoAmwNeLAbG8AyLd7W87IDNBYmFVumRvD7sgE2G4P7mdlZKU43gAqqHswGRjYnAjiN/OQDKlsgGMQMgAqWl5Zk+8T3l+5Ko0CbxkIByXhc656kmBTDvbuSiEe4h4SxfGVWa5b7JW16uA44kOS+YaoCCwrluSoLMHcvzFJpwwOc9bAAM2XW2ec01jtz3BiYGu2QaHivZdHKoaxj9XId2nUy73CuVdYFBl6ZIttd2s7Qw+p3U83yS6xhDpLckIk/h8MTY4pbTb6RR7dhpcbvUdYceyoNi4zgResmqvzMpoc+7GZpy9vMM6pWLiIWArJdMQSbNczNzsv6lOH1kS4OsqlQaGt9LK2sodGg7WMv8gXWwTVcvnoNQ8PDmJ2b195DWIgh1cOjI9pr+X51noQCiEWYJ0fSi1n5qt/zzFLVSLcyoj2YYONyUzZrPbveVL7rjghg95Eh1FSqWIadWaLErSbdNCj0Z58xUn1OiAKlpKiYmbmJc2fPi6EvkDMQUgad1COBgNSE7Hq5Lrwli4Ai2lj5eydbEgOLVAs7hZpY2s7yxNeGLGW5fz78kAMqAlQ3hwQAGFxJ0hTzNNx/C/Rpo1ktoVkvi+zC4G2qh6i+J2kqEIxiZbmImzNLAHOvOExmXkCNP9/IRyL30W5E+53ZaHJAbuon6wG1H0eYmWEAi9X+DAm28GrlEzAwWEQtDtNrZqusvEGCrwas8XffM3jrHGsrLVfFLHTMCYHvi/U717QnTfrBJi1uNJQPmx21v5f6Oa4v6WQwOlVTR63AfDQXFG5raQNo8DkZOt/dHtixp3bqHtZ8tOftSqV0LvOZovKBpA1zIjOrN/OTt37Ke9Pz+VauhLMrIkOfMwj+G74nXnepazwZVP1iG3HWfm5AbZ/RSH5+eO4Z+8px5JC/Y6NmBD/2w8yhaVULiKGO0uoaWrWyLJ2YNZFIprGyVuCEQqqLUKCJ3p4u2S7yXlcIYkTjWM2XUa40UKq3UGkA1WYAVVr8iswWRaNSE6jYduCW1CO0FWTfTOCMn4sKRTLxoxFMbJnQXqfoIcdqt6wkgvpcKwYC8Huk1G8aacCf9UaGNdCff+/PU4E4zk7Pu27IWk5D/bj12c6VQqC1p7o5hr2sdlxWgFSlemZsZsJ/68FtnV1B5j1VzJ7P1YUk9CrP0wUii4jranE/W+IewX9L1wuBe25/8hN9ZVC43qHzd259cc0S2ONn8/MfnTUdcMoCvfn3sljb1D9pbbr3wmuu679pX/Tk/k596LJjdRY6gqRlUNiz7+s8Dy6IqOysCu11SUi2LCcfgM0ZGut9s2I00rHUiJohOtV0u32r9dPHaf3kv89qE/583Us3h9I93kyA1v5lOTH+nvLz2bnqgGUPgnnShVNBuFS8zuUQQNWpfc2CSj/XWX36AtnvAb6E4vr1a9FbPErxyrNBa9bmbx5E4mcUIdzly/rP5i3jlJXoiXoi/9w6MHkfqHjv0cD7f/ozfAW2OJbnuz9CB0RwEjMvWfUorg8PtIAoG956KxnfRFmBycLc2G4e3VWx6AbvNuhomyzeebNZceLlzxsgiTwMHVNkc1gNGVPml2lMNR9kzdflwWK+jzZcIMuMrDEOk/ie7TA0z2B+ecaCGnSx/uyAYQGmA7tsgXgGPFiBI+lx0cJwjR1Gr0XaiJp/IRsTfnb/mTqHoGOweuWIpHA1O4h1EAnZtc9l/ah5NBJAELvHZTX4Dc5bNBCEINvFH6jcDIXoqhlncxtUloiacylB6OHIM9MOYxsSUGKbV7gkv3ggyxaqzWFWRYMj/q7BGA/DUBCVGv+bBS0bBdpqMbeCGzJVG6Y84a9PfvErHaCC/1jBcU6pUS2bBN4zWPh+WAT4e7kZqCDjnNebBVAmm1aRH4wEkevtkYqDsNTy/CLeeO01NbkeqCDjnUDFzl23yZu2byirPIdsOiuFw2agot0MdsK02Uz6ayqFAFnxZGbVKPNtKpxMQEU0hGKlojXRKK/j0okjaFeL8jGXhyUZlQzec/ZgvrihbRrZQmLBO6DC3wv+rhC5JnM8rMn3XvT2XIURSsTR18MhIodhBqqdPXMGp06exMjQAEbHhjWcY5g2WZSk0ZNNZXYWZmtjAaoWLhnrKDWSKgpqdXq42iCDAyQDL22tcsB46dIlbN++HUNDQ2al4YoZ/r1vJOyzWlbFnt37FKzN1sjikD1QYWxX/+Xl3fyd10DDtE4zYsNLX6A6LnkHyOF1YiG4urqI1w/+ELFIDalkBIMDo+gbGEOpVsF6aRXNegUTW7Yik+1DNJHB1RvzuDR1A8VaHS89/RSeePwx7LnjDvQPDkhB8sMfPIVnn3oa1VJBAIL2MOcj6i25BDh4docrFD3ga+yTNsLtBqKoYXJ0EFvGR+T7TzZqMp3UFYkEQxgZHsSO7dvEQt+5YxveOPwGRiYmEQwncGVqFs+/9CqiiS5E4126D7yfv/Zrv4YPf+Rjsgrg2mBj15uL45WXnsWRQ2+iWSqLMV6olFFg0HkwgN07t2GkL4csh7jpLlybvolCuYHVfBHlRgXZTDcCrTaK+XUM9PcgHGxhfHJEoNv83BpW12u4Nj0vO5IHHn4Av/Dk55FMppX5kBvow9uvH8JI7wC279iBlWIeud5uDeVnbs7htdfewEc/+gS+/m//Pf7qr74lP2V5zrs9djNQYSTwW4GKjYEhG/G2GJHcw8l2f+iDH8Q/+uqvyzbm7JljOHm6eafRAAAgAElEQVTsHUTadSRDQJz+3M7LOx5N8QQR2bzSiuDi9DIOnz6LcJpgXRKXLl7B7MyshiC0XuF1Vh4T6pgYH8Lv/M7/hg/c96AK8lg0gJHRPgQDVJqZzYTOQze41X8EAlgslPDjl97C7I1F3HP37Tiwf7elAgQImNAug2cTgXWCdAnwkjz11NP4sz/7Mw36f+M3fgNHjhzB1772tc6+IM9yP1xwgJl/lkylZWxG7Z0C720v0oCX751qs927O17qDz30ED772Z9XsDMzfGgfoeetFRCbmT+rDsc4rDfxzttvYebGFOq1Io6+86ZsREZHxzE3N4e5mVmdqaU8maIZJJIxMGSXP5tf165d095G+yxaZ+3ctQ0PP/wIHvvQ4wo/NzDeRlYB/swAQc4oLl4jUFHD3MIqzl24jP137REb2BjNzJiqiBlI8LhUpeVDAj09PYjHkho8dYCK1RUxz3ds3S427t98+y/x19/6z2g0mRtUNjuuTY2Nv64KTEVbDGgyz5n/MT8/i3g0ijTtMlpklnKIQ3VjFL29/di+Y5eUK30jIxgaGkW90UYi1WXKiwitDjjgaKrmYH/G+ufNNw/h33/932B5eR6tZg3JeBTd6Yz85wlYUOkiW656DWuFssChqjzNraFuOzWQfM43ffnhtL8PHqjg+jDlpilvuC17dp3fcw3kCMiihEM12rz49c7v0TPMf8uayA1iPQtSoK4UTTZY9T/fnxkcsCbTMYyOjmBseARjo2PozeV0LTjk2bt3r846DnvEhtzEMhyd3Klzlk0hGcAMZZUaiwP1JgfIwF9961s4c/6sGtAQm2vaWpFY4RUVHNbVK5b3EDO2f6ep9NYK/N0Pwt3yDLRtwEQFobeF4nkooGHT8MHvb1w7JLoQqCAxhXZ5rKtkH+CyWpV2QYBCmSVmg0qGsQZ9Cl517D6n4FCDy8GllJFWT3NzYY1DS6Y9u3dh185dZvtZqVqGkrIqnIrArY/llWUNanu6u3Wd3g1U+DPtVqBiBqtrqw6oiDlFRaSjqLAahoNbI1UoFLzFLIGYiAW0XWOfQICZ9ohUsZSLRangNEiNhKTUIxBCsgOf35Vr87IP0VBfIBvPPYZjsoewIGPv1e3ZmKwN+P0WMmrgAMcXGmAGef0JMFDVaYQLDnI55OB5ytqXn11EIBd+zZuhgayIUNwjbc3zNfywjddXrGgOifV8mSXGxhnhAtYDQdXYAoHcs+FVR2b9QuIIc4U4MDXrEwP/nFm1s+cxS7+Q5a6IlUtVjBsEc603akgno7J1o23iwGAvHvjEh7GytIyDf/sDs2+tVURA4aJcWy8hX6jh9/74nwuM+93/+fdUM8ua0NmdRBMMCK5gdGzM9S3c/8wiR2qOjle31a68CcqQYD8gZYlZ1/Jec+DnewK+gM8AoW0e7xPXEnsYAXvOQ55WOnxWFSy8iURCxYX1KzbgNLsXAxV1/QWE0GophSuXr+DM6TNSZrCHq1bq6qEIIFONnC/y/rN3JZmA150qNBuUkYVPohB7tHQ6pc/glUPaA2Vz6gJbnb0N+z8qVx544AGpDVlr02qzXCygqyuJQpGKceaxMBS7ruB7AhOE6gkyoVlDcW1FmSPttrGsg6EYYokcnj/4BrK5QSysrOp5Wl1dkfqBz6gshF09SjUMAXuqBvh+BocGpdqkRfHM7BxGhwd1ppgdcVhAMD+b2WkFcf/99wuQIUgi9SaBIg8KcMN1/TC3FoGItHfmEFxgLh0DDLziv/G++QJTuTc522afdcGznPeJDH2+Fhn0vMZGTmKNw/7fkcxEMOR7YmC52b141rwPGLbsJBviKuxX1rdmKyQ1hxwkvI2PAcHco6REcIRK3lu+d+1dfC6dDadnVPNZlgJKMwkjmonkxrBy2oA5MMdmBmYRpnmIC2nmetJ6e5eqSnWlyIFmt+SDif2+QjpOKhZGPNTCxHAfInQ94N6RTKPahGp95pP09+ZkFVsurqHVLEvlQ9vXao26Afb12ixRrDYQ68oqp4JB2iSzsc4KkIDF68LnwBEb2VsT4JTKUmHVLfFNaL/M/cFqAGPg+/BtXifa4Gmfq1ZkBSZFlbMkMrWYAfOsx3R/eJZ0Ap4NXObPseBjA6h51klV5vpsZRmKJc8cDJtldc4D1SzsIwxoNICkKQDAq8E4kOdZJPBF5ARmqRLUsbVjOUP27+zemqKS94j321v4+XmYbNGqNZ3PRpRwZA6X78LXE/jgMxnc2eCBPA9yCLRwn1VkV5dhxXNC8ysSINxreYBho4faUH3zYnCepLwo3lP13jYD0DMUj3f6DoJ1vC+dz+JUFPz53qaP/077NW3JCeyz7uqcWwbybe71NmdU3Plza06FarCSgVkWcu2BQO5bvH5mUWVnrmZxDvzz8xTVo6439+pHT6RhSaVZpgPAVYs6kNCD5qpTHXJu1lxWLDmoxbV3GyQevmP+XcdS34GxOpscScjcV4wF5/tbbztqbi1c5wbS+3ulvYqf1bmz6D28H6Z9S2/z/v/4H+AK/DSgQui1kxj6zUMPhw5XhjBZU8TNW2iyY0rY95oXqm0FBAdMsmmhoDZ8YgNhLK+gIb9icbB49Cw7Ux9YSLVZTpmEzWRRJm+zgCUxiGQb4IKHwvQNN8WE35iMob8hP7PGxRgc3vP/3Sg5Gzduoixo+D38nfszDxhZ4LgG0Qf1cTDGYS4LLDHg5AVOEMWkzRxQc8Mz9Yh9Lr6PTqAQGSq8FrQ5UvNjFlrajGQXQL/uLiQkdaXMzOT/tknZEIyfkwwW/35ZuPusDTLE1CDxHjpPYRXzbphFtpCCfmBFlrHnzRqC139tfc1lOaRVFPL6mD0WPzcDrg2QsHvO61rW2+JgjH9HSSj//Oee/NItQAUPZTbSbFQIIKkBcY2bZX5sFHAeOCI7UkCFO0CztH4qFwVU9Pb3qbFi7b40M4c3Dx1Sk3sLUBFPYMeOnVqTfcM5BQbmsjmBEu8FVPjGxgd4iekRaGu4Uak2/wFQweK9VFxHZX0FF04eBWoVRDR4YLPOBsWFiXq7C1c481narKjQoMjJPdkoEqjwAIeC7splXR8dyJEI+vv69GywuGcRxGbr6JEjGBroVUZFJtOtjIpGvYVoPK6GmwVguWw2O+Kqi7UZUtPPdRhNpLS2aL9gdmuWDmDgo6lC+OydPn1aw6MdO3YgnUlb8J+zuBALV+vbJJD8d9u37cTo6KSskvi9Ko+kqDA/bv/F16f3Pp9lDmclU3eKCgEgVFQ4Xodk277ZcKwFXqNKuYi3Xn0BxfUZJBMh9PUMYWx8u3zJC7SDqRXR3z+kYX88ldPg89zV64gmU/jxM0/hEx/9cAeouHjhAv7i//1TsZsbVPHIr9SKR3+/VEg6VqtvlNVMuIF1R2LKwVitjEQkgD07t6Evl8WlixekcODnpqULraom/3/23ju68qu8Gt5Xt0j3SlddGo2mSKPp3WN7DLaJwca4427cAdOCeUOAUN6EBAfC+yXrg0AoocUxYAzGYDAGjI0buI1nPJ7m6VWaGWlGvV/drnvftfdzzpVgQb7v32RZa82apnLv73d+5zzP3vvZu71NkxsEkHft3oF5CzuQL5ZhYHgCzzy/SZ6x1XUNsibieti4cSM++am/xfDIqMbzeR+rK0OYHOlXOHjvyZOYHB/XpMrE1CQiFeVYu3IFKsuDqK0iqVGDg4c7kaBlSjIjQqe+th5DAwMiZhbOb9UkQXtHm4iJ4109qIw34khnN/oHh1EWCeLm227Gtddcj3Qxj8bWFrzy0stoqWuUmvd4X498+UkeDAwM4cUXN6G9fTE+/jcfR09Pr6mdSiqnYomsVIGsKnWGyPLnk0A/Wc/7dUyHfwg85kTKHXfeietvuQ4nOo9g3/atmOjvQwWmUUUFM8e9g+VIpacQipVjJFHA0Z5RPL9tJ4oVZbpOnFjgzydYxUeA+5TOFLBRLeKGG96B97/3L7V3RkJFzF/QAhRJVPxhmHYJjKVaeSqF55/bit6eQZyxdgU2nr1GmSYikzNJ7Z/ZDO37Yigvj+LggcP4xje+he07t+Piiy/WM7h582YcPXq0FLLomzgR8WoCzDLR1qEFuNqkHoHBCv3uG3x7f8ztaZKCnet4zZo1uPba61DX3KrnlN/LyMaIwqP5vOXKrHmgVQv9wn//9NPYsuVFpJOTmBwbQ3Njk86Mgb5+e5YLRWVP8GysinNfM9Cot7dP/8/XFa+uRHNzvV7HhRdehKuvvlrPvz60VxUwHeBkWEQTUGOTGfQPjuPA4aM464y1AouMHKIFREZEBV8DLQLpbd/Q0KCMA4Ze8/0Mj4xgbJTWTzEsX7IEB/ftwWf+/m8x2N+DYBknAO0cs6bVyNHZH2UBO995/+pqawTcEIykDzgnK4x8pp1SBHPmtCiEmlZXFXW1iNfUipziu+KebFN8VF9yXzYydnR4DA/84Pv4zWOPKsi+ooJTQAa8c9KJ9hBxWrVM5zE0MobB0QkLKeb+6vZc1UysTZxy1e9Js4kK3gcRFZqso5iBT6KbqNBU68y4vBeuyDKnQDAvKYDBWwn472u5CXZ2qa50/tNm4xl24c0G3rnCTb+xtonXxkTocJpiTvMcNNbV6cfyda5du1YAKtc89z0j0W3dVze2SgnKT05NEUyjhSSnF1iU2HP1gx8+gKNdnQIqQuVhnQfMQyi4moOToAQMed1IVJAIJiCj88zlEBj46xpuH2ooosKAFNZgAg6oZJ+etmB2iWq8damtZSpJx0aoGswjTLW0iG/+j78mTkQQimhqQkQFxQ5uSovXxLJcZizmpsts0oM1KQkLiRMqY7q2zEbasH691mJeOR/MhMk6mwbXZHOPGhmWvz8tRux9sIa3qYtS8/1fTlTMIiq0v1iYtoF/JCrs/CepJKIik8XI0JDs/QhEcjpiIjGh2pAThhoUiQRl2UHbl2AxpEnY0a5eVw/y+ti6kqApb/eH798EBdzDCGT43Ap7lqWsdTYUnGSh+IQTpv7+mjjL9kfzszalqgfLBUKVLErsefGiKVNIm7WqJxRmwAYDs3zPJUUqQVLX3/A55N3wE268d/wc399YzWE/m5/DDBe+D07+WP4Za69pJCbGtafmchpF1brgteR6j5UHkU8nUR+PobmlEVfe+Q59v8cfehQjA4Mo5ni/uPcF0XNqADt27MPDzz2q93T3bR/D8MgY2jraZRlFAJJ7OAHwNWtXqxbkc8T9WNMGnPJxY3Q2wcW1b0T17e++Dmefsw4/fuBX2LJpZwnYU73t7Fp870iSide+tq5WYpTEVALjY+NoaZ2r986fa/WmeX7z9TMTzvaIoEhrr85mZgenEAzINNsQnqm0e7QJFtoP0iopr7p5KmUkEa+HWbDxXHUgt4ArO2s5ncczgYSArGfc2el74RJw5sAmkhtnnX0Wmputh+F9owDKCDDetqCFlFfXaLKI9ywWYbWQR6hYwHA/7c+4A9BVgAHNRQQravH7l3Zh/ZlvwJ79BzXZ19t7CitXrUBvX6++Z2JqCk2Nzbo2tAqkUGB4eBjNc5o0Ld22cAFOnT6leo25EVyfk+MJ1DU0ONKNU3ghnL1xo0RwPPusZzAC2UgaJ9Zwk2Gy1HGqYQ/88ms4icOv4TlM4ZZyWhjo7nz3SwA+LcKYf8L8EAfeSnDhJnKszjLAlt/PxJDWe+tcog2b3CFs4sFbKPsJEp4nvD/cr9nH0G7YCxstENycG3h2GIlpdleysHLgO0kLESGu7idAzueTH3xP8vh3UxNcYzO1mk0I8BylA4IyWLh3Owso9nec6JEgzeVdaOd3+RoedLU92irjfHoKhcwUgoU0slPjiJWThA2htrEZU+mcpkNWLl+KEA/HaU6rMAPJyKUIA7Ongc7j3UhMZZWLVwxGMMXel/ZJlXHZjAkIp30X91pXp8nKjYA3cycJkJNTo/1YrAL1DbRHNUcNXUtXxJv4gKJFm37gPi/Sx/VZXljq+8pSnTHLlkj7J9l74h4ij8qEWWiNuIlG1rC6R+584D2WzaVT6Fu/Yc+1v6behlVTd5wSIU7iXDv4M21vNutu239MvWC5FiZ+ZV/n93O/v2vCSkB+VvuGERVWp3sCwuMfXAvqddy68mA3f1eGarBMZB2Be369nkEvVpB1gjljmIDE6gvVcP5jVmnrrY5MXGeCY7l1ONtvt7xs5ssRJ0bcOts+N9XAr2VdLwzFZcx61wM/LeCnKvyUxr4n60sviRkVXoAlrI9WYVxnzgLRf6IIQGeNOdtiU3bvwjU5ZWeEjUg193zyLPEiHKs9jXQWuuYmm/n6vNihROzMspj3T5v/3a8jj13q7y6o3Mi5meuk68s9kh0lz0knfDQM0M52c6xx198RKqpdaDHoPl4nKmaW8et/+h9yBf4rosJvinyrfIj4QFDpZSp/a1bpYUxQ1oLiZj6PDzT/jYUEN20f+GPFQ9EADtc0cGPmAe3tUlgschNQ2KAbDfNsrlcsyTpFxZ0F1Zo9gSNPvGrPqYv8hmJhbZ615fnlR1/LLCNBh6w1ufKODYcFvNqmxdHYvA4RAhu2t5t6yvwAacFko+UaHVemBdVpZuNjkxWm+Cs1IPQi1sFm4If9Hxl3eogSBDNAiYWUBTlFpWxR88oNjWG9rngTYeCKJJ9DwZF5vi6+h8FBju9PqOCiosAC5vIKcKTqkworboAsinhoKPSuaCSKVCBi/8MqRlncqRGUAsFUKDo4GMobNAUUb4eUKAVrEKjM8BZQb7vuRnlU2rh3QAHfCt8j6M5ixoFAvB78uX5ygESRX5MsKEhU8HXw8GlsrFczGyoPqbgmwEPP5cToGDa98CKy6RQ6Fi/DnNZWelMpz2Ep1YQIoHlenYAMWkrEKqs0DUHLmrHxcRTyVA0QzDfFB++hZ/wLmEYZPeQJetADNBhUsB2tn0jSnOo5gcmRARw/dEDhZQz0ZWEk0NCRb6Z8MMKH64RkDe/RH6vzBVprhBhSmWjc06k0eI957fIsZKU8MW9pFn/9ff3oOnZMGRWNTQ2oYigaPTkLZgnGdcD7LrKDRYizcjLgq1LEDRVcGrl3IJ15g1oRRaWtb6qphj558iQ2bNiA6ppqBbYST/aKSw9S+cKoqbEFq1evx3SBII+zQPMZEy4skF/D9zowMKDvQ3CRTYIBHdbcsoHkdZzJK7Dii7/4nljQJJMT2LdrCzqPvIaaeDlq4g1oa1sqn9TxxCimUpOoq2tCoRhEebQWew8fw6ET3WhbvAQvPvk4rrzkYixdQd/7Gmzd9DLu+4//lAqVqmb3k21/dECECh4q/Nx4v98/Pbik18WGRgpeeqKn0dpUjw1rV2JiZFDvl++JQE2sMor581rVmC5dugR9A6cVzJsvBFEIluPJZ57H6f5hNDTN1XVhTgGv07ve/R6cvfEcKb5sTHYaVdEQJoaH8cyTT+L4saMCbicnx5UF0D5/LsoKGbQvaJVt0v5DR9E3PIZUroAyqoYyWfSc6EZDXa2mP4LBIjoWL9QztHfvQdTWN6MYKseefQeRpiqxuhpf+uKXUN3ciKa5c7Br2w40xmuwdNkyJDIpDI0M6/mnYuvkyVN46smn8fTTvxMoRoU4f/nr5tcMldECLJwiUffdZRCVwCMHhvpnwFThQVlT/OgXD4n4iYWCOH3sMDr370Ygk0SEVgPTnBpKIVvIYWyqgM07j+HZzVsxlp5QerdvPExl68fzScIXEAkCHYsX48N/9dc4941vUPZCS0ujrY0yex++iC+dAYUCBsYnsfWVPeg50Ye1q5binI1rtR/zOc9qIs1swhhoyMmThx9+BI899hsMDPWXQkJ5zz0ZLUWfm0Ljz+OzyffPn8m9xcjFGds4v2ZLgIkjKvh3Thw0Nzdj6dKluOOOO7Fw8XKMjo3rvZvFjJGonBQoi1nWBwF1qucOHziAxx97FNkMJ3f6kFVoYRn6TvdqaoJTAASYqRSivQCBEq9A5P8LWAgGUFsX11rmdMVNN92EK666UhZLBGT5/7kCkdhyHO8ZwOhEFr39Izh8rEtEhfy1nWiCZB3POirDM5wOqqlW/kZVZTUmJhK6twMDg7KriZVHsWL5Mnz33u/ggfvuRaFIJT6bBLuHpV7uj4gKxyioxmCdNLelWZMVPP84ZdE6b77VM8Ew6uvqsX79eixbvgLFqE2scWrGAj4rRYJxT7fmPIDxsUmc6OzCV7/6b5hKjOuMyWYTUvtzMqWi3AI2WcOMjIxI9VwsY0CpBTpqYkHgt/nk81w3sGZG4GD1GO13CG7atKl89XVMG7goH11HBGuPVXPlMk7yDA2mwtnWo7fO8Oo3E+FZPoWJLe2MEkAjfyPfaTllmpreAGoaYpjbYkRFc1Oz8oQ8OU5SnGuUr0N1goQ0ZaiqrkE4ViNygOc2ryVD0TW+L2UJFdwZfO/++9Hb3ysAPxgJyWaJwC3cRAVrFjtObYqQzxAtLlR3+hwCR+yz6SUAY3sW6yMXKOpUrgw15/UneGBEuzu/pFU1ooJh86l0UmtcdZgD/ByU4NTyJGAdKU7wTX7MNoVok89ucsvlXfG/qHClXZKm62KsUSpQHo3IPuvMDRtQEYoo54Ph9eaN7vPPyjA+NoaJyQlZtlmdZ1O3vg7iddDe5sB7XqtTp0+7jIqo9ilNTrFmkV1MTjWkFy3o3zWtw0mFcjXpg/0Deo6Y8RKriGIyOSlgj/lIsqVkRlIFM75CCJcx5yuCieP9WqP8eSQD/XvgfdDEhgOd+PPkre+IBgJOqiOdell7YrnVadyH+J75NUY8cA+wZ4l1hamiLTBUXvfMJJKVmd1bv875+nzPoD3Y1Wi+7veAlLeOlHLX9wuOFDNlqgFPXlHtATv+H59/P/Grny0hk1kHkWTjNJi6MfVKZhPCvirAnJsADfQKqK6MIpDPaxJ3dGwMa9esQayyQpZNBEsYlD0wMIqtr+7Gr17+jaYW7r7t4+g5fQrrNpyJzs5OWT/x+rHuWLFiuep7hcuSgFfGgLPqmTUtydfD9/Cu996IM89eg5/86DFs2bRDe1d5mLYh5g9PUJrXnkCtTXMb6GbnRVCh3KzJOfWgyXJN1ZmVkN+7PTit/U6ZDEnVkLIsymQsYDmZRuexo5hMTEmgQNKFa0pq4PKoQGKdd3zdqtcteNlPD5DM415oQoOMSJqi7PYMGNNkjFNre9KJRFc6k8QZ69dj/oJW24do2VMw+yo+w9x7tKdpHRYRISFSyKA8UEQ8FgVyaUSCtNrh+g5gMplHFjH8/qUdWLh0DQ4d69K5NznBfL1qTb2QFJ8Yn1BvwPVsfatpQXjvRkeGJSbgJID+Pjrmzhoq6c1eiwQuz/MVK1doCoyiJp2/rr9VZqGIWXsmeLbIStdZ9nCv48/mv6ez7PkyynqSAC7ng2uNlOd1NXCbREdea83nuLCeFfldChP254qJRSxDzghjO8qtRuJ74z+YoJHPEsPMTXnPz+W+ZP2O7cQ25RoxIZab7uZr8tNyXIueOOfPJCCp3L5Amb5OhKiz1OHXmQW1ZW1wfXNtsxe3vUKIpKvh7TXKv75IHMUssLz1s4kqzVefr1eApwgaSAyVmRpHIJdCbmpcQqDEVAZFTtQUbU2mEgmE3VqKV4dRV8/ePCxrypr6BowMjYFuUQMj48gXgxhNpJQBlS2QlMoKW9AZ6KYABUBzLeWnwcxEvm7ec14LEpoL29tEdCnHxU22Ef/xJIefDiaYb/urkfMeB/B74Ww4zp5rTkjwuqYRkE2ekZMSXbje0uoaOxP5NXx2RXjxvHCCWI9zea0AwX6/VjzepJQ0l+ni62gT3vAe2BoXFuZyt2Q16jAOn3ehWsJhbLPXo8K7KcCY5UogkY47P9wRU8K+RASJ/PW5US4LTFOINj3NNSHMoZxn0kwv4N/PTIFrf7KJFJtM8NNMpX3CTYgKr5uVySJyShNuFDW7PZI5IXTO4B4tu3cjeNUblWo/9ydn+fvHYdpG9th0i98HLP9ixqLeT3aqPnVWj3Y+uDwOJxKWgwmntBxZ6EkDL2DQa5MQzQgX7Yveykp2ee5Fz8q7milhHT3orKF83exJL0/2+P3EExpu5LAUZl6aINSUpxGh/hzzz4hp9maYpdeJitm7wet//h9xBf4r6ye+QQ9C+qZKzSf9JDUCTi81F3xdYgZdCJobpXX1sgvGNi99fi8WIB5c8RuvGgf3wU2Fh6+NYNlD70ErbvpkUvkhBbpXaLgASD6zPCj0s11DVXq4HTiugFlu2gye0wiqNbR+0+LG5NWmbE45FcD3a9MHVHQxTDovS4nqOAkBU7WzeLSf5QIQ5QpgDYMOI+fLbL+bqsPCvGi7YyO4BibZpq5vU0Y/2Lj8r8fGR3Q9WNDRmocbNkMG/SgrQRAWhQxcpfqU18esk2yig3/2I5TuVeo9iVV2Y4q+QJNns4orG5OlYokHONW2fG0WSJZUwaSpCmVEsDBPIRgyNX06lZQlFJsTFuEEu9/y9mtLRAU36koFx5nPIxV9XiWhdeKUkrMbMxEYVI7RdkWEWBkaGhswlUrIg7m5pRmp5BQKtL8YGsWmF19ALp3GIhIVc1sFoNPKhRMVZFYaW2qRTk6hrqZejY1sm1JpjE1OIp8p/AFR4ZtrHfDUkmj9e6KiTI1eNMLAwRHsfm070pOjKOO4cSZljRqtShR6aYCQV+Z6z1I1py5wScFIzjLIExW0neG4JccsPbnBdSWbsGhU35ckDp8tWhTRE562Vy3Njaipq0ZlZVwFYoAKMn6fWMxNFZm9FiEPXuvKaFR+vAQ0opWcjuCzQjLD1KVGVNDyjQSKqfYIkNOGhor5JUuXChywgKgZT8xSgYMiqqpqsX7dRoRCMTXPUoQq6NWUjR4g4Psk+EYQT3Yt9KdN87WYupGiGa9K4nPASZfZRAULkFRqEieO7cPu115GVTSIWKQKra2L0DynGclMAmOT44hG4xgcmRk2eZcAACAASURBVMD4RArFSBRV9c0YS0zhd4//EtdedQUWLFwo0PRrX/437Nv5mmzTuC8UYWoGD/R5qw9ZeLl77H1J+XlS9LjnXIUKLd1yKcRCRZy/8QzMbarHia7jAsX4/+Ewrc2qBeguWb5UwAJfY7SyBvlABM+9uBmdJ05rooJEKoP1aM02p6UV99xzj0A77nN8JmklwOezIliGrS+/rFDe8bFR1MWrsKR9Hua1NiAWKkNNTRw79x7EkRPdUk6xmB8aHMbpnlNYtGAB2tvmSbm3sGMBQmUR7Ny1C+HyGOa1deBo13GNklN1ePcHPojLrnk7mltb8OqWVzCnpl7AN6csJqam1HRt3rwVv/rlr3Hw4FGRT1R20bqNo+kKeHagD++xQPhUWr63/jyYqXEdCCBVnTW3WtNuIom5C1/7z29j4byFAjpqK6OYGh1E14E9mBzuR3i6qBDBiakJbNm+D5u3HcSB4yeRmk5Jac1Winv9goX0xQ/g6NFj1jAph6UgS4Vb3vEO3HHn7WhpahRhSnCINa1561qT9cdExbat+9B9otcRFesEUhI4SaQY3E01WB6HDx/Do7/4FbZu3aapAzaDCsx1gJYnUPn9ua/z3/nLT1eIvHT2gWxk/Vr1CiLfYPkz0wNejY3MklmL226/A2e94Xyk0sxoKGpqj7eFE21seEKV5Sijv3JZWAQ6rZ1e2bwJxzuP4lT3MXQeO6wzo/vESVlJNDc02tRXmHZSsRL4Fo/HcfjwYa0L2mAEw5ANRkMDSZMGvPvd78Ybz30D6uuZA0F1HsHlCI6dYJj2tAi7w8eO4+wNa5wHuxX2tHdKTE7JAiibzyjTiCRCVWWNgoKpPO4fGMDI8IjucfuC+fjU33wUO7dvEUkB0H/aLCP+3Ic1HdZwR8IhXPCm89EypxlHjh5FtLICbQsXaipGYGo0ihXLVmLtunWoamhCKstcBFMk0r6J5yD3b5KdtNXgGMSjj/4Sv3v2KYSCJC6GUURG5He8ulp7IQEdvr/x8UmEIuUIkwApmjWFD0pV40iAR7SuvVaR0K7J1NSHE2tY7WdEBcEKNfAuIFvvlVuXC8jWZZnOmiVhxmoOP23hiQo/su7PPN+kCcTV/KP7cLYC1swB1fUxtM6di3lzW9HaMldEhfzM83nMaWnB/Hnz9FwRKCHozDOpuqYWwfIqZXNIXZ5MiqhQdpaQKmBifAr3ff97GB0bFYhNMpYAiwBdFzovooKTk2q4CwIued7Nfm58bcnzmoIFqSsd8cLfeb95ZgdDJnjgLwPErLaS9zMt54rTmJqYFHFMcIt1merUUl3sxTiseZz1E2s31/TzeTAcbaaO5vuSxQEBDEnDXf5VOIyqeEzPAEm5tnkLdZ9JKHId6hx1xJUnKpj54q1HfV3tz73ZRAVfRI+IijFN+VREbaKC5IIRFbYv+T1LpJNeJ58Ls7UZ6u/XfaqtrtE+wak/Al0xp1BnJg6JFipto2ESnuUYPnoK0XLLPSKzLIAhUKZnTYIJTa+abaoBm1RM2nSPamB3bug9ugm0T3/+I3r9J7tOYfmqxeo7OJn1/LOv4He/fUnPVUWsHDfeegXWrF+h98jvzfDixx55Gn2nB7Fh42rccNtVON3Trz1p3oI5Wuh9vYP45U+f1Oe6ZkXAKPf8lWuW4uY7r8bkREIgaWNzve5Hz8lePPKTJ3DkwDGsWrsct991HRKJpMQMDBd/9okX8fgvn8VFl74JF77tPFTXxvV1g/3DeOKXz2Dnq7tx/a1X49wLzsaLv9uK3z72O5QV81iwsBl3fuB2JBNJbHr8WVx0/RVITEzgvn/5GiqiEbQtW4wLr7kCc+a36rk/tO8QmpqbMDGZwF+96+9EVFx82cV4x51XYQOnAqm4n0zgBf2MFwWUfvqfPoRYrAInunqwYtVSiZ54LZ964gV0Hj2B9959q8BzdzFw+lQf7vnUlyREUuaD83Hn/9NC1ULdC6qFBwYHMTQ4qOf8RHc3lq1ajRUrlumcYt3DXs1IHsvIUd9F+xjnAKDnSfmFBkZzXezZs0ckhSbh2Ztxj+XPq4prT9UZ6zJX9Bz4SRcC3tOmZubZNjXFfIsAQqz95YzjVff8u+0B7BsF4qWTWLNmNRYtasPIcL/CjAmc8WexZ1Euop5zBhfnUR4sIhTII5dMoCIYRG0lCZEkcmnmDQCBcCVS0+V4/NnNaGxdjCkGC6hHS6K+oU7ZMyLZsjlUMEMpEJBoQEr26azlouQylnGmgPIq1eHcSrjOWYsT4OV158TVsuXL9IxkMySNbRqNVb0cEEQssBY3e1/bX7iPOVtBR4DrjHXBwPwcgdGyhDIi0+oYE06KLBTRO5MzIRsfGJlo1tQF59xg55PseVwgMskUnmsiBijacna1IiDdOrH7zExIswnT+pA1FDEAI11570UyunXA889sxQyxZ/1Nm1Mfpi1i0eVTeOspZWmlUvq+FNopYwtFAbsirR3Iz7OOjgJ8vXxtvq4UIeemjriOTRRheUVyNcgkURePoq21CYF8Btl0Epksr18Q3af6JRhimPZ0OokQs5oKKdTUxpBIWMZmXW0dElM5CSA4ZV1eWYO+wVEk0zmksnnQbk0ZCeGQyAFZ0rBm4GvksyWA3iyheDySaF60eHGJaDGbTk47WKg8nwcB8k457oV5ElE6K29PVPhJBk8W+Rqb5zEn6YgXiKiSG4jZL5IQYUalSGiXz6aejVkbbmKthNlwDwiSZLLnQCC7E7DKmpElhUSdM/au3K88me2V9AL6SdSJwDOjYn7w+8qSzAH0suEWLmT4hiyvKBD0faYj2fn/fjp29tQEiS8KDVkTyZlDOaaWl2Pvaeb7CYz/E9MU/rUpn4OEvZtUssxSwxxEHMpdxMh83z/4zCDlsxEr1GSRTTT5MHvWuqWQayskZkB4N/Fx8JmmUlm4+tIRm0BwUwmlnsbltfq91L8/YYDOxlz2ig5T0POi51gFgr5/qZ51Qmr/PoS/ORzRXFDsefLWWaqtuLa9MKH0amf+oDXqvtbwE/aAtgdxHfr9rJSJ40LlVac7vFB9nc8Z8dM+GrEzm0c/yanX/br105+4C6//03/rK/DniArfRJpay9hebjTlAlFY5JeZ8nX2JIMLzZ3Njpoi2kaueQh7lpVgEw9kA+lnABw98Cza3IiWBQoZkG7Y/wxpwQvvRye16ZesLYxh9VMe/gbZ4WVgFjcYkiyeCOGBwlFhAi/eTsdbX+lwkb2v+akq/Eg+w+a7bBuNKX40BugOD702V5RaGWsbj4EFBiYpWNsxtT4czzPxnjQh+EjrCJIho2MjoM0RR5zZ/DE8mVeEh2KwzMgbfp4mOAgasPCJUL3C6QjzC2XzyA+qMfizWVQRANZ7d+AoDziN6ZGgoV9seUSKV4GFGarIzbuQhw3vl0YnmX9RBim4crLJoEep5VLQMoPhSSx+33rN9ci7EXm9niqbqBBRwckUqc8MhPZEhVeTeZUZCw/6z5v5QBF19XXIUE1UEZGvqgKn8zmM9A9iy0sv6Zos6liKOS1zpdyLVsWxuGMxguEIGufWCMSgtQ2VNARQGRDIEedclvkkBjD4EX+vppxNVMi+KxhUiGxFOICpyRH5syfHRkyhUhFBBUO8qCzJOEWQAyC4Vnlt/Xuj2sSDOSpEnJcp/8388c1uieuN91CEGom1eFxqHfOvLaD39Cls37ZdKrHWuc1qZGkhQ6IiHKJ3bVREBQ94n3tBsII/k6GV/L5sRMIVMZfhYpZeNiJtORGyCXGqbd4/KurYtDAIl5MYXvmj6SunXPHqwbJABOvXb0Q83ihFrcO+UKR/qn65CYVwSGQcp4K4Ti0o0ywk+Ds9qE3pQCXPDEkhMkCfw/DOJPp7O7F1yzOoCDGbgNYvrZi/cD6mkdM95+LdsXMfXt2xBx3LV2Pt2ecoTPu5xx/FDdddg/kLFqCvrxdf+/JXUKAHLvecgMruUrHDe2QTVAaQ01LJExP+npaug3JbrDhj0F1wOosVi1pxzhlrkRiftMY7lVSjSLUfAZNFHe1orK/DeCKJuvoWBdq9sPlVHDzShWhltfZS2i6woWT43XnnnY933XUXqmvqkJUqy8gKZnLQKqDzyEE8/OMHkU8mcNlFb0IokEM6MaHpsK27dqPzVB9CFZXaE4cGRzA8NIIli9rQvrAVsWgYLXMbUR2vxeYtm5ErAh1Ll2NkbFK2UZnstCZC7vvhA6hvasTOV7ehKmLBmgc7j2L7rl3Yv/8gensHBCKHQmatR1CAllqEoXVPnRrSWz9wr2ZT5TN6fKHpwTM2AWrkPTHsxpH/4oIL8Ol7/hFNc1rU9PN8qI1HESxk0dd9HAMnOjE8eEpKyk2bX8W+gz0Yo61hLIT5bW2YTKSwaNEinHXW2RgZHsUPf/igMl/oIT0+NiRLvoUL5uGee/4BG9atQ1NTs8IwCwE2swxhnZlukEKnUMBwIolXt+5Fz8l+rFregXPOXqOJCp4VtNChcvOZZ57Fj3/8ME6f6sXkZNJUa7RIkwrblLc+KNQmDJ3+mrkyjujlNTKShCph7s32daYUnmkQfEHsQVTuAbQRu/TSy3DuBRchzpwSBmQmppBkmHYRAsqDUdodMtwzgnCRwBIwNjqM/fv2Yvfurdi7Z6eaxd5Tp6S2JtjM85fPCPcgvg4C81TH8zkfHByQcrtQzBlRVx0XUfGGN56Da665Wo38ypVr0TRnPqaLIXR192N8MjeLqHATFa5uSCbTjqhI6PsSwCMpUlVFdSknKkKyIBsaHFLGw9zmRnzgrndioL8HgQAnKszzekbZPlOLaP1Zn6WziH+jRcb1116NxoYGDI8MK/ckGjV1L+kBNsMkdM/YcCbiDU0CU7jHEZRlnTExOqY1w32NqmVmV/3LP/8LhocHMTo8KEuxysqIa0YzmKJ/eTGAFCcSQxFU8KzmuU8lZzZn2Vd6DnjNLatAggVnweQBD4F5ThlqRIXZkMl/mu/OWRz4+tADRrJuKBI4JMGU1hngmzcDkWxKQpNds8hrfh+zuTIAwaY1Zq4tb19VrYVpt7e1i6yoJ1EhG9GcQOj2tjazytT0XE7nFi1JCkGCbZY3wDqIGRUCIKTwBIYHR3Hvd++TgpfPDxet3h/BNQJaCv60iQrVo9M57YNUNRuJYnVrqdFl8+4mRQVIyi7KzmcKSDit54EGTcq46Vp7/kigFDTZOTI8KHCVoAqJCgFvEgjNIioE8Lm61NkolGxoZhMVzgpRgA+FD7JgtfDbAPM/olGRP6uWLddapT2H1JBOsUlQaHx0DOOT4wq1NvDRBwS7rAG3f/ypiQpOAUejtIiL2pSCC+DVtK0Lm5blkUAFO+NsoqJf4DSnOLQ3TI6LRKGAQsHYJN1jrGFIVFD9HMbE8QGzKivjnhLVNZf1B60U8qbgNXKE/YSFa/MMEZhH8og1nLPpYl3K9f+xv3u/rJAmJ6bwyks7NBmy8dwzNFX9w/t+gdOnBnDHe67DyrVL0HW0G1s37xTJQNKi6+hJfO87P8Ha9Stw/a1XGFF7/BS2vbIbq9cuw/LVi3Fg71H85zce1J7ONcbXy/p62arFuO2u66RgP7z/GPbtOYy1Z6zA0hWLcLyzB9/56gPoWLIQN7/zatV1A31D+vd9rx3S673s6guVDUQygtfi/Lds1Nr/2Y9+rTPg5ndeh77T/fj3f71PYdqXXvUWXHT5Rdjz6i4c2b0fl9z0du1HJCqaW+fgxvffifrmRhzecxC7tu3CWeefg2WrluFEZzf+8raPY2xyAvf+6CtYsWoxXnjuFezdfRjX3ngp5s5txi9+9hRe+v2r+PvP/y/MaWnS69r0wqt6XW88/0wB1z/54WOqcdafuRJr1i3DU4+/iBPHT+l9E1Dk+klMJvQ1IkHGx7V2malGNX9PT48ET69u3YY58+eqPtr4hnO0Zm1/puUbAVuzGRZQR4CcoKGmEG3ahN+T5AZ/3/TSyzqDuU4YQh0O21QQa4+0U9ob8Wjh7NreHAhG6xtaIDGvQYIk9oEZA8lN5Md+0aywVC+K3DbAfOXKZehYskjTuhRcMeOCNR1FMtk8z28TxjBbJBxg8DcnKwqIR8tRlssgl55EQ11c62hiKoeJTAh7j/QgEm9C//CYrIcGBntFUrJ+MJ955iZUSATC/Yifw2vF3mxoaFD2Wuw545WVEudx0on77VQyqetOcQyf7+Urlmn/53smyUsBk+RHXvWs6Reb/vFTR+ynee28xz3BYw/cstbjupWgin0KP9cJ4+QioOklm3TnNSWY7m1i/f7M68BzguQv75NsWNwUjgROLpvL287x2vr8Cr5uhsGzH+Y5YoS1kc/CM9xZKQuxYqGEDVC0QrBYU2BRE4PxunBf4RSbVPkSfzHPgDhIXtecn+Mnz7lOeH15LUS4sM7j3kscxuU48hxRHqAL+tXaluiA68mCxXkfOX3KvnRiqN/sn4p51Mbj6tHYC2fzRWWTnHvO2SjQcixHrIZrI4yR4WG9Pk5V9nT3IZcvw/D4FIqBCEYmphCMRJFkX8opGVki86gyAJX7KesZPsNk6dTPkuihMLOcYdo2UcHXr1qAWRxuyoa/W89rIlA++7o+ro8UKOvwKf4b93LVJY7kMkKj4CyKDFTXs+esxj3ZoIwUOhqUhzXJw3OX54UFYRs5wL1B+aScQFOoPScDkiY8oLWUJijYl3N/SJcm3rzYzt9TA8TZs9o5SrLKE/Yi0RwhJpeOnJ1NNrHqLIpEUDL4iFWZC213ziQ2PRPSdArPU2IZXPsS9RZhZBynKByZJWGtu4aqQWaD9lqdNq3myQ0jdY00lfDNgfbai5ytleWo2n0TVpTNav2qH+PUuvZKszASeavMjpkJmhmszsiDg8/OEBUrLmbda3kTwolczosPz+bP8v0L751qJgfu+ykaiQgDQHIqqR9FYYRwPl13+z+RReqVeZlnRB9ajz5v0AV02/UxPM/q3T+cCNG3C5AYNuLayCTrufTncgbdG5bma0l+T02ZuvqI74PvTd/ZWbn5+QmbcuY9MWG2zqDXiQq/jF7//X/KFVioEdSCHh4x1xwb82wyN0c39mRB2dbkKOCPD5ebIpD3nyxbTL3F7+VBfvnqKzvCRhi9PxsPavP2dDOCjrXkU+sVySUWwI/Yz2KT9eC6RlEqbOeX61XoGq11vqcG3sxY0Agkkm8emzdroO2wMEWCZy7Juno1rrd0siA3A129Ktpbj3CjM1bXRgr9xu6ben8Q+U2cf1c4F22DOPapJtDtN95/zvk6m4LAGF3eA1kuFBiYVq5Dkz/bij9Tg8lOwakkeUDpXZaZdYF5g9u4ugUumcp3OmeBqFbIE8iyJt17Jkox4gLPDLExUFgbJRtC/t90VoWj93bmBqwR6ADB4rTAtUuuv8nGYN3IKwMRqRxVOOAs8IxFqs+oUEAtFSTuPXH9RMvNX50HN6cFCCQQGG6d16og1GIhh8G+Przy0iaBNe0dS6TAJFERq6pGR8diqUCaW+swNWlEBZuHscmEGpHxxCQKOQuflAoym9WBYQeKkjikIubjwsKA3rZVtDgIlyGdHMfe117FGG0lclmUB+jFHjf1MZXHKqxyKvr5QbAvlTZLMY0rqiC2QowHPNeHinEqYKQksqKE95zEE/9c3dDggsIs0+PUqVM4sG+/1Bv1ddUq9Pj+gpEIyiO0fogpjJLTLryeXh3ANc6mgYWz1lcFGyreVwvaNLLQAioJMvmJHF4bKnr37d2HNWvXoGVeq1P0GCjrSUVTaxNoKmLVyvVoal6A6Wm+TwfzFalQyuuAp2UBrzeDHbtPnkBdXZ2CZwk2sGEzX2nLpRDo5sFErmfnfcxrwWmeoYHj2LrldyibzqAiGEFNdSPaFy1Ceawc44kJKT337DmArdt246xz/wKLV69HMp3FE4/+BNdfczUWL+7ALx75OZ579lmFxhVzfI2ln6hHgq9VKiL3Z6m0HJhlgJb5UXNv4DOgxoP7qrx+kphbV4n1q5dgXstc9Pf3CpAdHBrU/SSYx2d3UccClAUjqKubg1whiM3bd2Lf4S6EmSXCsHutKelJNVnx1re9DTe94xaUx6qUuWEe3VlEqfhJJnFw924c2L0Da1e0Y3zkNDJTkyKhX9mxC2NTKYQqGGiXxUD/EPr7hrC4vQ1LFs1HTbwCtXVVaGpuxXMvPI/xyUksaF+E2vpGHD95Cj2n+qQs/tBHPoxrb7wRv3/6WTz9+BPY9dprGJtKICdVHK+ZEamyp5F9CNXEBMHMdsPvswShVBSzEM9aiKbsA2ZNT3Bt0t/d7U6m1HVr9pZbb8UNN9+G9o6lqK2rx1Qyrf2sMhZBVUUYieFBHN6zHXt2b8funXuUeXC0uwd9owOappk7dz46OjpkIdfXN4B7770PZ569UQDDjm2viAyrrY7j3DduxB233op1a9dpMoX8scbxaUnhSCweD6yFJ1JpvPrqfpw40Y/lS9qxccMqERVc24eOHcWjj/4KTzzxW9kTkduVopLnLAPDZatoBJ3ft9ksqQFz4+1s7AlMG3lpzYKAA5F35hnMNcNzk+cR16oUzlQfFYsCWUlaXnLpZfiLi96Gjee8EeEw13RIr0kBlhVhxJkdwclGBDVRIYEBref6e7Fz16t46cXfC2BPJyZx+OBBAUjypeZUZoTh0g0Y6B+QtSGbcE5dkGwO0CdZ51wY1dWVmD+vBZ/73D9ibutc9PcOY/W6DUCoAl3dQxgjUdE3jCOdx3D2meslkFBQ8zRtr1Ja0yRYCB5V11SJqGCY5KRIsrAIkqGhAVRFq9BQW4t33XELUlP0yuf56dVvMxMVXjTha0HrbWx/XLduDa647DIFaathptuQgl+zuk7cF1rnzsOadesRq67R6+NzyylJBsFPkSQnoaT1D+zcsRNf+MIXkKPnd5bEZQiVMfr9puXHbs4QVB1X2JRbrMKAd6cCzhCAYn/LMGaC3wSrnVLXT1OIAFcIpOVqmcWZrTHWE9axz6j6pOAsPV/c3Bh4SjA/aQHgAondl7kQXTWQLhtA05o+q4ljRy5+xppM67pEVNRVYVF7u4KfSQDVcO24Rp7PLwlkTkJ60o7Nf0NjEwplYa2v6Zyds1lNYhmIQz3J6dP9+N793zdyQflIbhqPr0uqToJf5oNuYKYBTaaC+0OiQnUzyXtN1BIQsWwKs4mys5zTPzRt4r2S9ZZv6HWNWDfSHiODocE+U1jrHnBCmeeFBfD6CyqiwZ3DBmKYNZdNVJklDb+rVxHK9pRWNSKoeP+DAor4Zyp3F85fgGVLl8g7W7W6I4xYV06MTcgSjYCpgF4f5ul+hu8NPIDH18jag5lmlVUxqaCppOfaIlFB0EsTFS6g2ogKqjot/Jr2U9wLWH9Tpc3XMD4xpkmdqhgnJqwP4RRBRawCwYBNdSZOMuTXLLPsWrgMD6kpC6iIWritJpw5OapwV8uJ4/VhDWWWrTZZzXv6iX+4G9U1cfz8od9g365Deobfc/et6FjWhkd+/LjuwTU3XYq+3gF8+6s/UH3GGvWDH30XlixfhCd//ZyA+RtuuxJDAyP42he+p+/Rtmge7nzfDaoBv/hP37J7Ocvukl97y7uvwejIOL755fu1f4ciQXzoY+9G67xmPPLQb6X2Z6YD9+Gvf/G7bsI1iL/+1HtRUxvHT3/4a7y2fZ/WO4mIS696Mw4f6MR/fvNB/PUn34u6hlo89L2HcezgUbz7Q3eiY9ki/PanjwnQuvJmTnNM4Dv/z5dx0dsvxZsuuxjH9h/Ez7/3U3Sd6EYmX8S/3fdlTU3cfccncOk1F+FDH3sPXn1lFz75vz6Lquoq/MVFb8TH//ZuTYF8898ewN997kO6lg8/+Bts3bJL07rv/sCNWLp8EX7+0OPYtmW3JlPOesM6/OzHv8HWl3c5oYIte4KH0QrbH2nryoDh6WwO/X19NomOIo51Hcc0bUE4jVNXh3M2nqN91Lzp2RPaVDzz7AhSiaB14KmJ8gLIpo0A3fTSJmRJ8MriifueTR5EY5UYHh1FOUGuHAlsAwy5X/pcg1KN59TG3FN1zjrbVF87C0gMs4+x/jSXZw7ZUixcON8IZU4us3+IhDTFwdqI9lsi/QhkBqYRKuYRmM6gIU7brhQCnPDksU6LKDBHIITnXt6JeYtWYHBsQhNak1OTCugW0O0sZ0mks2+z6ZNyPW/MZ2DPyGtFooLCE6r1VSM4EQnPWX1OrALLli3TnymiY1/MXELWHJ404PWJVsQsd1Dh9TNK4ZmJJhNA8TlR3+5EbRIeOjVxCQA17M6AUCdqtDwuywMQAW2Ft2XAOMsl/ixOhpglW0H9EPNBRBqQtNIeYWcQrwkBVU426HwMsFfldFfM8g2YN5BJi9Qh6SYwm0pzkqC06yojQWJWiJqYjMeRcrWXLKwddqH8E+c4wbXKWoE/l6+bwCrrIgHvzmbHchwyZukjDZLtZV7xJQW8m8TIZlMIM28il0J6coLIKbKpjCYqKGjIqn+XJxaa6uIKaY/FIgiFA9r3a2prUdvUhIFT/UhmiugfmEC2EEI6X0QilUHK5UewPsiz/59l0SQClpaCJHu8vVcuI5CeokJv+S0Bm3Px4L1Xpov2RD6zlifA54zXmhiTZZyYTZk/SyRW8mIKlrp0BnW2Pd5ezGNBurvOBs9sgExsyi9iL67Q7bwRjSZwsLOdQl3WdGZ1ZdPbvHb8fK5VPtOGk5lgTfk6HsJ2jiQGorvK0eU2sSa0a2B4mp/qUJ1MLMbdSw9c2x7jMSsvBKF1pdkcsfbzpJ6fZuLrsfwGCxv3zxPfO8WosuDmBI+b6BSJNEtkaPuV4Vy819ozGQyeTmvPtMknI//44f8sUYbrVfxUuV6Lcxfwn+eJEL5n1of7n5rJqFjxtiFHZFnf77Nf9Ll+OpVCRZcB4XEsvnfL1rTanK/fnEVMgOP3lz/AdNUTWY0sAal7L34/BiOQ8QAAIABJREFUsjNh1hSXs4Qy0bWzF/PWpnyWnS2anwTyWTf23Lr8NoWVs4b2bjA2+Wf5bm4NzbQfs16uz0Bk70YBSss5M0ZQf/CuXv/L61fgv+cVWOwKEgFsDlAjCGSWE6YS94ueeyuLBRYh3ERZkPiAKvnuuY2TD5Y/UAl0ZGb5+nOzEBngVC2eFJCSlo2FaxjYEAmck/echT8qF8EBK149ywdbr6cUNmPBoAGBng5UlbuKFS8eCPab5GwWVp/vVH3a3Nw4mxVBdnBwU5Qnd8BAf/86+H+ezfWssvd/9hukf69eMeA3Kb4HKUPc2PFsZZoP7DJlysxoJ09nWhI4i1azr3LXVgeqgHUDhD1Tzu/Fhp3qfQsv8rYDdkgTWPJjkF61wUKZYBT/n4UR1Ut8/3wP8tp01ixSozCEkvr06ZyaA9llMVxbn5N3f57GZTfc5KZJgvJIpWcyD0ivnPBqPpElVARL5WfMvALWXciUVyjz75VxKm5YQJdLeUk7Byo8B/pPYeuml1DIFrBoMYkKN1FRGUfHkiUCYFrnN2vMXWHakQpMMIw8n5VHLzMqpCx1Ck6vPNV7cgVsPu/D0sjQh1EeCSKXSeLQnu3o7zmKMga2BWLKxSiUcVw6hMpolRRMeo9sjGkpQCucWd6OfqKG99WPXFNVyb9zvfk1R7KC9zteV6uDnP/P0eBjR4/hxPHjqK+tRZ1snxjISyCL4Zq0YrCpiXSWqn0e3AZ+EOgg8MN1Eq6ISInIe+D9NKVgcGFe9L1mQakRUJIZBFgPHdQ9P/ucsxAlsCBloz1dsuwgQE+FDsrQMmc+lixZhXyBhztfuxWC9PVHsCiVC611Bnp7cWDPHk2BbNx4rtT32Qy9TrU7oBCwoHYqaEsfjqyQmimTwmSiHzu2bkJypB9VYQZwVmLBwg7UNTTKNowKuJGRcew/dAwbNp6P5vkd6Dk9gF/97EFce/VVWNS2AF/60hfRe6pHajZadUix4XTUXiUiP3enurLsGNtbvfpYqmL+XaAfm+icVOihacYCp/HGjSvQWBdHpCIkb/CR0VGkprKYmqRSp4jmefVoqm9CvKoeFdFqbH9tH/bToomNTL4o8I/7HBtbNoU1NbW48cabcMlllyFcEUVlTRxJkmLTBdTGKpEan8CxQ/uQSQ5gZOgk8qkUTp8exGs79qEQBHKFtFRTp08PoPf0ADra2rBowVw01sVQE49iTtsSvPTyyzhx4iTmtrYKOOQ937N3LxLpabQtWoK77noPvn//D7Dl5c16XbLCoypIgKkBAQTibM2HUBbkHmYwJ8M/uS4VEkcASmSxedLLV13WNjPBp6EKU8aoGC8FdRbxkY99DOdf+FZ0LOpAfXWdGnmta06XVcZQWREB0lN47olf4dCeXegd6MW2ffuxt7MTi9oX4aK3XISqeA3mti7AseMn8ZOf/hwXvPlCLFnSgdN93SKwkpPjaJ3TgAvOOxerVizD4o4OLFzULpsFqpk4HcAbREqNzwzVm6/sOoKuk4NY2t6GjetWIZfL4MWXX8GPHnoI27ZtU+NheT6lrlzPu2x63Lqabd0j4YDOPMuREWBAIJXkPJ9ukc/0NabFFv+N4gI75zO6xga08ozmns9vRhvBa99xE6644hq0zmtHRSwu4Gh0YkT7Pv2t6eGt8W9ZL5q1IUHPkyd68NSTT+DQ3p2oCBRw5MB+OwtoqsS9scKIismxcb1mTk1RxT08Poa0QBeTwEcjZWhqqMXVV12Bv/pff4V4dQPlsMgggs6TVH1Po7evH8e6DmLDmRv0WsxCsiDPcYJqUjVm0wLMqCi1XIiUgJn+/gH0D5xGTVUN4hVxfOA9tyGV7EcgkHFtpgfQ/1ytZ/eIhPCb3/xmnH/++foZnpDh9acal/eA++vChe3KNSFQwD2BanZdt2kqM02Vx3VN4PBzn/ucrEg8cadGV/fVhS266VLaNbKx5nkicI25BdNUoqZlvcCzQdN4bpJmRmxhQI72KtphcE93TRJ/lvn88zJY7of/8GSFnlROiOVtooKv2ZNnaliN7ygp3Hxjqe/NyTPX1LMds/dmBAdfQ7y2GsuXr8Da1au1Tiorq3TmyAM8l8GcFk4LMlzWRBW8tsqt4OcQHGEeArOuNFHBegRIZwo41nkCP/3Zz8xigfWVUwsK4pdQI2+TXWVWF6UoXGBzHXbWAZLxGCFMkFl0R8iU+vbLrB4JxlktagSHgBNv8WndvO55oZgXADsyPIA8ySieUQTGeG28qMfZnvjrRkJDoJxTKPJn+PrR15ule+UUhn4fCVXEBEjwvXGdLlmyGPPmL7DvxxDxaWbQlSMxRjvEUVRWsv7K6Fpxj/YNfilAUveS77FMRMXY2GiJqKAq2UJraedp+RQiRmf5uvN7EhjlnmwZFQERFVyXzB9jvU1w1cRIkNVelJZzZeWysZzs7C9lrOkc0bnLZt/1MLwPJCU4IeSEDgTLCXxJ2clnMEeveIKV9px+4jN3S1H90P2/xInOHn3uLe+8FuvPXIVf/OQJNHGvf+u5eGXTDjz60yds2risDBdf/he49KoLsWvbPhw52Ikbbr0SJ4+fwn987UEH8gTwqX+8W7fi//3sN1QvWE9kE9eLl7Xhlruu06TEt7/yA6ubpqdx/c2XY+N5Z+D3T23C0YNduP29N+hz7v36j3Rtlyxvx213XS9y5Cv/cq+rs4D2xQvxrg/cpOtOYuSq69+K8y7YiGcffw5H9h/GnR+8Xdf9/i//B+a0NuOG990mcchXPv05vOcTf42VG9ZhyzMv4KWnXlD+zWu79+G7v/iuvt/ffOAevP8j78RFl7wJD//o17j/P36sHLSOxW34u3/6iF73v37+O/jkPR9Ur/b9ex9G17Fuvbbb3n0NzjpnHX7+4ON4/nebcdcHbsaGjWvw4/sfFVFhoG9QwCFrYNVchWmUsy/N5dFz/KSeM9aXk8kkegf6wTvHrCySU6tXr0RL8xyRpyS7zbnOakYTAhlIpH7V2/TkaOsTxqZNm93ErvWNXNcUVFBUNEkSXZYotk5Ye3KCx09Fz7aA0bMqqzrRYAKTlP+Xo7iJ+6l55BuwlsHiJe3o6GjDVCqJmniliGn2UpxuJrbow39JGATyWUQjAU1UxIJFBWtPZ5PavyoqKpErhDCamMaLW3Zj0fK16Dx5Ss8vMySYWcfezuYEHdBaoE1eSpNM7BV5HVijEFxnT8GJP28nyXvBfoLVDEUFnG5avnyZqcLDDBLOOIvBmVrMLJ9MYczPITFAEJ4EAteG7+98iLJem7s2Ihmd6NArsS242gDskvWLsAQDkJWx6PJPLHPJ9l4WQbJQDhnJwiJQ1kp0fpjiPhM3N4A832O5shb580nqcm/wJIrEXSRCSbrIecEBm5qWs8ktli+q34RnGLCrLBPle9B6yXAVri0BtlKe2+v0Z6EyIt0e4IWKynUIMl+TGZMu/0NriL284TdcMDZ5ApQV04iGAliycAESw8PaC+kcQNvJ4fFxWTtXEixPT6GMVsJcSwXr33necoJtZDQjF4JguArZ6RCGxiZRCASRFGbEXjki+8OKypgEAKwjZcVHmyXVXnYPeb2q62rROm+eXX93vVS3z9oH/bNpz7izEXKB2IaHGAnmn1/hN24t6D5rYsphNayZXV6dJ7D4fZV7w+lHTUtldB5rEoS2m8mUelizMjKLMsuksfVl9aWRVcKIHInH1+aJBhNe+GlIs9z0WQu8pzadYKSIXq8jAfU9uEeQSMqSAKNNma0LZf6ELafSyALb17iejbwhZmXck027esU/2y4Dv72olc8ShQ8ULGoSh5O4tI11od5+YkEkAid0Xc6pdg2XX+onkES0uSmM0r7qrI98Pghfr9/vTDRs9nf+7PN4Ga/fwWcbS7XmiouHHGDPusTEx39Q28j5xdxeWHMJh3NrhffHpliNwDSBrZGRfxLUL7Vb3lrJ/QN7Gzfhb1iJW28uO0NkocugknMCcQ8J8ox8tWxdKxuNPMrrdfh7ppqtVCq7deNyLkpk1x+3Hy53RWQQ39PrRMWfa9Be//f/rldgEcf1HIPnfeQEToABu2kpKKyXcoeBQDZrtnTgOD9BNaou/NhUw1RmOf9XFiRUkrqJCx4G3m/RyAdTIHi2kYc/izkVAG4cTlMabhzbb5RGiEwjnbNDnCFhViBlkU6mZ3yAuZ34EEd7oeqcbQyNIIRt6H5agluXxmE5BqiAPSuqbGrPDhmrn8wjnM2Qik5ng6MGTMFnLryIBYMriqXYUfC2TZ14EFPfRxu6eW+aTYMFXOlg1EikY5JdpkQ6RVVMVUkVY+pkY5f5elnE+UAvHuSyrcrZz1bGAT+Hh5or1Fmo8DXLG5OqTnmR0teRMXsF/bumM+Rx6tQETGrI5hCrjCGZTqoQ54FL0qD052kCbQTNaFGSxRU33azCgq+Ho9Whcnrg21ryxZmuswtCJshAz26uAamOXMAhr51n0+M1VQK/aH9FUJEKPKry+/t6sPWll1DMFUVUNJOoAMM2a9He0aHX0NLaKOsnERXlFZicSuk6jY6PIZ+1MTx+ngBDZyVgxca0+3cWAVYwV0QZlhlCPpPC4b070N99mOgfKspiCDEgHVTGlSEaYQZETPefxE95Jb1sp8zbe1ZIp99XWAjw2vP9ichxzxvXNV8fi5tKWrAIZLR1fejgIZEVNXGqhzk9wYmKqFun5YhFTb2czEypQffgCkNyOTbK10UANxBmEe0UJVS2sRnXNBILfQu75oHPNVHIFzA8PIQ9u1/D+Rech3nz6R/O0XZOEFghxU9W0VAIaKph+Yo1CASobOLzYvY0IioCBYWjkxTo7urCi88/p2bmbZdciXh1PXKZohQ6Io3KvPfsH+7EBlRPI52l8ngEe3duxWB3J2JhC7WdO2+hfqUyU7pm1dV1CJXH0DBnASbTBezdfwSPPvwj3Hzj9bI1+c53voV0KuHyE2aICtsjDYjyRSkBEb8nlBRoTn0ToOKFxVQgI4uyMMKIsllJjuANZy1Hcw19txmAGlAw9fDQGMbGEkilsswORnNDM2qq6hGrrMGBzhPo6huQkz4nLfg8Grk6A5q1ty/Ce9/3fqxetxbVdTUCvmQLR9CmCIwN9eHY4e040bUfoWIR3cdP4+jRkwhGgphIjgqYPnGyF4MDI+hob0Pb3GY01RPcD6F95Vps274DBw8dlg3A/AULMX/+Qpzs6cbeQ53IZKbV+B0/fsIppAzAJjBEdbd54nNay8hTG6cmqWXENG1xNEHjiVenuFZIbpLqbSNd9J75XCj42pRo/vzgM/GPn/0s1p51tuxj6nifqbjO5pDkpBcB0WgU8XAZXnz81+jpPIyu7i68dvgwXt2/H3PmzMWVl1+O5jmtqK6tx/ade3Dg4FGce9752HD2WWiZNwcPPnA/fv/0UwhM55FNTSJSFkB7exvWrluD8990vrIVmprqXTivWRwmp3J4dc8xdJ8exaL5C9DW0ohnnn4SD/7kpzjcZRkYJYJr1tLm+2Rj5a2b/OfM2PVY4e8bmdlTF3xWqdLk+c7fqczk92KBT9sFNX20E1SAqPnKstlrap2DG268GW+9+ErMb1ssUjiZSWGK159KJTfV55sO/9ppK7v15c149qnfoJBKYGxoAD09J5GlslpNX5kAaK5bEsYETdnUDIwMYyKVRDDA85A+x7QSi2BxRzs+8w+fwdlnvQHTnFQoq8CJnkmMjE+jt78fXccPKajaCwrYr9ILncpjgieeqCD4EglHnWd2Bfr6+tDXfxrVVdWoq6zFB997JxKTPUDAVLMyf1QC45/7sHDLdevW4eKL34q2trYZW7ysAfhsVKIVlfq8lpa5Uv0WpOS3MXPBldzTBGST2MjgxRdfwFe/+lWXNeVyedy+x25UTbNTvfEs1X4sgYk1Utz/eIbmMwY6aHLC5V/5s8ar5vh1JDs80CvfXFeLmIcuQwSdVacDRUqWVyQLSRbncphITJZAUt+YmbjCGjtfdHGtGDHmFGoiNWY+h/8Xq4ljxcqVWL92neyJqqviTgU8hXwmrSwYTo5RnCJyNhpDc/McFDlJxIkrWsVlqCBNm6qTIcl5YM++Q/jlr39tY/ecLisFIPvag1/rrRMIYBGcpGLTakUjWAMIulB51kg5Ba7b/5mqn3WsiQcCHK3yINqsKSj5mmu/tukPTh5l08zCCKFcmSFGVPiV5xtSD1BYyLsjTbiGFIxqNa9NQc/K/3BLV00vrWxUexm51djUhBXLl8sClc8cLRWDZREkxsYxPk7SgfZaGYEaIir+yJfZyBNHVJw+jbGxEYkjKGIxooIgygxR4fcmP50cQMjsXzIZDPQP6rWTqOD7pAKc9RGJCs+3kKigips1Deu25MlRyzIQ4WZ+8jxHSNbJmiNouWq09Mplp7XP0E6Itapqf6dWpDKaNT/rGU9U/PC+n+Pk8dO6ptfdfBnWn7UaP3/wMSxd0YEzz1mH3z35En7769+L+CUAue7MFbjhliuxa/t+HD/WjWtvvkw5F//5jYdcrlYBf/u5D+me/p+//4oCw0tBrQAWL2vHbe+7HgN9w/jml74vUp+A3nU3Xo4LLz0fm1/YjsMHjinHglkX3/q3+7WGzjnvDNxw61Xo6jyJr3/hPv0b62a+v7/9p7/S8/9/Pv1lkQM33nE1TnaexPEjXbj47Rdj3449ePaRxzG/bT6uuvMGjI2M4huf/Wfc9qH3Y8WGdXj8x49gz/Y9yhJ55ZUduPdn96p/uPuOT+KTn/sw3nLx+X9yYxwfm8T3/+Oneq2s3x564Nc4sPeIasB3vu9GbDhrNR75yW+xY+seXH/L5TjznDX45cO0i3pF14fnEJ9jA8ZDOiMaa2uQnUqjr+eUiKfR8QkEwmF0dZ/ANAU3FfTWT2hC7/xzz1Mwc4ZnVSIhG1r2TQScTeRjkxIWGmth9Px98+YtIhdYI9iUJzMk0tpfZBdX6scMeCPYaCIqU/ELZHa/e7KMfQKFCGaHzDqFv9v0v/38LBa2zcOy5Yv1bE4xO40kHK3X4nHkmQvlfPKZu8dcoHg0LKuemmgY9fEKZJKW58J7ns4FMJkO4PebdmL5mrPQOzisfW5oZBALFszXNeI9tKByIyZ45hjwmENDfYMscPkMSilOW1gJy8owMTGuf6+tq8HY+JiU98z9k8hQ1qdGBkwmJksT/Hw2mRfF98TajGIHfvDvPHNodSSgz2WS8LrK5kWTBq73dqtMdlr0fHdBusQXvJ0N+0lON3ACmfsG7xmfTX6+ahxzQXX2l+Xqcf1ZmE5lVDvIYlP3M2fWyuyreIZzsofh6K7/5z5DvICiOxHaGZu80/5sykg3YWe2nMQKfI9O0JNnPcVNfl+33temXv0kCjEH1lcGLhuZyT2O95m1l02rmxpA5IcTPzLHkfd3amIMTfVV6O48gkAui8pIGDVVVaiurUVNQ6PyGHv7+3DG2jWoqYwik5wC8YXE1JjeMy352GN2HT+FVKaIRLKAVBZIZguyfOX+y+vKvY+kcmV1XJOenDphPcOcxDBt+dx1TGYzqIxXyuGAYgKzvbManrWoJpNc4WDnisOC3BSn2Q+rC3bY1Ky14awjbUiNdlIz/bKfqOO9FLlTKJYmVfjdbIrFLHr85ICRYDMTArLpi9hEET+P95KEt+Yihb0YVsX3JfGt2ALngkHCw+Fn3tLWcomsv2EH48k8nlUkSoyMIqFh4l2tS9YKLkuK54a3DNTUojAdC5z2YgU7M83Kie/ZLKzYs5uTCMkQ7gseW+D6488T2O4AcC+wFU4ogZSJSvgc8yylm4LHY7zoeYZIceQIhVGuvtPkt4Z4DN8yAtSEzNqXAwHs+W1N6UzhRIVf1xJ+aP80goX7hc7eWNSuoyz2iDtYvVzC22QV5wlBq7m8oPiPDy+f/eEJB5u8dHWYIzpMVOvqN4cN8r7Y3jdzz719vT27NmnDD+0t7u9eCG2r2v7fnyH2MxzJ8Ucv1Nd+JvwIvE5U/Bcd2uv/9d/0CrROm3JVhYADe9SS04MxnSop77znGzceFozyMXYEQ4mW5KZD1R6JhpCpSwR6kA13oInAe7G2xrwKoFcwoI1pWq7BtAvgi2p8TTZPtsc6n0kbo+QDbgCLAfwiKJiPwDAaNoizWFex+rMUtlItcKy+FDLKA4IHpGUryGpHnrUMiDLwxjYeU27ww28wOvS4ATvyQ+AYy3mXUWE+ubbpqCEt2kbsVRL8vlSVyDfXhfzY4WAFiDYgV/SWRvq5KTMYN2eenQQIabdA1Y2fZhFoykY/yhyCgggdhSK5wCDvRcxCiffLDhdTgliDGZVvOD9PLLs88+xQEyggK6eisxAJqECjKtCKCKrbOd5vh49ZBjDjII+3XXudFfahkHIrGL7lFWPej1HAmiPBZhMVVkyQ+Z9RgPJ+1NTVmJ90ICSiYmJyXP7mfb09eHXTHxIV08UAamvrsaC9XSDAnLkNSCdp21Jr7zkxM1FBokIKVY6hujVshwzfuZEtzLFQSBJ9QCvCiJQHUcilpSDuP3kIxXQW0WAlylgAFTgODJSHLayaa4KKjYALCjSg0QdeWQioV00L+BM27kAIN3YpsoPBtLGoSCdPCh47ehRHjxxBNQvS6ko1+cyo4DPI60RlKomGZCYp5QzXM4tfKqN5Hfjeqqrj5ofPMDE30UMwRWufa5rvmSopqkm4tvJmQ7Nr53ZU1VRi4znnCEjgOiRA5EEuU54R3Ixh9ZozECmnbRGbBSq5ieZMa0oiGGGY6zR6urrwzFNPqoi5+G2XY8HCReDSyjnVMSdVZMblQky5Trz6WARqNo1UehxH9u9C95F9qAxbM9rY3CLFP9ctn7Pa2gY0z50PRCpxenAC+w8cxRO//Bluu+Um7H5tB554/Dea1IE8tR0w7ohQP5HC96Xn3REVmmBRkKOBx3q2CaRIwWXK9rJiCBUBjkiPYdWSuVg5vxUVTKvmaH9FOYaGRzAyPonhkXF9PUNGy8srEYlUondoFH2jY5ig6qoiJp96I5YJVBmAxfv5pgsuwO133ImFbQs1du2nZKi+y0xN4LXtz+PQwR1gQkL38V4MD09iKp1AWYSKwHIcOHgMickUFrS2YkFLI+a11CESLGDZ6nU4cuwY9h88JKusltZ5UjTH4jXYtnM3jhzpUnOqZ54EDac9uM+yMSmzYpOgd0V51E158TfaGxigyrqb682aDBdmZuiegIPJiUkpCKWOoXIoYDZjfCZ4zbkO6HH8pS99CQsWdaCmuhrxGPNcogJzJ1NJ5ArTqCgLIpzP4pXfPYnsxCiOdx/H7sOHsWnnLinPbrrpRqxduwHxmjoMDI/RDBQNjc1omb8AdU0NGOjrxTe//jUc2L1LVgxTEwxpZiNfLSuHSy65GDfccC3mtjQZWQFaEhWw60A3untHMae2Dkf2vYaf/uTHONzVhXTe/KL9fi6wsxRya/Y8XgXv/92mLGwySg2WI8ZERqvQNeWubOQyaeUJpVNJNYpscgTa0As5Z2P4tILxln/hWBnmzV+ISy69GtdcdzNa5i6UdzefQT59PA94zf115/2ycMegFNK/+sXDOHHsELLJBE50dWJ8fEznJM+GpqYmTYONjoyosaWiM5FKYXBsRN799FFnZkl5Oe31orj+hhvw4Q9/WMq9QjiGru4JjIwX0dc/gBMnjyiQlPuqPorM1EjK+okgDC266OteFa9CeZj2F7af9fX1Y2CoD7XxWkTLynH3+9+FdKr3/zdRwbORQfFXX/12WYTxXiifgIRZoaifTdCwurpGk3sEy3QUM+y1MC2wUnYBLmuBe//o6Ai+853vYOvWraX9w+8hurfOr5v3mveJ02/am7U3OfW+C+nOZ2ar2M0ixxSg5u3MrxPg4TLBRCA6kFtnkkgFAz19Qeb3WJ3b3ENd/glVuF4AY7XPTPPFv0ucUgLx/ITCTGPmGzmux2hlJVauWoUzN2wQUcG9j9eW052FXAYNjfUiKhQcXpqoIFFhimeFlHMyM2UTWARU6LO9c+duPPH0U1aHUe0vxsWIHas9ciKkBRIwNFXWjGb5KCBN5yVtN0mysn7NI1dmpKrI1j8iKgjwaqLJTUH5hlRWBSopplHIk6gYQio5qSknhb0GIyiWArVnVKQGYlkQb4kgl3LS6gO/X3gxTKnpdSrC6cBMhhKvJ/dIeobT4pCkAs9y5khNjoyKqKiKVwhI5dnFX14JWbpX/x9EBYOm2WPwHmmPcUIdT1SQYa4U0MBJ2H6dXQSY+UERTCIxqbrUGvaibPVirGnKqzQFlOgcRCRs618TYS5wXH0DVams0dyUTnHaAD27NgY+WKC3iSi4xAlwkaig7c1D9z+qyQje41vfdT3Wn7VK1k/NLQ244KI3YvOL2xWe7a3BLrnyzXjrpW/CtldeQ+eRk8qoIFHx7a884AiuIj7xmQ/qufjC575Zsqnl80bgacGiVtx613WyWqT1E7PXCBQT7N/4xvV49smXcPTQcdzx3uvR3zuEf//X7+qer1yzDLfddS2GBkdlByXAKliG+W1zcddfvkN70Bc++3WB5R/9u7tRV1+LnhPdWLx8MZ76+W9wcMduLFm3Cpe6MO1//8znceuHP4gV69fhhcefwsvPvITp6QC2bNmOe39xn+7h+2/+KD7693fj4svfjB/f/wi6T/Ro8pX9QmNjg6ZkNr+8Dff889+ItOJEBYkKbgDv+cAtOOOslXjw+49i3+4juOamt+Gcc8/Azx96Apuee7VkdyuRVpHZBUHk0yn0dncjm0wjotxETu3nNS3a2dNN1BS5IgGpgkBu3r+G+nrMnz8PjU2NIqp4do6NjpaIfu1HtMJT4GwEBKu3bHlFZykJdU7g8Fln0DTXF88tkl/aC42pRT7ngSRT685YEdin8HuZYMtyEqTHYT1E3ZuzNy8ih/nz52LFyqUmHEjTdpD9mZHRfLbdZqocKO65lZH2X3PLAAAgAElEQVQy1Rs1FSFkJkck7KljKHkgKKIikQni1Z0HMWf+Yhw81qX8HlqhEnwmgcvnuKa6VnlofOaGhoZ135TrErJJb9rWkuQxAV9K71cZhrTCDZWpT+TUaFt7m+oVP+nH/6PAygsqrFeetlBiZ5tVcmAogc82WcTvTQKD65rPlWoaB/QRm+DP5z5tpKQBBAJprfg2kl6Ttxmrb5x6nQIr1iw26W/9Ei35vFjRbAutf+f3lT2WbPisBo1FmelhQcciXtIpAfA63519js5Vt9+Y/SJtninWdFMSznee91giTQ+uO6GO9lb2/6pfScDYNAHXFPdOAcLejkih3zaJ4dXqmqrlN3XXg7XTdDaBuqoKpGkrOZVAaiqFZDKPLMmvaACJZAaRYBFNtAkuj2BOcwOqayvVy7O/rq1vQH/vIAaHJpFIFTCRyGEqO43RyQRyzkZIWUFTU6isrhKZR3yGVn4hvo+8iRh0bYrTqK2vk6WULK9oZeZshkwwZ8JY1TjCWkz0STDdwGIjgHwvbuffjA2qF0AIe3GZF6xtuB9IqMF7KStly6fgWW/2Tdw3Zix9bN8x0JjvxZMpvobx9uKmL3H5DE7I4R0rSkC/KV3V33oMie+PWQv8XNbN7Mm09nM54TY2vRESluJdQZRDMSvA2U/asI72hN5s0kvAuZuSFsHB2t5Nskrg5K+p+JSZCQd9DwofXHaFsmci5aV9UhOoBP2dOMDXgtrb6Gzgpjz8pIRIOk3T27qWkMAJoPm7MhtcIDe/hgTZ0RfmlpBVTlTwpVimC2szm2LifmJCYhJdJE4Mo2Q/XlpHjgTzUw2yyHW5VH9qpsI7qth5YBOxZtVpeVYlG+xZdZlcJVzOlc4Dl+MhMsQ5tMgOzom2fSC3uZhYrzbbUso7vPjr6CfL/hTUzPddIoVen6j4b4rGv/6y/+wVWOJGn2csj2wU1k8m6PB3bLLG/8nsO1bcmluSEAXz0HMen6buNEWAAF53CKt5c8CZATAWyiPwyY3gUkFshzzV8c7vXV6WtoGSgLDwGAP8ZsAbN4ngwsxU/HnlnlPpzYzfmfUGv7+p0mbGzrhpsXjzh54f7dJYp3WWNmrMn0+QhUUsbQPcv/sLbapgAwn9BIYx7nZt+D1kp0RCxykg/PX7g5sluy3bjP2Gb42dFVrRCgPj9NJ0PWg9EZM6xpTI9Pmv0MaeymbEOPPA5dcQCKEnNl8Hva79hq9DoEBP36i9PykhzHKFartEckoWPzwY/b0w26ppeZJqmkK2OEURFfTDtxFXvoccLr3+BhsPjkRU+NO/m+/Jg2v+/bNw4cFGooK2GD6EyPsLelCf16W6tlo/l++5o2ORlEIEeXtPG1ERmC6iffESNDW30HQFNSQqqHilP3pTrZQpDXUNAtVp/URrHKpCMykLfvNEhbdY8RMVPHTIwehQCgUUHFkeDSOXmsKRfTs1UVFMZ1AZrhbYmytkECgrIBKiZzOtYMKg1y1XE98X76EHuPhz+Xd+bzYL/EVbJq/u8Gp9riVOE5VXWlirDr5CASdPnMCe3Xtk3ybrp6qYmjp+X4KHbCC55tLZFKaLMxNBVFGy4GSDF6O60BUz8uAkQE/SQiregkgreurzNYmkdLZuzJPYd3AvLrzwQjQ3t0iFWXAZFDOFFVUPFVi6bLUmJALguiSQbSPyxTIGYEYEUI7092PTiy/InuXNb3krFnUss4kK9xzycwUhSQ1ne8EfEBUMGcwncfLoARzdux3RoAGkBJ3bFy816wcSfpU1mDN3PoLRapw4NYwDh47hmd/+Cnfc8g488vOHsX/fHkjB6r3+/YCWii63hjVyS/DN9hev7vfPKH9Xg8rCOmAFaKAQRJhK2PwUWptjOHv5EsxprMfE6BBqG+vkAUs1XG8/QSwLuuf0B4HDyVQW/aOjGEtMIRyrwkRiygFVtt8a/laG6ppa3H77Hbj8isvR2NBouR5Sbk1jOjuFfTtfxoH92zExOoz+nkF0dw8AoSIq41GwB9+z9xCymWn593csmIsFc+tRhhyWrVyFwZFhdB4/idO9A4jFqzW5FCmPYe+Bw+jpOe3AKWcPSAsFjhCzoeU+JlI3LKJCBJn2RoJFzEhgEW8hdda4WDNKgkyTbFThTyY0Vu49S13mbAkk5n1dvHgxvv3tbylkeGJiEtPZvKx3OMbOa5vlfkelVC6Lbc8/jeTwIE739mB/Zyeef3Ubenp7cdVVV+Git16K5jlz0dTSipPdvZqKqa5vRDROG6EwnvrNr/GD796LaT5TVNZlUgiXc0qtSoH2111zJe6481ZZOvDcSGcDOHR8CEe6+tF38iQe+9lDOHhwP6YIIARs6sKvG52nLk/IN2IEDrz3Lv+PTY+F73JSJai9k4eALHqkFmWjxOtPUjEv0IFTKXyuSbQSGFVDqGfZRv75i0hKJErsI4S29qW46uobcN31t6C8ohokfotBa0L4wabTTyLqCA6EMDk+ia7OI/jNrx6RPVb38U70nepWYc99jwr4aHk5JsbGtHfHae9THlFOEEnGcJAgBe0SIgIN2trm4+N/81Gc/+bzkQ/GcLI3hbFx4NTpPnT3dMryQyP7Gv/n9FBGlhaaWstYTpO3fiKJxmaQGRXDI4Oojddg6PQg/vHTn0A+NwSUZTSFZ5JrI6lnfxhxbGeYBY9fov2Yzz6bTz6r3Pt5PXl/amtoA2akHNV7Y5PjAjpqq6sFWKWmpmSzwfN5//59+N73vofR0VGnXqPQwAgrAypIHthEBolnTUSwUXRWSzyzeX5ICZo19Z9vUv1amq1sV1ig1GJmV2eAu9mMGUFhNm2+5vB7LdcVATLLjMlLgMC9ZeaKeYsiW4vWbNuHX8u+gfXAgK8HYvFKrFixQn7zTY1NqInH9dpo1ceJCip6Oe3JdS0VZ8yUmmCuBC0oc6wjjKjgRAXrndx0EC+/vAXPvfii6j0pJN3rMUEASQOz3mKgNe8HCSRzefI2pEawmn2LAVO5gDWlfpLCAq6dVD/gg1hniB6dU2JXGZKZk63N+NgIEhNjFoAaCSMULucFm1XjOZWupo55/cw7W6pC+VLbz/NggK1P9xq81zIb6QCnPy1jyk/ZEDhauXI55jLLi+dGMaSJCk5HxCrZUHMPN6syZYw43evMfWSPEMDp3l59jc+cYQg19xauXYJ9/DV73fHfbZKzAvksJ2FJVHDislrvhUSFfPBpz+eeQdq3MYuBZKPudc+41gAnSrgva7IlaJkr/Prq6ir1LhRakFzidBXFSeotlA9A8cHMNA+B8U/e8yHla/zkgV/hyIFOfd4t77zGrJ9++lu9h+vecTn6+wbx3W89JIUq18y7//IWLFuxCE8+9hymEilc845LNaX4ra884O5NGT5xz1/q6n3x898233DlZhiIZNZP12J0eBxf++J3S6KlD37kTrTOm4NfPvwkhgZHcPt7SFQMKlxb/Vg4hI/87/fpujALYv+uwzpfL7zkPFz69jfj0P5j+M5XvodYRTkuefuFOO8tb9T+MDIwhIe+dT8KuaxIi8tuu0GTC1/+3/+At99+C8679G04tu8AHvnuQ6qxBkZG8ZkvfVaq9Q+/61O49rarcNtdN+Ll57fiC//0dfUZ3Gsvvuwt6h9OdJ3Cpz//Yd3fH373ERw5fNwmKt5zAzacvUbXd/sru3HLO6/Gmcyo+NFj2LJpp6maNRHGvIQw0skEGBxXE4uhmM2j88gRJBIpxKriqG+eg4OdnchSCKHs3xCqa6qVtUEwedXqVVi4cAFG/i97bx5l+VmWiz57rr13zXN1Vc9Dku50Z+hMJMyDiCDEgMho8ICCoAg4oOjVJehBr8fjcrpeFJxBDyIgkyEEggTI0J2kO+l0ekxX1zxPu2rPw13P877frkqAdf+WlWaF7nSqau/9+32/73vf95kWFrX/c4HzPZiNkNvl0pInmVaN8OCDBIeNec11lYhbTpyY7NxT1fOa13vINnCss6nOb9rukhAoZjXXuavxdTbx2TS7NlP21DE8MqicCuU71A1cYz/FmpyECdZCsoChjR3VGdE6WlMxy6io5AVeEHzmGRNLZDE2s4pjJ85ieOcBTC8sqR/nGUjrpw0/E3lfmItF8Hxubg7d3T1iSFPFwWskxQUJYnxO46YgUc6cArczsnnr6e1B/2C/e+Dza1wN6rZaFqjtmWRU11ftM2nvdFtCWgQTJQy5eyQeWq5FWkPbrRmSfJBCiKz42j6otnPD7Lq4h0g1ns/jyDXX4PLlUSwsLQmo4LpnL2RABG11LP+R9qlSkJSN8KOzQWvAAq35M7kOeMbLflTZXm7nJ7DT/+fEHDLqFYAsC0XafW5YKDdBeFrdef4fzxFje1PBbkPb0P+J5OPZF/xvrJP5u7KTqhYkzrOYtUbId5ANsBP+tI4aZbS3xNFJm1NmK3oGFrPrmOtFO7OBvl4kI0Ahl5NFcSabwuLSgt53R1eXbFjzRVrttuDS2CxKBNviSRT0Xqi2jMjWKSgUpXZRf2ODWBE+Wd83arJ+GhoaEpBlbhamDOTa5bW2nAcbynOfDTamfNZEcFUGkdnpWM9o52Jw3FA+GdeTOxSEekc9kZN1FKDstTGvsWyJqzXNUKT48awMfS72vj7nUW3sFknhDBewteX84J/DvMBe22yHjIVvParuodQklrngIhH9LlBPFsksYY1IItWlbCKNyBrOdsvyYH/g2ayusrHXMNWyfW7WGgaqSA0qu3WCXJzVUIljPQbXJj+vqfGsduC1CLWjBvg8S5VnZQBRmIMJtHHgyq6tze9Cfxb+LpB/pSTQa5pS1+6tzTlOfbWzWSceeMlcMxBdP8OJo6p13OGFpKNY3GoEDf491yOoYsLspFl78np8H5W0ruvW2V0on0KmRFNFYVVjAIb43u25DWoJt39yfXNQTTT3KN2zTeu/rX1FU1XhdvQ/CKhw/Ks5C33W+mnrVXz2zz8UV2DEPwUPGW5MfDj1Zw6hvcEJAAX/3ew0zFqkuXm5ksA2edt0xB5xJFuZRg4IBDYAB06B4Sl/RiopGOiTNJkvD6mQl6BwoMAyd3Q4PPDGODDQgpuTye7ZrGyGHZqM0pD5gFgSCAlhSSH0KCgfWIwRgBFbXkN7Y1eY4sDYGgqq8twIA0DsehjTgsoPs88KShIhpu6ZqB/hRQqHwcbSyKiY4j+8vmI2enC3wBi/xiy6BA7J/zGqoY4NH0xmayFDJiO1AGZrfHTwsLEkS4ebuYKo6gpKDQoFY+j5Z5RN19OtpMyWxT6jhceZ969lDlA5wT9T9suiiQNIAybsd8ptqZap4Ed+4o6nARX0djZP7E17gzCIMSYjgQoL0AqNbjgwDZGvKbyPLFI2ijt37hK7l0DF1OQ4jn+XQAV9eg2ooI1CW3snduzarUFRb3+HhhgEKhLJFHJk3xYL8uwkUMGiJQAVJk+0X3VYqFy1woKEB2QU6UxSORUMLDv92HEsTl1ErFJDJtGGCD1sG6aoIFDBZ4mDRtorkdHNgo3/6DmglVPWciLYPPC+MGA2t7ah19bwywdJ/HcCSPFUi0AoFr881M6eO4sTj5wQmMUwbVo/kcnLz8OJC9mHeobFkjTWuliiURtK8XWTBKsIOrEJdl9OhdYp2C4ixYOkp2QxeKYMn6eV5SU8cOx+DI+M4OjRG83DU8n1VoDy2WOTG420YMfOvRgc3M4YNTTo28NKKkKgom4ZGbQ9WF3F6VOPY3xsHDfdcpsCnAlUkB0rrm7MBt5UVASAQgMnBy04sCpXCpifHMW5xx5CrF7UntOSyWBk5y60trbrOWpr68LA0HZEklk8NTGHp54ax1e/8nm84XV34BMf/5jk7vTpjqojtYJRFitiG9salpJbrBEbHvFe2qDP3puef5cD1yMc7JH5FEOsEUUqVkW2pYqjB/dhuL8PKBfR1pYWmDUxM4e5xWXML65jaXkVre0dqEjlS+ZwTQx0JFIo1yy/YTNUVTuf1vrI8Aje90vvw8033qQhFZvtGoeskSomnzqNRx++D2effAKLs2u4eHEMbQyDZuxAJIrHHj+roW9bJiugYtdIH2KRKraNMPcliqnpWSysrGF+cRXpVg4Tkzjx+Ck1N1zrbITDQI2XTwApbeF0TbgmjNXLfYugE6+vCuyoDQS1v1Tr1jDEGJod84B5s3exhod5O8Z2YxMaGDrMWCDQQPCVXv9t2Ta8/wMfwODwMCL0pmXDEI0hWavi/ru/glpuFfPzsxhfXMC3jz2MR06cxE033YjXv/5NOHTkGjx68hTuv/84fvSVr0J7Vy9au7rFgL507gx++0MfFOszWq9qH+IAk+qYjvY0hgZ68AvveSde/ZpXKmOoUkvi4tQaHjl5Fp//9L/h2LfvRbFIhUdDQEUYdPCzh2JYe48z8wSiet4Qh3D6vO5zGlRqm2C+yarBZ4TAshinJeQ3LLuBTK943DJ5+N84MORQRT+fqpR2ejVXte6279yDO+/8Odx624sQi7eg7rYD2pfZNOhstLOZL7m+UVDjf+KR4zhx/EGMXjiHsYvnkM+vS+3AXAqGJJM1zMaYhASueRIKcrk1b/J4TlhdwKDHl//I8/HeD/wSOvt3YGyqgOVVYGJiGmMTl3D4yEHdfxuW02u4KK9tnq8cfjBMm0AFbZiYUcF6ZXFxUa9NRcW5U2fwJ3/0e6iWFwRUhDBVo74+/Veoi4aHt+Hmm2/C0aPXKxdGKstgzZdMaV/mfq4BEj+f7AKiGJ0YQ7atVZZGZltZEHDO9fy5z30W9913n6kqnXUWai9J/x0zYdPIn80DWixN+WXboIZfR3s0KirC/sN7GmT6oU4T8O82UsFfx5SrZqOmesRzFpqqv6ZdkrGXOWzneyUBQesunJXKdLJwz9CEh6uor/FaMzT61ijax0u3ZbF33z7cdstzFKZNIILvi/eR4EhHR7vuJfc7nim0YegfGJRKUVlZlaqGQbQsrLqiolqL4hv33of7H3pQe4gGTf6GuPYl+3fWLZc21Rvk0AgEor+92zuJ/UlLJ+5NzAyhj54GAAStN0Fiq8HsXA3q3kDmsWKCr8lBSA3ra6tYXV4UGG72bilEZJkY/LeNBKT7YrTqpopDaj4NP421qPsYfjkoEuwcIK9xKkJswKS6QpZkA7jm6kPo6uqWNV05nxeAl067wi9OwMLqvmcCFcoeggEVVAPRDoZgANnbllHxdKCC7zPYItL6KZ1OoVapN4GK9rY2rQNazHFwyowf1rnc6wRUtLcCUXrdp7B8ZgoTlydQKtPqkTlpptrluccahvtqX08Pbr31ZiwvrWBkeBhLi/O6Vvx+w4tI0KEqcUN1zfs+9LN6T5/6u8/h4rlRnZm3v/5HceR6U1Q88dhZvOXtr8WBq/bgqfOX8eixUzhwcC+uPnIFxi9P4eN/+Skcue5gE6j46z/7pOpt7s0f9IwK5jdocBWA5GhUWRNveNvtskc5c+o8zj55EYeOXKHXuXRhDB/7809iz94deOOdr5H101/+77+3nLBKGT/64y/Cy3/8RcqpeOC+R7S2n//im7UXfu5fv4LTJ0+jVNzADTdeg594y+2qP7/5lXtw/N5v69zaf+hK/OibXieg4s9/83ew+4oDuP1/vA3d/b148pHHMT05iwOHr8TOfbswdmkCP/fG96FvqA+/98cfwvD2ITzw7eN49OEncNXV+3HbC27C6MUJ/MlH/xof/l+/KuLBP3z8Mzh/9pLWzlt+5g5ce/Qg/u2TX8Ijx07h9te/HM994Y14/MQZnDl1Ed/91jG87k0/hisP7cPXvvR1HP/OMTz2yDG8/MUvxvryMi6ePW/M/5Ysdu7fj2MnHkOG6oASbWRJCDHblYWFBSmvtg1vQ1dHp1tQsle1PtV6LPZG7MVasby0jAcfOmb5M0EdS1tNgZei0WhArIBkWulkaBdmw2LbztwOyvspGyQ3QFURLai4fxJYpsqPRAyztyLbu4Hh4QEcuHKfLE3SKfrm5wXiW1/MZ9D6Te5Prczjqhb1z3B3B8q5ZZGluEepRE1kMTm7iocfu4B0Wy+W1/OW+0aSWyaNldVVnafcM3neUJm/tLiErq4eU4lHY1haWtTfc1+hCnFhaUHgDnvR1dU1tLZlMD8/j+07RtBHxUoIkSVrOWI5YHw9DteDDZN63Kh9bgIg2nuYBaE5wKY1S2BES5HibG/aQ3V3d+ksl61euH++h3GPDkoJ1g7ci7nHPfd5z8WZJ89gcWVZtrXcT/j9CgJO+eCf+R3Fsvqy0EdrCO7Mcb6WnYURqXlVlyno3YOw1YNY2DI3Lg13mX8hf3ojJvL1MnRA8BwqDWfDwFJuFFRnMDeHvSXXMUPk2e+Zio3Kl2w64+qAuLk3kMyomYA5MGhQTKDGZy8ielTyKG+sYnV+CWkC7gSKUgnEkylkOzswPT2Naw4fFGEnnaQlMRWhJDKWkG5rlT3W4sIyZhdWsbRSwOTMssK0Vzc29Ixp2M7zkMHjUtrY/eWMga8l20Xe20RM5LeOzg509/ZoXfMX37cCw52Eas/d5vkVBujsUZkVFAgPqjvCsNp9/23eZIScQDJlbROCimUTJtWKZU0Yec4Y+lJ2eI/GmYOsrP09hbmDuUwwG4Qglc1bLK+T18BeW+Sg5t/ZAJ43RXuOHCbsjFZdH4vr2VBIuM/KCJAGopuyVhyAC2HYAmh8IG+zmU3Sra6HAyeB4CSMItg7EZRxiyJZjrNOdhVLsIYKIEsIpw7kZb7/oGQw4rH90mzPQV/Nchy0C3Ur8YBw/cKeu5V4FYgLUg/5TPDs1/uaP/+Kl8xr9sU1wb4qDPh5TptSxwAXs2C2fklzJNZVvovbPsRsUDqwkKD0/e1cw/cagGzEFN7QoNgyxab186rH3ZopkKHDTFJ1Mu+xqzFCJkWYrYZanr/zuVcN4meIlKOhfnO155ZqbrOsEynF1qDe97OKis2a99k//XBcgSHfDJsNr0vyQ1YAhzdsMOQFR59j3/jJ0Nv6S2wPSTyt2eVmr83f2dc2wDNE2cKizJPO5PH01LegG/rDMvlpfSOnRj5I/3gwaLiu5txtlcJm6AoF25QckFCQZEOFFRt/bmJiNHpoMYsAIuL0ALTBaQiX3lRpCNGmt62z//ieuW/IWop2RWQlVCsqWIzFHrwMTdmwFRHlvwVLDr4vCyS3YCJeK36/bZ48dBtozTJs2SRuAWgJXsd2aLJZtimFvsc3ZQ70LM/CZKDhuot5zppdBVMAdqxBDkOLcNiEIYGh4mYHpQGXTw7itCQgaNCoq2iS7YoKJfM75CZNeTOBCWlXaJ3FoEiGbdafAVSQeelMMA0pwpHijFGzKDE2pBgbfiBaMxBsFGrIZNMCKjgMpe2GZY/UMDk59n2BCobi7tqzV+tikNZPhQK6O7vFVjJFRVEMk3LR2BVseHmf5J3pDNoGMxTETLFDOpGMCaSg/VNueRGPPXw/1pemkKAvebwV1XoEjWgV8UQEqUSLbKf4s6laYOPDwoDF8yb4ZGwgDvFopaMhbLmG2dlZfd1WOyECXgQqWOzzZ7KwPX/uPI4fO47Ojnb09XY5o5ADAw7IaLvkSogGQRazUrOiniqdqH4OrUTKYnWZLDYMcWxQFZFtFwGrMDRj4cXCgUXA2fNnMDE5jhe+8KXo7Or0JstC7jm044AwggR6+oawd++Vsn4iUKF46hhtgeoqajMtSQU8z05NYm5+Abt270Mq1YpSyYCCAFRIsdQw5ZXYMMw8caaRWLSVIlYXp/DkI99FvZTTIJzPw+DwdgwMbFNz0N7ejaGRnahHWwRUjE/O4mtf/g+86AW34Z///u80OG3UadUUgAobslmRaAzkYP0UBkYBqAjFmxU3kF0FgQqxYapxRKtAa4ZD4TXs3zuE7f196M60oCUaQX9fP+bWljAzv4SZhTzOPzWq1y2SiRaJiaXNgQwZThsF2tuUDBhoBr5yeEUVTQuec9PN+K0P/aY8yTcqZO4TQqpi5vJZPPjde3Dh7JMorFVx7sIo4sk4ipUNlGsNjI3PWAg7WfXbBrB7e58Aju6eDnR392N2cRFrG0WcvTiK3EYJpVoNi4tLUoBYlo55mxqgEzPbH/e0Z21G8JpDOa5PPksM1LYiOyFQzYLK7Hv4sVi08lwgSMGvy62uWZGnwZ09O3xG5LdcqcjeLTQgtIL4wC//Cl72ilcg2dqKOO3dCFTUa7j3C/+O6toK1nMrWCtX8NBjp3DP17+BHdu3493veS+uv+Em/PvnvoC//cQ/4LbnvQCvfM0dWkMEI9aW5vGB9/4CCmsrsiyiXUmDUvNYBO2tLUi3xHDNkSvx4d/9Hezfv4fxNThzeQGf/uxd+D//+E9Ym59SeHSxUkfVP0fY60JxG0AK/s61FQbJQWGVYMPvOUpsFgNDSYUs5ygKrvew6wpD2nMCK3S2s6smZOhBcCqMvalhcC2Dr+sRsxo8ePW1eMtb345rr79JA2wOUcSq8l+BEUgwkRZRZBbzLDjx8EM4e/I4jj/4HcxMT8s2gkOM7o5O7TG0hAqybr7eKsFBqfQC+F5Ee1sWIyMdeN+vvB/PffErMTZJoCKCialZjI1dwOFrDgmosGF5DIWNoobnBCs4+CHjmLVBW7ZD2RXc+7hWF5bmFLR+7DsP4m/+6s9Qc0XF/x9QQebp7be/Wgoy3odgi2E1E9V2CV0z2j5xX+DnJZixsLiImfl5dPV0S93I4UuFgx0q4sbG8Ld/+wllZ4Tz3QZldn7LCsCt7qjUkFKOwJ4ChAlg2rBCoaJkbZYNRAjAiuob3x/DGtIz5n7GoX6QHSCHM1zRZKqztmqqVK11EmBLlU7N2J1UIKh5DPx37dPGplTz7YBFaCj5ewA/+OdQx/HcTaYJZu/A85/7PGwfGUGa55fy0IqI0Pax04AKXgveX4LxQ9u2IZK0MO2GrK/MbojWT9wzCuUGvnLX1/D4449JSSGQ29dtOD3BHC8AACAASURBVOPMWotsQOi+EKjgkFwAosCAkEVBsII2fjU0EgZOWK1mli+WV8F7wjDfTSsF3cPQlLpdAZ+ejY015VQQhOHZSlvEOFWwwaY02KiyZlX/7MGQej+8T9YcCwzf8ssaaqudDVQx+y/WwlK08rmXXVlKqtSrrz6Mei2K/FoOy0vzSLWwOa/rnOGP+kGKCr4pKSqWl0zF+QOAigC+hdqX948ZFVzXVFRwgCLwTSBQTaoiqkzYB/BnUkmTzTLM19Sfa+dmpGygFRJZvvVGFCWegRwqSBRGO400nnPLTearzZwCAVkcENNeg2zIlDG9BYgAH/jNdwpk+dTffw6Xzo/pvbzuza8SUEFVw8MPnBS5irkQBBJYs/NnE0z4yue/jpmpeRy9+Qh+/LUvU5g2MyqkPqo3NhUVH/4rG6hUaxpksq6WouJtt2tv4mfr7evSM8+cjC9+5m48deEydu/fgTt/9icxN7uIj9FSyj30udZe+orn47YX3qh9jt/HbKl777oP3/3WQ0i3JNFgOHMqjne87x3o6evBP/7lxzA/Pi2lxfY9O/GKN79eQMVf/NbvoKevD8O79+AFr3kVBka26Ro8dfYi2js7pFR7z52/KhXntUcP441vuwPX33hEvRV7OgI5d3/pW/rsv/3R9+ta0vrpzBMXdC6/6W2349rrD+Izn/oyjt1/Evuv3IWffPOr0D/Yi+nJOXzkQ3+Cd773rTh4eD/u/uLXcfd/fBmr8/O4Yu8urC8tY3F+AVOTsxjasQv1eAKT84uIJlIoMI/H1WQra6vqXcjE3r5zBwYGBozdK0Z/XKA4CRO8TuzB2ls7MD4xgcdOPq7aQ9ZBCQLNGeRy60YAo/ohRmA0bwNOtyKWPS4VbrJUtiBWe+bN+pQ9G89AMW9TKdmcUVFhhBb2wXn09XfjyJFDIgVQpUnwl48yv5/9NM9wKaBiUaQTMdSooqgW0cf6QvmBG1KjytayWMdGOYbjj55BS1uPiC206KX1IXtYArv8ubQCZSA2QeDFhQX09fUjt7YuAhTPRfaYIkNxcFurNsPN9T3ZDObmZjE8sk0gpxjzeqZosWOzgJCrwWtsari8ciPYbxEUUq0m6+WS9dsEAgoMtSZA0tDZLYcF1nzKf+DPtn6Qswr2bxyScr4g8hjnGq76kgokWBg6QY/uAk3feqoSaEXq64FkGO4v/Lnci7gfsp+x/sdVqd6fsnfl68mKKp0W6KL36BbW7OML6xvWY3vPxGdd4EimRecTQS7ZEcpyzuYk/GxGujHQQbbQAr9tQ+d75fnE6yYHCioZNd9gRp39HK5x9s4iTfL9lHLoak2jg9kHa6tYnJ+TTSwVSHxeRDCsRJCIABkdsXWBFZ2dHbjiyn26X7NzSyhXgY0Se/8GcsUy1gvsIbg+aStE3wR3rEhwDygpE26N1rQrlmmi+j0WQVr1ULuUs8H2R9Y4coywuQRJqmYRaMNxG35b+Hiw1wmDdK4zs+ZxGxw/a2W75WecgLKWtIF+Ig9Y7xoC2QVE+eBbahr/cxii871IZSAbKquh5W7qVmNW7xhZlPdFuQZNtQ+vjL13IyW41aRIR0beM4shI9yGmkj2lXIy2bRT530Prh68z5at4c+DK8BIFgrkOFNKmMqf8yoSIII1kd6xgwhhcB4+h9XP1rMb8S6olRoC92RNTfKGP9fBPl6zNWZqeh6aakERgC03MNR6QUHBn7v173VGooEz92wJ034ZrZ+srtE6cSWCSBlui2b3wmozXp+gAtlaW26WREEd/X3IR1sAMn39FkVFsIESKOf7UfiZytAI7iBOIA5fr2vrswLVi1w//ncC5LasISNDm3pGuWjhBZ4BXFju76bTi2y8ngUqnlb3PvsvPwRXYBs3MLcuCs2h7CFCo9O0VzJpnhDhLQE7ypTY4hEXvDl5YPLrOMjmYWCHjTVs3FT5S7JF94e292DDcG5QGjqqKDNwQeg3vdbph++h3eE9hqCgsMlyQ1cwpasraG1hw1m4VNMKPw0LXSlh4AkbMUPxzcrIbrCpIzab5zBw5GfiLx1e8tazBkTNrAeShiZfwx5Z6NgPJTOUBTAHGvwlaanQVytsA1IbNnbtRQriMqmgrpLuk21SLMJteGHIvgLdFNxIyZ8dyLyuJpu0oY++R9Y5pn7j5zB1Bv1542Kd0EopsJLt4ITYJiwcdZiw4VWRRKsnAylkwSNQgkCFqSgEVrBAr1fw8tfS+slenwcdrVqamzuvkYMQ8olmAUdfcfru68Nuyil1HT1Xgx6+ChqrN3Dw4CEV3Y1GxYGK70hRwTDt3r5BXhQxvvnv/HlDw30aYnY5UJHLF3SY076ikK94eBxVAxUVXoG5wItG9ki5bLZHDNGmXDbVEsPK3Cwee/gBhSOzsssmWq1pjvN7IgryZdHPRpyFfoQeqAnzgyV7k7/zM/OasliXuiKdQUdnl9YMG4yFxQV9rZjkHJBzvUc4BGtBf1+fvv/YQw9pVM0QX1ofcIhjAEdMLCquM9k+Jc1eh88MGzK+MAtThrOyIFMYlJ6BusmYnVHJoWiM66RCFgSVTLwnBgrOLkzjidOnsWvnbhy59lo1fQZoWfhYmU0aeL3acdXBIwItIhE+awQqGmgwQDdGGXiLhmC5lRWFpbaksxr6lClB1jvhQuefad9ggI/WjRe5XOss9rgm82vzOHPiQZQ3liSzp3c82bd79h7AxvoGstl2bNuxG/VYGqNT85icXsDX/vM/MNTbjfv+615jdDCjJ8i7fai3ObQSh0nrMCixpM5ykC0MjwQksrHi5+RPq8UQqUaQaSHDZh3dPWn0tbdi71A/OtMt8uNOpTO4eHkMY7NruDQ2qTyI9SKVIvS/TWJgYFAZFfRr1rrIm6WNVVkGAvL+tGdb8dY3vQU/9/PvRJlB43Xaq+Ux+uRJPHbiAV2XbEsHvvnN7+Dy2CUUK3n519JigU01Ex13jQxi364hpBINdHZk0dHRjUojgunZeYxOTuPcU2MoVciytvtgMmxnXNHXnUAx93KBi2S/cphoAYRch3yWCJ4ZGMmv5zozEEjPOaXQVP7pew3MpbxcgW4JD6/dwgbn9TbrNAvH5Pp7yct+BL/xW7+F/uFtiGr/jiGTjOFPf/93ccPVB9HX24uZpSXc9Y178dW77pLP9a/+2m8qfP3MuQv49Kf/HScffRSvvuO1uP21r9PzRe/s3/z1DyInC6FWhUzWBcYTwIsg2qigLRPHz7/rHXjPL7wbjVgLjp+6iP/5B3+C+7/1LUSqFvbcIEvbG9OwZrayb8Qu3BK2yDNBzbBfVwsot4aPDaTYaFI4kInpigyjASmjIre2Iisdrm3t8wR6kmYxYcqLskDd9s5W7RcCG7NtuOrgNfjpt71DoEU60+YqSD5vlvtA0JL++nzWi2yGUcP89CQunz+DE8cfwAPf+Q7m5+b0vHZJ4WA+vXwWuecwhJf7FVmcygxAwywJayXsHG7Hj73mlfiZd/4SltZiWFgEJqbmcPnyORw+ckj7Kq9ZFDaQ4RCblh4cBnHIyf/e0dYtVijX4+LiMuYWZtHd3ol77/4a/uUfP456jVkkrFc4nGfR8L1NDa/V4NAg3v2ed+H666/fZDQSVC+XZTnFfaatnQP1DrGfstk2DSHGxyfEcO3q7tF1Z61CW0U+rXfddRe++MUvNK0ouc8Zw9J8hUWMMPcnWWXI61h2CAZWaEf0obbOdh/WC6ggoUSWkj4I0fc50LpVReEqy6C0bDTYTG/+Cg2gag+FPdrey8wtUx96F+/7pQbissmymkq1DwdCPpgIBItApmDDm2xJCXh40QteiN27d8snmWcQGce0gSEQ39Heob2BViZsAoeGtunsolKKFmd85htONOBwKJ+v4LOf/xLOnD9nQ0vVnd6Putc5v0/PHu0sPSeMZ4hGMSpVzXqCyjExf1lD0YLQwQndGPerFjuXQLYz85oDBAcq5JEtRmwE+fWcFBXMkOG/p5hdkmwxlQx8KBUsGnT+mFWJASI29LThiCv3/DobTmFfq0w3tzHgcNxqAqruWJeYVd0NR4+iv38Y66urUh6kUhwC2SCHjwHBju+1frLzZnp6RooK5mKRRU5ijqyf3G6Ha8POBbNHE0u92hA5ggNkZlTwZ7cpx6Wuc2JpaQnxOK0UYxoecoCWYshrPKmadPbEU2Bw8/LyGqo1WnHxAhDMiQEx3t2awMCbb7rBBn8aGpsVGmtR1s68n2HYzLqV1yIA4mH/lerIBxJWc7ufvBOEQu9g5Cez4COxizV4YNAam9dAF9loOOmKQzA+P7v2bceb3/5azM8u4uN/8SmRZnjeBZuu8MwYA9M+g4FhxggOVir878oDUOAog7U5mKvQQBTZdALJOO1VoliYmUJbNuSXRQRcT01NiiHf2dNtOQqNqIaU9UgSj514QrX07MISCEdOzUxj+/btAp0ZRMyMivVcDgNDQ6CaUZZbHj7Ls4n7iWxdKxWdM/xHTHPPzuLPUMiwBnusL6mqXkc6GcX60jxG+vtQKxaxvLCIqak5XHH4Wpy9NIpcqYokA3xBZncSa+urCvrl8z2/MI9t20dEOBDzlr1dlGdDoWlFx+va3taJS5dG8fjjTxiAoL3KbNVsYEnLxrJUg+YKYOS1QBCzod2W89cZ2lJaxZX0po1GYF+VA0TakNHOh4P6PAaG+nDttVdbmG0sItsrque5vxeKZKXXjfhRLKBa3FCYdiraQGsMyCZoHZjT68iaJZrC7EoJDx1/Ajv2XIXRsUl0dHVibW1FQL2G/MWS+eH7oJcgA4EFqj04SF6YXzBSS34DCSovmF3pWQxktvNZXFxaxODQgLItFGAsxrEx+mU/5JaD/D2dydq5pEBgy0fUQJEAj9QJFR0b/F2KUV/Xof8NrPt8oWB9xJaMJalA3A+eJERepxDWa6G7rp7yYbaGngRVIuzjzMqL+zbXgYGWRq7hG+I+yf6Pr7+xbkRK1lZSC/PraFPmdqZc4yHzQwAwex/ONJRlaTUu3xc/L6+7nccEqmhhahZU6nnVS9meHYBtzSOcgBDO0EAQ4cyED6sG3VybttRkIRZrlJFADS0EgJMJ1Vq8/+nWdkzNzmJpeQkj24aQTSVQyK2p3qdaidctk4miUMxjYXFDfWY9QjJMAiVmiNYbUkjwPmrf4Vmqo4+qjBTyuXXV5lLaMo+TzxvDvLu70Nvfp+eevwiW0aYtZJypBvB5StjPApATCBcBgGoOa/x68lpJ1cIsGZ+ZBCKr8u68jw+ZAzaQh4egGwFSeRb8TCHXiDmMrtJXJliYC6mHts9PgIlAIOsTG+A3+Z1uTWXVk+6Jn8XhHoa5jyZQIYvOiaVUj/L5DzavgbiiXBIfygdCrZQQoUNVLeKkBR/iW2YHnzl3wZB1mVm4i5DiNudhBiV7J+alNK3b3bpOwKv9Pc8g/sxA5AzvJZCqwjkZyEv89zATDOdqqAHDOufPfvIeq4v56+DLLb+OdXMA8sxOzsb4IkX79QrKVREZfU71tMLVb4LC7r/nP2wpcMMfn2H9xG9RPs8WV4twL8JsMdS+ll9qNvZG5LW6o0nK1Xsxqyn+Yo8ji8GoqccNMFU46dPfmM9m7XsNRNJz8SxQ8X1u4LN/9d/6CgyJPeRIrMKS7XHh5mMhmtYYcfNMMtiWAXedHWL5qGmukWVunrOWWWBIMAOpZJvEzdiBjVBc8wkNiLD9XGOLWTBRXewCeZfzMFARYKoGvhfZUnhz0JRleYETiiHze/VAYoUphYG2Md8zGQ467LMGVipBGDawLLCMkWEB1kEZYUFPm5Ybaqgd4RfjwTf3sLnw9QMgEIqMYEXDzZOFeWDT8e95qGqoJJ/czXyN4KHIQojFpAp3HSrWRMtfvmZggn2/XzeFjJtHOT8Xf47kejxoZcFgtlb8UCwGw6FkfuTW4HJdWD6J22vVzXePl1bsaDbEcYZkmWqCvvHy+XWgolqn1QRVIyWBFeZZWsGL7ni1riWLNa4dNtcBHaf/s4FSJk3lPzz8+DnC2mrKMIU020HJJpi1GRuyw4cPmUVPvYrJiQk8zFC8RkQKiq6eXnmqt3f1YNeePfqZA9u6NMjq6+1XscgCvVSqYG11FaVy3TMqEipcdIB4CCml37RGYtPC98Sgv0xLQs3U3OWLOPPYI2qmkhwARONSjhCUUVip/OSTyGSzllPBgb/WUBTFUhlrq2t6fbFjPOSL96m9pwNdXV1iPhFsyJdKkrWTNcb3x+EKn4+WJL3QOzAxPoHlxUVJpTks4OsEpix/ng42DbZsSBUOXv4uywmyX8myTDqgJmaHe6fyM6etodQzoM/pPpPVCtY2VnH6ydMaQNxyy3M0pKPFggoSWiEx1K7McPYUDh66Buk02X8R0AlJZ7evQ0qH+ZnY+JL5xnBpsTxY7Li6iL+z4aLihOvFnjULsVMRw+e5XsHa2gLOnj6B9ZUFxMker0PX6qpDV1r5GI1j94GDQKoVFyfnMDkzj3u+8jmUc2uYnphAQmwYG5yoGNf6cyDAAd5mbcMhO5tyL9D1VQ6Mmn2RXSt+TrFo3GKOYd1k3ndmEuhrS+LqAzuRbUlIWTNPu4Oxacwt5bG0XMLaehUruQ15mHZ0taGny1RBk5OTqChLz+Sjth+apR0HF9wvPvr7v49bbr5FMmqGpY5fvqQim40+95Gv3v1VfPWuL6NM2xiGVIg1zWeyhG1Dvbj64D5UShvo7+lTjgiHGktkOeYKOPb4Wcws5rQeWVwaccSaLm4pWv+09dK6NyA7MLC13ikbF6uVBVjcQ9z4/cbk5TGjZsLBKAM0YlojvCsa4gvwNVk3X48MvXx+CeIcR2IY2b4L73r3L+JVt9+B1o52VMt1efL+3v/8sNbj4YPXYWJ0FJNj53Hft7+BxeUV/MZv/x4N3zA5Pq2Q2T/9X3+IUimHH3/NK/G6178Bp588h49+9A+QX11De4ZDpzIKZbOts+K6jmwmge0j/fibj/81eof24f4HjuGXf/lXpJQy2TuVQnaNDGNSEnETmBYoFnxg3e8/qOL0WWmVlTRLKBtibdpQhCYgNDpq3jwDp5BnwOKagT5szBXmm0RC52sdhZLlMXHoZAPlmEI29+7dh7fc+TbccsutaKV9EVUvBCzZuKVa1NhK4cMzIxrFytISJsfHMTs3i4cfegCnTjyK6anLyGTiiJBpyqFBgXL7uoLcQyA1GdXWhHHQHUF7exwveMnz8J73/jIi0R4sLgMT04u4NPYUrrvucLPh5frJbxS0rxPAK5XzCpHlELy7q09ABZus5eUVKbb6urvw//z5/40Hv303UKcyz4btgVtmBAkyzOzsSyXj2H9gL177Uz+JK664Al2dnW6FZwPuUrGC9WJF14Z2OpT5J1vSatgnJ6fQ0daKgYF+PXME9nhtGez9t5/4Wzz62KPut22bYtjzNNis1Y0xmeT50aJniX/mw6Fhh55/Y5XxHw2HadupHCOzaOA9UY0mCbydp2LZO9BlDnVue6nPnbAm2FkcAQyzIEPLp+LP5OCdIfcGXNs6Nn9yO/vCYCE05IH00Ry4elPG6iOWTGJk+wied+ttyqqgypcqKlmQRmqyfqJfOM9ODne47/d092h4zSGWiDccppSNaED27MpGCf/n05/D6Phls+WQx7U9a1azEAHyPaRMtikHm8wCsTBt2/lp3WCfR+AAG0Xw+1xtqABeG9wLvNCQ0tmJQR3hw1gqBlhDRWmNVMojt7KMEoFDkksSVDWndGbyvvJzVBR0zaGQ2XoGpUYgUfDfNYz31/STqmllo/Y8avkYPBvsHlswuBSzJDsMDgisIAC1tLigYanWRsyGa2ZBQxs586sPVodcC7Mzc1haWkBrR6vZUaZTAuSYS7Q1o0IDQFn9kXDJZ50gVANzMzNa762ZrB4/7ju0vuQwl7UebWsy6ZRYyel0q/aamUfOYz2Xx8zMAmKsVxhCrnqKZy2Hx0Z8uvHodeju7mwy1UMmX7hPdj6xVjYgRXUKB6nOetQ9qNLOL2VKIg8j1d4dLCd4ZWRLYzWIEZhsHw7PjMoNgoXu/c1vpsUPf8auvSN4/Z2vwfzsAmgXFXzwud8YXmqDVLOlcFWTA9eypHEiEut+s9KIoKogU9Y8VQHSna1pneXJeARL83Po6etW/cUajkSfaQEVfVLDGkGAvuUx1KMJnHzklGxUJ2fm0IjHlOnGmnQtt6Yzo6ev1+2AdmhYbEGz5rPPfT3Y6vDamqWoDZz493xtgtFUZfH5oQKENomNagmpeAPLs5MY7OoAn6y1pVWcOXsB+w8dxpNPjSGWZrZRCvlCSQQOPtfcD7meN0oFAcrbtm0z0hcHwQTKkkl9ran9G+ig9d/58zj9xJPKhzE2simNeR9ZZ/IRpwKHwz4Oy8022AOMde/tmQw9n9m8EB6yPZJnqHqgeFI1K/cP9gMrqwsYGuzDtdcdQalSQmdHm8hkhcKGW8wYuGwwaQPJGNRvUFHRS3s11JBbW0ZLJmVWLrEWjM+s4vEnL6G9ewhTs/MCjizzgrZLZfWHzIJRf8LPVygq24O/s5ZkfagcnmgEBe7ttDBKJrC6sqrnkK/F2oV7NDNA5LbgNRytJaWS8rXJM5xqQhuIWq+l68/QczHdSYiw+UAALFjb83oRDFL/66oDvoaRoozNb9u3g3+WiKwelqQHC9tm/c1eh/s9+wTrrXiPMumszmoBKS1pqdpJDhORzn8OFV4EtZiHxD6zs6MTtKHi9eEa01CWeySzwXy/CDa5Ifg6rHv+d85QuP70tR7aHQa5XGd877wHtl6YJWR1l2YuJDlSOeuKSKuJDFTVBXSLPeVRKqujjnqlgHopj3Iuhypts2Rf1kCdoFrSQLeu9jZkkgm0+31VTmGmBd2D/SIkToxPYXWtiLWNChaWN7BOSXA0jnzZrXhqtBKuSXXL/U/20FQXcW3Jgrsuu1kS8whUMFBb900zG+j6BmVwmE8IAHQLpTB3CXVDc0jtNkbh783i28PVfZ4S1qApkswmyGq5aDMonnuR5buQSLeZVRoG7mGNaU1wHfmcyqy7TOVj994+k77Ph+J6T66itOG+q66cxGpErpBpZbOpQAqWgsMJpiHLIgR5h3xXzQ9cRWQ9kJ1NIi155kNQVmh25JkxFiie0POv6+dnFtdUmAkElwLukc33KDs2UwZwHQYLR14b/hNmfGFmEj6PZk1OoGJtH+ZwmkVsmaby9bcCFVe8dN7zbzyjNpB+/VzVOSeg35QuYQ3YvQv27FsQB9eKPGP83wQLnoZf+BeFDE5egwBU2Hxh06YrzKd03jeHAfaH0H+FmaGtDfvh4X0Esne4r9xfNI+R9XnQ/Tq8ojrc1vCzQMWWxfPsH3+4rsCwo7p8cGQR4Wg+LUJ6e3uFGtO7mag3B2UsTOhZubS4KMY1C1k+sGQ7iZHg2RIBxCATljJI/uKGIW99bm5uz8KhikJR3aZFAxR5v1kQDpmCgcVONhQPMiHBvgMIueXXP4PpSGl+kKuFoXxorvkZgszMLHvYANrBYcoKC3sNsjQO5W0YaRuSHYZWvFrjbSBLGJZp8FZhU2x2VpY3EdBS8+zkv/JasBgKnp4stshW4bWTKkShshWTLYpdawHY3AAFLvmBwMJFDEUNTs2XkYWNABf6U3Oji8Qs/ElSRAtc5vCfTDLKU/lnXh82NiwWeXgJiHHJn6kVTDkgWwkPTS5VeS/ss+u+6HtMUUHQwcCJshp8DmD53p7/mh9zcIVMLw6vzEZLzYP8IA2EYWHDwegPAipC08evVQhshHYQBQ0zWNgHoOLRB4+BfOIAVNSZUdHRLaCCa4cZFSxK6MvKe0rQggzg9bV15AtWQAd/xsACkNyWKiHKVrmWa1WkElGkk3GkU1GMnT2FS2eeQKNE9hpDMenvzgLOi2X3k5e9kuwWWuyeSxpp7G8OehisqrUkdk0E7d3t8vYkg51fW6KPvIMMZF0Q2OAzwkEOi1QW6WQsc5jG1+A/YZgRGmYCiWwgQwESFDSmJDIGkiTGbrsVvKYlNZb/qGWSaMilPAFjzTKke3JqEpdHx3Do0NXYuXO3B3kb48Yktpre48CBg7IP4mCBBZOtZGOCUJovoIIhyCwQ0wRQDKzj+uHexM9uGS+0lzG1URgMWCHEMDkOzxZx/uwp5NeWkGRdx+IwEsOO3TvE3qw2ohjetReZ7n5cmJjD5DSBis9ibWFOoaIypmLBHVhDwRv1GYOnZn1C9pSuL0O1nCEoabto6zbk4hDaPWUNrKJCKoaWWA2ZWBXXM69ioAtJggypFjw1PYvp+TWsrlUxt7CBxZU1ec3WIzXZogwODInZuLiy6nYDHLZYmBtfjIM+3uurDx7CRz78u7KVYvApm672zm7kCkUFyX/9G/fgXz/5z1hdXpCKIkq7E9kAFTHY34Ujh69EPr+KgZ5+VIp5DG8bFANrbHoBJ568iKn5FQNgPPhNCKfAXmeVuCKJgBnXF5vDMEDnWhdYoewaY1+bp3FCDC8qFPg9fB7N5s2aWw4RQtHI38WE9sEr9ycCFXUy1hsRJFNpvOCFL8WvfPDXsWPPXrQkMkhmEjh+8hGcvzCG9dUy1hbmcfDAdhTLq1hYXsGPvOoOrLBJm13itA5fv+tL+PSn/h6tbSm87WfejtXcOv75nz6FUiGPNgW/1mQjx/euplG87Soy6Rg++Ou/htf+1Nvxp3/2F/jYxz5mHv9ezNo5GCxcnl5zqCj1QbEGu97cBHk7lSEMlAvPrDVFZgUYyAKh8QqNkO2xBWysrYrVp3Bt2mVwzSljJSabsa0sqMCAInC6e+9+/Mzb34Hrrz+KTFuHho7MThGitKVg5/NDpuPK8rIsjWgvcuHsWXzz3q9iZWkG5XzOzMo4FJNlVE17Bs9J/jvrDNURabLYK7jxOdfjve//VfT07sPcYg1jEwu4PHFZQAXPBK7zRj2qfYFDEYISWy1+fwAAIABJREFU5WoBXd0kW6TR0dYllUUAKuYXltCebcGf/vFHcOrE/QZUiP5mTYfgCgcqgn0I2ee33nYLnvvC5ykUnMobvl8OmIKlRL5MO4kWARVtVFXE41hdy2Fubh6d7W3o6+3R5ysWCXrXcd9938E//P0/SOGhx8bvd/hdTYkDAgKTyGJmsLrXQxoac1YjFrNlNMgCisN9qhlbDLwLrLpgmWDsT2MDG2jAf2y/UMnVoDJg05bA/j6w1mqyfyR4wrqKVg96zghKxzYJMGEdhlXNzyQ1r5Nk7Pp66CT/THu+wUE855ZbcPjqwyKv8BpZnWBAhSy1CIjRyqJSRW9Pn9l3eC3BPZY1DZWTXOsruSI+/Zn/wCUHKrjYeZ4J+JZdpdVJqgWL7oGteBeztVCtpRw0qgx8SM+vbbjExWCMLfZQZtO0FajYek9VGzRqYrpTSbGxuoIiVaE1goM2xDRGpdUHNji3eyJLT7Ed3T4g5GAwy8EBKJ6r5idt1my6lzbL8YwlA295FnLYlmhpkc3bwUOHMDI0qIBvDju4H3DobV7fTgbaAlTYz25gdnYOCwvzyoKxTBkCaRYayrXIXiHU0hpwiPVouUKsa2enprXmSc4JKgKC7wQqCGYQ+GAdL6VGogVR9imPX8Lc3AKWl9bQkm3H8tq6lJeJVFrrL5GIyCLm4JUHsGvndlQrBRsY61AyAjLrPt4jMpz5PeoDfBAS6omQp2dKBVsbGoo6GzVY/ahf4PeH4HiuQVeaaZgjjbNZuHHoyPXGr+c5cNXhA/ipO1+DuZkFfOzP/tmuj2eAhd6J60FqDvdlD8+MBkICrKPaf7je21qNxc4avDWdQrTBPK40GpWC7NOmx0YVrsxajDUd7femJicxONSPjvZORKIkjPH5IFCRxKPHH0P/wDaMT03ykNA9NVZuTX0GWfN89to7OgQOGJPc+5l4Umd408/duaQ6x0VgSoiMw1qI+z0vTK1SQiLaQEu8gXoxh962LGqFPOan5zE6NoVrb7oFpy5cwmqRQGxUgC/Z3LT46ezuxlp+QxamOqt27Va+RMqVnSQ3KFvFWcy00Tx16rSsU6nWYU2j/omqTtoWFYoCefkZpIpPm+f5JhFjU3UXzlkpns35Q5ajYuFXrG8rFanGJoGIWU5rGBkZlPUT96RKqSD7J657sdHzJZGbeHbQiq4lEUWsUUGStR9T83LLqjnaOlrVl5QbcUzMrGB0ahmZtl6s5wt6/x3tWbN/qwG59XWBF6yj2dMzq4BALz9PsOQxMJv7TVTM+3Q2LRXb8sqysmIW5ufR19+LnTt3GHlEyom0+kqew3zuQn/B68Bak709Z42si9hL8XlazdG+s6ZhL79XALTnXHAP1HPjQ3gqIs322NZMGDpz3XGvN7ssghymUuI+IgUJe90oZL2oMGwqKqKWucHzgwNB2l0JYGvUTRVqO63yK7j/iYQJCITRkFq9WEnneui/+XX8eeyp9Uw6cMU9jiSF8P5477mncC0p1Jx1T6WqGkJqYZ9tiBDmYdSs/zItGT0fJItJsexfJwDbAeGUvzaJRDFUMdjTif6ODlSo3F9dVj9VKFdxaWxciplMkjSeBuJijBNAsUHq4FCXFA9ruQKi8TRiySxy+SqK1ToasbgUXwSAFAjO87xR1/rjeUErQp67tODmGlbv3Kihd6BfQEWwGQ9DXJ5j3AvYq4Y9VvkNrOekEjbwN1g+2XDd5izhXGFfHeoKgV8O5PD1uTaoFFLNy6wJ30eD2kOAvKu++AwYGdTmQcZ0t+G85iW+7myvt3pV67AZxGz5BXz+RWZ1UCLsNfZMmO1tqPkNgrQMCdXnrsSR9RND6DWzMuAqWLvq2m0Bykk6EF6lXFQblpktk5FUpbJ2e7CgIJRC0klNmr+x36K1kbuhhLpMcxpeBwKvrpZSZeNKXJ73vF9yFvFQbc4T9We3Kg+ztEA8DrVQmE2E19oaps2MCl7MMJdTSLt/Bv08EbysPg9jf/0cz5Kw6/B0oMLHek9vsLxACu9J/3Hrt/lX6/pxH3fr9VC/hv5TJAQHl7xEMJWrZ4mEeYD9/E24JABQISw+ECWeBm6EGi70BU7+e1ZR8b238tm/+SG4AgQquJGqUfQBtiyZXHoUBuxhYwmbdvB/lnevB09zUxBDXvYzZtEktM9ZxAFpDcWFCgOxnw0c0MBFnn88ADjYs2AiKRm8+AiSO75WyLjg8I2NXkB/9Tra+A1MCMW8HRTGyFV7piGiBYtx41UmhhcD/D2wG8ImHNQOLGT4y9i89PdnfoEdKnxfKtbVnISG2/4usAb1PslmUaaHFV9Cg8m0JJggH2orZrl/yX9QSH3Z/BGDxMsbVGv4ODezw5OfI7BRguWMUF4FdbFosq/jgatQNEehDbzZfK/yxvMwUIEUztZnwRiAomK5aJNH3g/mUuj+GTuQnpdyyubwQooKKmWqeOHtr1KRLums/CHJVjKgokzPfAfMOOjhwP0HARV8P5sKAR5IvFYF7Ny5UwNZspnZbJ04dlws6qcBFZ3d2LV7j8aGXT1WELa1tatxYPFCFcB6zoAKWSB5sPozgQolY6sgZlBaFC3JGJKxOs4/9jCmRi8iQlu0CId9SWOaiM5hYbMskPj+eVhbyCoZsZT68XOU5B3PRpPrhAc/GeHRRATdPd3YNjSiIOjllVU1LXwPLJo729tV4EmNwoyAhUWMXb6s4trsF2z9BDBC64ANNgvKLYqKUHQY08sADhU7WpcuaXXPS1trXpC5B6dC1ytF5NZzuPQU2dJZXH/9DSoQBeSxYJKFhFliDI/sxODAiAdimQQ8ABVhsL66vKKGOZ5JSzLOn83htmyyyiW3hjG2a/AJNbs6AypQK2FtdREXzp1CcX1FRTlVQY1qHX0DvehjDkgsgb7hHWjtHsRTU/OYml3APf/5OcyNXRZo1mAmBAFNByq414XiKlyfrceCFCk+KA97qAXtWbi9GPAspgLw6kNnshRpAxSvbmDfSD8O7t+OVJxWGBlUkimcPncZufUa1tZKUn3Q5YKMXTr3tLfRuzuL+aVledBa8caBmsuAhZFEJWW/4zWvwc+/+936mgrVVdk2LK3lFLJ45syT+Phf/xXOnj6FOPdSUTn5aFXR3dmKQ1ftx+rqAgb6BlArF9HX04l0miHk03j83CjmlnLGLNrC+rBhmSm75GkL814N54mG0wIXbEhqw3drxALzjRJ0MSG5DzFoNZ/XutRwWEW0sdL5Z1mqCPixry0UlxWszIeMlkB9A0N4x8+9E6++4w6kkh3o7u9ENBXF0soGvvyFb+CRB76DPTsGcPToIXTwudt1AMvrHJivIb++gZX5GXzsL/4ITzx2DMPDw4jGE5gYH9eQuiVBYCWmAUm5VLWwbllvlNGSjuHoDUfxux/5Y/zaB38DJ0+e1Hu1zBUbTOv0DKG4vqgCUyucSVaUm3WeNVdsbCzYnXtZOJP0nHvonwAcP+8NCDK2EZvj/PqqGK3lYtFAdp0ZxuhW8+nXM1xf/s5719Pbj337D+DOO/8Hrrn+qBQD/G6qoxpRgkK0aImL5a+BfL6Aufl5rK/mpB771r1349Rjj2B+bsKYf7IEMasLXgjuPxwc8PXlVc89qF7E7gPb8b5f/hUcvPpWLCw1MDaxiEuXL+HoDddqn+L64UflPae/OBUVBCrkb9/aitZsO9ZzG7pWBDHmFxaRjEXxv//wt3Hh/Amg+oOBCj239QaOHr0Ob3jjT2Fg2Ji6vCMc4hDgMfChJG9w7qOdnV2yearU6hrW8J+WeBytHCSSbVgyMOZf/uVfcc/Xvo5KrWSmSSIl2P4baiIOcviXstlMmf2NGlvLV7bhq0vsWSuFM1zqv5SpWDXw9joiNIey//GaLQw/BS7oPXCg50qwp+Ug0KqPg8yKABT+XGXGOOFDlnluH2ADPQvX3vq5gv9waNq0r3JlxuOyFLnpxhtx/bXXad9qXot4owlU8OfyWrNe6uvt06BM65yv5YQHgt20rcwXa/iPL96F0bFRU7PyDHeJvewsaZVBAgAb4LKpFMUKZX0jqZ8hBAJxJOl32x2qLXgDmkBFIADwnLOzSOQPH36HZ51nAVMyWDVWykUU13MCDWsastQFVBBYo3KAFjTa1wSebfoeBwaf3UcHduMe7CkV1tOBCioqfJOx88GVZlK8yHIqhZ7eXhzYt0cgOQc4BLGoJpKy1k5oU4vo+002w2vFZ3t+fhatHqbN2oOKCq6hAFRoiOIDJJGEIsyoyGjtzkxNGSDJ7JWWtK7XxMSEART6x0CKlgyVwyTlJDF/4iImJqb0vDOUgjk/iTSzwWgjQ5YslTgV7Nw5jINXHUCpmLdwbp7FFbOuoAUhWe6cGpM0xM/StD71YM5NFa/ZFXEwb3YOxp7V53KmroVoGkAs+yAPCjXrB9qfMoPACEAceHDAxl8CGWidpnViQziri405Gb4mDOPELncWMc8/np3s4XhdrP+hkIKMVeaNUdEdR7RWRqReQiaVwMLsNLZtG0KZCrFsm6zHpiYnMLRt0Ozq4mS989yIoRZN4MTxxzG0bQSXJyYZeYQCwZC2NtWo9JwnQMF9jDUVz0We0XZNzGs/WOjwcxAY5z0WiOMs5Y11Zh9kfRhJiyaCbg1UC6toFNfR05bVsJVr5eRjZzC8ey8mF9cwv5rDFVcdxPjlcbOnjUaQ7WwXkDWzMI8D+/djYGjQ8gC4dtm3UV3ubgJcn12dPThx4gRGL41JSSJCRIWEr4rep2olDqCcqS3LnqIxysPzbOQ0v+9SknE4aAQu9Z56VDgQ5doh8Gd7JyJV9A/04rprDyujwu4VsxRNUUEbOJ4wulbs1YoFJKI1tMSA3nQStUIO6RZmJuTVb8Ra2rCwWsJDj55BMs2hv50PVE+a/WaLlIS01iMxivU51RG8bwycZ6/B85n7t2yFHKTmoH1gcED2YNybafPW3duN4ZFh7RHKXhT47KxuDXlNScJHITwHHFKrt6W6wcHiVMpskFjbcw8Oocx8hvi8cV/i86J6W4NXs64TiZFDVXeDkLd/va49hf9NQAv38Ahz3My+SgAMral5QOvZpTLe3CLYG4s1TTs12b26XU/E7Or4NQq9TpLcV9H9osKU94Z9q2YB1SoyvGc8hwWebA4kA2OdvTHPhZZMWgoKDd59JiDrF80WbEiua0gQlXMM/3dmh6iWdlsifm/Iw+A5rlck8QQVrC3OoVYoIRtLoL09q/eb7WjH6PiY9tSR4SFoNE5F/OqKaj6S+GjfR8Lj7OwKitwHkEClEUMuX5KC1up45iZY7p/UmswBam8XqbUtndE14T2oNvgslTA4Mqx1trC0aPWG5yTprPU5SrAZ5uwm5D6w1+PX8P3K8cOVMIFMGPpb3pswqFYtIdeOmogyrJW070uJYTkqxsDnPbb5iK2NzZxP/ntzLkSwzHNYpDLYYs1lSmZTaAo04v7tZ0Agflq+hQ2tzRrNaoPgzGE9q6k0DCSx89tyoez7DIwzm3LZEbqKPNhQqn8IlH4tXmsilF3iWSB2dtMmsarZTSCsGPfE6xzvQzRn8pmWwr0bpq4IZ/gmideIJ6qfwufeQqzSfMwdRLQ0vRcJX9+clUWArWHasn7yexAcFczW3FQgskwiaVfWaGYtZX3S5pnpbVTzt1CpPfPvjXyz5W83H9umTXqYkZjC39UyXtMGsEpKY79+qnubtXwAVJ75ykYuCrX4purHVcxNtNu/rwm+2BxChIBnrZ++96I++zf/va/AARaIAgEskDlsPMExLXi8bTZWm08vD3H6HLLQsCwKK8zC8JiHKlnKLKx4aMhDmWGB7j8dgnfEVeBGo03IrC/4iz9Hf6fBv7G7jaFiMsdwSHFHYVGmA1rFItFoQ5I54NAwgIMWL4rEhvDPqsJZQ49N2V1ooFjsWyPvns+OCG8d+hhD3UIc7TBl82/DNgvxMqZbyKcI/nUstsReDBu2Ay92qFlBtXUD5/vga/HgX1lZ8QCvvPuOOyATVCUcaARZo9s0yLMvWFXJC9lAFX5WgiqyPpBHb2DJuYeey8x1wHmgtKxJ+O/O4FPQNv9GhSZLFs8HqHFIygLKMyo8XPv5r/4xP/AJVJC5SxY+2Y/O+AzBUfRjLZfVBHCtBesnvhcDu+z+qkGOWjYIgYodO3aIncTCn9ZPJx46LsseZlJ0dveAxy2Z4zt27ZZ1Qmd3Rr69mSw91k3lwWHARm4dhULVBgRuTxPQcr4HPjcMaqQlA4s4SujZ9KFawOkTD2FxakJWDinKxtkMeY4HB3f06OT6DhYbHLKy8OIzwvfH+03pOwcsLF5LhQLWcqvYKG6I4TMysgPbRjjYj2F+YUH+u/T3bM1k0NPTg442hos2MHrpkgrFDJv6FmOE8b6zIW4OKzks9+CtUGQF0EIFdJqBmAQqtuwPBDvIROGz58W8znYFv7E4q6FQYnMKyYXn5+Zxw403Y9euXWbfJkUBgcK0+be3dVt+iKw0LGyZIIIalUhUzy8bKYIaiCXESKJqgA2vCjQVohq3GqfTCyMBdNpX6NFexOL8NJ449QiKG6uyPuDwuFqqoL2zDf0DA4jGWzAwsgPtfdswOrOAmYVlfPOrX8DEhfOSUzfIxnc/c372wOgIzUUocEOxHYCKcN2bNnF8VnwAwfcQzJmaBTVDUdkcVTbQmmjg2qv2Yqi3HVEyIgcGMLeYw9kLl1FvJLC4ksPc4rIKIoZO8x+uq1Qmi6XlFRXjHBiTPUIAwCxLTB6+bXAQ73rXu/Dil74MNRZ0iZSY8zNzc1hcnMe/fvKfcM/d/4lIuaDClN/DciuTiuPgwX1YXlqQFL5aLmLPzm1q5J8am8Kp85exmucwIIhHLMxbgYAa2HAYWBOzMcimxQz34S6Lbw0LGaYbZ9Ci2X8xY4XPOP97+HqeLRzckfEllVCtrsaRv5RrEGww+JxW1vVcVQsV95FN4NCRI/il938ABw/egHRHVmDFRrGCh757End94QuolVbx4hfehIOHj6B/+x6sFhpYXi2o4alXi/ivr30Rn/y7j2Fpad6KTB9H0vtbzxMVaFUOIMnq4yJlMxxVOOWb3/qz+Md/+qTAtrBWrbjetNcJRWtYUwYs2NdoMXpDxQJd57dC3Q0oD8o8G07bebr1dcLP0c+UWqakpp4ezAQrpNYTKGTWD9qj2Yh7cxGalDaybiMxXH/0BrzxzT+NG2++RXsjrwafSLFs02kN9rkv8b6s5XKYnZ5DMV/G2OWL+O6378WZ0yexvDAlSzEyLk2MaQ2RvMxTKT33BgzH0NIexRve/Ea84pVvQLHSirHxBTw1Ovo0oIK2ZcVCWcxRZpiUq7S2aNVgjbYxBCq4llZW1pRTkUxE8Ycf+RBGL50CqrSx2FRUBPWgniXu4wB+4idux0/f+dPKnOEQlucVG29mCrEe4HlSrkOAdzbbqv2UOTIcpHHAkCFA7Tk2HJSeOnUKf/2xv8Ho6GUwXCnsKbwSttcZU433gfdNYF4qKTBOxAdvSqmACt8T7hl/52BQKlIpPzlQsWsc9h4Ok7Tv+lkRgFid8nXPQgjhpIEdpvBDkhOMXMDX2WAeSNHCUZVxpAfDhpVb1w/3IzER3dYyrG++K635REJgxHXXXicrIg5+zCqSTFYyY9uRbW3TZ2DzTsYww2AJVFg9VkFFGSUbKBdLOjuK5QY+/6W7cGn0kuc72Xtj3SSbSuUyxbVeOWDiQEwKFQ7eIm4T5UCFAqz5uVhfSR7ng3sO7z0rzVKvnVLtTW94njXEEomhKqCCBIvyxjryBNW015EMExMxQWQaDrY1nLGBRVC7yIrM1a02EPa8EoEpJFRQiWWMVoFODNx1e0VlKVDdzIwLWUjQkpEEiozyrnaMDCNNVQdrQOWQsC5mc25rx4COzW5+dm5OQAVDe/nMyrKpJal6Qc9DUFSwDPC1xBUgUAIRARX8jFQIBgCaiopslgAFFXhk7dPKMqH8jlQqjdlHz2F8bAKRaBK59TzSbZ0oljhUi1pUhUkXMTjQi2uuuRrVCofLBrZwUCqrsDKHqRZQu7X+Dj2B7pVsPo3hzmGqLDSpfPGaOtQeYZ1zwCQvex9kq19xm4ugxjZbF7NxCmpuMpx5pvFeSb2lXshsZnWvXTkRzjg/FDSs0FnguVCByGTBzLQHLWNgsBfFVaoLS4ihhunJMdVmHMa3tLVjZWkRM1OTGmDTso4KPdqhVkksiaVw4vhjGN6+U0xsdgrFSsmHkks61xi0TRtIghRtHW3NIZqyQPhMycLPAlrDHsW9K4SksjZQz5My1QqBlXp5Q4qKJCqIVkpoYXh4voSHjp3EoeuO4uzlCawWyqrxCxsF5UPRmpXnb2tHB2bn53DlVVehf6BfPzPBnDOy4Dngkd2hZThRWf3oI49ifHxSKhCzzeQwzO1cuPeyrnTGfsgZCTlctp1u7r0aaBEw1/CSpDwPjpUFHi1YtPu6cq6CbDaFF77oeeqpSWrgWcI9wayRGMLdYsx/gpC1MpLxhkK0OxIRlNaocGjF+voasm1t2Cg3cHlqCRfH5tDa2Y/l1ZwPRysaUlN9RrvDXTt3YWVl1XMjGZzdoX6it68XY2PjsjnS/RJQWkcuZ/+NvSh7iZWVZYzsGBawEXJ4ZFMSgeqtjs5O/Z5tzUqVEPY+foHZdNq6F1OdllY+K1CfJcDNQH8+O3wGCCJQ+W69tYGJ3JNow8Xv5/O8ZTtqzhNk2yW+je19PEv5dyRFBJcADtFFNORgketCfbMBmcFKVmvWg25le8csEYInPpuQzaXnz2gOQMLJluGz5hhR2tIVpchRdpjb+3AvkPWc9oiQl2mKlgBU8plnXyRmu2eRUfnOs91qOVN58ev43Ee5h6CCFC2gShUUVldRLuZRIjmGn4Ugf7mK1kwLMgnWLlZLpDMpWWUPb9+m/XFmdh65jTJyG1Ws5StYWl1HkfeN4LXAHruf7InDPZYqkepPJzDwevK86x8aQltne1MBHcBL1SrVWhMg3tpzq6bnYN7PveC2YXMru1ZGrohJZS+CjWf46Fr58FzAQFDuu8pD60qAkAWQs69QHUQlGPf3kNFAhZeTKZtD8i0qfq1RD3DXPMtDpM0W26wORe7zWiiQfrR/yJrbgGq1yK7iUNi3B2IH0DrUhXwvnAkIJHIySJg3BdVJEzT1n81rIpursuXA0L5atpYenh16DqnZFExvIIksJX1tUgUiZ44yCbSmOpI6w2dFJBcbcWozrzH0H3y+FHjv+RYhuzUAN9pCo1E8cbdZg/EXFRWhrglAJe9Jsy6OMUOJoeJGSuPrm+XTpiK5+cP8D1trlmf+t+8LVDiww8fLMkysxvMXaa55kXDc6rA5MXXyWXidLdiHfXt4TyJOGMjC9RhmsM2e0JXH4XsMQLV+8FlFxffcxWf/4ofhCtw8OOhhLZbBwMKDNZYYHmqGbPM2ZiKHzuYjF9gGZCVwMEoWBhsYbi5k/VsYFBFts+vgYSqGEItaFgZi5ZuHOw8bbjiheeYGI0/Kag3ZDP1NOVwJQT/czOk9WtOQkRsCCwsNbeT1bl8ndoFnP5jfZVUByXzf5hvJ0GDLqmDTwQEDgyyN5WI+qgEwkf+l5wQYUmx2VRr0M7jaNxV+rwpfR+ipjlDgo/PreJCyeeYGxuG3hYmbT6autXuPau7umR1izpB9z2BTHxwE1rGaqTrDrow5YjkHDOQq+T2y4s5AHfdr52dlkJQzsMQY8SEQN0QyoniQio1INmiphHYWvIUCmBWgALQa70tW946yacm4dY0IYHD4WNJhz/fNoaIpKywcmSwEAhX8xaGjgCBYHoJZfdhgkcVvgYGcHNLL33zTFoWfJwRwKXxRDDYDWXj9DxzYj0qlJBYd2c20fkrG4tjjQAW9+zu6ejGyc4eG4j19bXoNSoE5CCDoREUFWV35AgEiAyps/dvhGhpW+XDSE5dhVwyzSydRzq/hiUcfxOrCDBKIooUgGwtRVR4RsTfJOGExznvP+6ZQbQ4ieI19cEMlBe8Br4MsbghWbKzqfbW3d8q6qr9/UGw2AhUz09PKo+C9HRkeUTNDoIbNXms23VRT8P3ztQyEiyCVbjFromAD588Q7xELnkym1YaMLu0MTA9Tf1hDaR/NwrT583X9a2YHsDC/iPPnL2DPnn244YYbLDDTLSuSiYya42Qqi57eAbEO6Qusolw+28biZCHEQS8nU2Re8nkWs0YCFfORNisFG7zZ0MYYMLx2XD+F3CpGL53Ho8fvR6W0jr6uDmN/8fVbEhgaGkKiJYuewWF0DW7H6Mwi5pfX8K2vfQljF84aSOFNh6XpGCsisG7CYCIUnrx+sh3aoijTPsX9gMMgvmdXNomV44WrijUO9fnfqyVEKgXsHu7Dof270KgWkchmkEhnceHSOJaW1tGIJTG/5MoaekzHGDbaglSm1QanpbKaOQ4RVcj6UJJrsiWZxKFDh/DuX/xF7Nl3hWTc/GeO4NfcLL517z347L9/GivzU5Jw05KHRFxalOzbtxP5fE4FVqWUxzUHr0BPVxfOXbqMR584h2LVh+ieHyGbP7GW3EuVe6f7m4bhOZ8FA7ojKJZo81cxINPtxwjC8Jxh8DOve5Bwy1ogbvZmpooyaxH9XC8YtYYiFXlT53MbChdW4ZtM4qU/8nK8/32/ge6BHnRSVRFrweLcGr5z73/h/OmHsa2vFUPbhnDri1+BUiSNfKkhKyEOuxZmxvE3f/Wn+O5931S4rwKpZfFmgZIMn07EkqiUqKojK5aKwYjA9+Ht+zAxMWlKhXD/A1PdPVilbHMpuUAmgh/O0hKD2Zte7lFmP2I5FUHRF5SL4Xzg+gz/hCF0UPaw2Sdoy4Bt7jMM8tTzrimzNULh2gaFBn/PpFt13Qn2XnnoMN729nfg6sNHUCFCxnMrHrU9TkxEFvG0OKlonS0tregMfer8GXzr61/FmdMnkFtbUPgX9ztAAAAgAElEQVQx7Q1Yl4RhBj+fzoaCgVPRVAVHrj+Mt9z58xgavhqXxxdxaXQcR2+4xq3DjCXN4QgVFRwsVmpFZFszGqhlWjjUsTOPzFICFcwZ+oOPfAgXL56UqmkrUGFaLwP9+Lmv2LdXQMXzX/B8xKVkrArg4XmSTppaToPQekMMYa1NMjH5XHKYEU+gtYWWZQUBJ3wvX/rSl/CZf/uswLa6zsOtAd5mi9n063Z7NALfPE+4/gNQYXoA+2XqTwMQeA2CvYFUqSHPwK0ELOPCQoDD0EnDD4FnbFTNVkbXwRmHUqVyCCrCQ01rhEAFwTytLdVLYX5ntYj2wS0DPV5oPqP8mWpiA1gXZ/h4FlddeRVuPHoDujq7mgq/OBUVnR1SExJC5Tpa38ijp6fXrA5TDC2tNYPEpRrK57GyXsJnPvsFXBodDUhqc2DOusHY6HHUqc7y5ltz7iZQYXCkXbugqODBYwJTEi/MRsGeXf2Zvt0epm3guQHsuj8E0pm/pAa7gmqxgMJ6ThZy9HnnGiS5hZY6pjAmA9sYj6ZEtpUZ1kq4L7TIY71qYIr7l2uYVNMzaR/eVBE8GcyLPopo0ggN3DPaW7PYtXMHBvv6BF5QPWdDC/PotkHuFqZ/JAoCFXNzBCqyqj8IUtBKiiuZa4P/BMaj6lrZt1KJndZnmZuaskF1SxqtWdoI1ZRRwXBus8uMoYVB2hyqZdpUg22cZYYFh6Y5tLV34eKlCcwsLHpmD1nIVVx/w3UolTawbXjQ1NCeOcVrKYWnZ60IOGA95EMIAyJMSWqEqGD/YddcrHB+rhLVciQvGdnIbGCMoMU/K1fCnw8TwxijVvWL/+zQC4Vnx+xoYwZmeXhveG4MmLYzwKxajMUtJjZ7plhCuVMEfGoNDrWjqFWKGOjtRjG/hmJuVXalVFQwDLlaj0gNR9s21pP9/b3o7O1HOV80G6RaBNVGBCcfO43evgHMLy5jo1TSe+N9IjhBljTPCQKCtFoa3DbUZFPzszB4N9g+sVekLR/7A75/go4EynkxZJnlSt3O9ixyy7Noa4mimFtCK/PgEkkF/p45exGDI7vw1MQMUtlWxFMZLK2sWe3a2iq7I14jDoW3b9+BHbt2mtVOIa99hY+AMriYtFWvo79vAF/96tewsLCktcN1yPtm/WVDlmDcuwk4U3XDNWI9iTG9DUiyQbP2PuUQsNbgmWHnt/pTOchRje/OAxoUlpHJJnDrrTcjFmcmQl7KPAsV5rkPtGSyUj1GG3Wk4nVTVESBDO2fYg0x7dVTx1JIZTtx4fIMnrw4hr6hHcjxbCpTdVbAwYOHMDM7q+tOy1beBz5vfM62DY+IUU+QamZmWrbPskFSz1wV2ZCqmcUls0hiNgnzKZhtwTqcvTwVf+xzeF24Xmn/wh5b2Xck5glMiIrMyOtDIhJVjlQm8GLzuvF7+WeC/EZitPOM109nLK3iqKot8r3bzw9Wctx39DN8PsDXZE/EwSl7WgEL7rBgfbZdZ/aRIa9SaiQSFvlM8ec5CcB6VQMSVK+jIRIC+0+dbXxeSfJwR4dSoWj9eTSuGQvfN19TzH727OWi9kkNe11Zy/dKMIlDe9bwQdnFZ57PCM8n3TvPGGUvy9eXUwL7C/ZxbjdUphq/VkRfZzt6OtqkkOa64uvTrnRyekYKmp07RrQ/zFLRBqo+izoLu7tbtYcT7iiU6ihVoyjVjNhUIimUIdIFKtDMvk5B7dWa2RQRZKrUNCuQNSX79EoZfYODSFNJ6sREns283nLBCCx1nReWcxIA3PWNdQuTd7JiUAXz2SURJfS2wZaJf69hvsAsc2EgedXUJry3zC0NYfKmVBDIJNUnFcWWO8FfIcQ5MPhVFTspNLxOcB/g+payvwmOGOnEailXTfv3itDhRCNdQ58zaNYg9YaBcPzFdW8B5xkrTY2zb/WU13t21pjylOue9aLZ79mcLFhtW//p5AUBLFZrNoEKH4Irt0uzJLNJF7E17NFueyXLIp7jdJGgYrdhajkqhbgWDGgxhU8ToHaXDg3hXSEloN9zH8/c09usYfe/eMZqGFllmWLD6p6nq9DDLIzribaZQX0rNYZnSqk/E7Nxk9RoIIiRLwLho/ni/gcDVGhL7Gqrpu12sTlfCfuTwEgBLkbKbAINTqiWVZwrDO2MSVpelROk9aw4YMPrxXVq729TYR0EWqam8TXwrKLimbft2X//734F9kn6bEWVGC3ezLLRYmEh6bCrGsTgCWiqbEviOhhCEa8QIjYazjTRgdXaqkHn9PSMNlaxY9xbXAV/3DztZVmgcB4bcorxQnZ7yT3GYyavJPNbrEb6KHpOA983N3TaO3Bj5IbAAaQdIIbMCmEOFgd8+BuW08DijEU1X58HjPndG5LOYjqg6xbozaLTmjdrPEw5IWCArG8yI5zBzd0ueEyymeMhY6xGGxKFwRyLHx7Ckik6Y1KHoq4NWY/GmGOhooBHbfJW7PJ1s202ROa1NCDIimkV0Mra8O9xtYs1MOajaNd8k63F/8b3SSaPWXrRb7Nqg+W65SZkqS5gBgFBJh9m0IvYivGigrOTHNaXimaTIIaf/iRWUKVawm2v+lG9TwIVyv+gNRIbKTZwFSv2ee1K+aK8LTlk5mcLtih8LX52fh2HO1b0kwHJtVPG4cNXK6OCP2t8fByPPPAgktGnAxVdPX0YGhkRC5UZFRwU9fT06ZrbAJKF1To28ibHt+Jpk8UaBg08hdgkEwSLResacq2vzOP0ow8pByEVjSNNay02kTw0xV7ZBCrsOiT1nEhVQel/3MLcVbgx6HZ9w4PemMlQxOISM2PKagj37jugAoeNAiXaczPTGB0dxbbBIR16K8srCsqjosKyI+ww5loPDBNeg1jChi3hnnNNWSHIAYmxGM1aZlPqyX8vabBpBT8Lv2DXxPfpRDQsLS4LqGCje9ttt8lvnEoWPo9UVNAGJZVqxfYdu7UmOLDQ0NYBPgIWGjrTniGVRJTsbmcTuXeFDxjINtwcfnHtamC2saEieW6aeRkXcPb0SfNr7e1WA1+hvUy0IX/5THsnuvoG0b1tJybmVzC3tCqgYvzCObMLcqYS37+FaXtA7BZmRxgC8zNwrW61UQkDBv0Yz3rR80z1yBYbKQEXVHrx66oVtKVi2LtjCH1dbQpZbPDZrgPTs4uo1GKoNKJYXVtX881njwU1m3YOtsgk57CWmx73rxBSTqCXzQzX3kte9lK89W0/g46uHplDcJA6PjGGYw98B1/+wudx4ewp8y+n9QubZoZxdrRyBo0Nhi5GG9i7cxj79+5RwOaxE6eQKxqoHYZ5xjg1L3QV4LqGVhwHQIn32fZiG0Lx7wsFAp8mF+YgKqkGzYp1AhV8FsnW07PE/TRjftzy+vWwQZ0JiThqZBHX6iiub6BEyygHodkQvulNb8M73/1OIBVFZ/cgUI1jeXYWTzx6P4rLkwLeb33Jj6FjcBdypTry3J+KBY798J9f+gL+4RP/L3Ir8/KVZ5NXl389h5vczwlEsXlnM0Z2ljXELemO5pmgwZgXtGoUAlDhwMVWpq7GKq5+E3PNGWayeuJQMmoDknDGBvZ9aKJsz3Qlkq6NeTwHb34qkHhNtf9WygIvyEYOQEX4Xv587l9UvVBVYe8riRtveQ7e9Oa3ym6vruRzOzc728h8J1ORzLGGvI3pZ1/kPc4XcOrkCVmzXR49h4vnnmw+b1LeOTue+3FbK8M+yyg3VtHV3443vPln8fwX3Y6x8WU8dWkc1x89okbN7ACoSittASo4AMg0FRUb6xxuJDVk43CqNduCP/ro/4Vzp48jUndmpgKSm0RZ9VGdnR14z8+/C9ccOSJ2Ke1RWGfwWgs4cyWI7BZJjKDCQl7WFf1DS0z+HYOTOZDiHksW78c//gmcO3d+k025JUDPmk5TtLAWaoJTibjID2KiuvWTFFDNxtWsOGQpyJBaB1oEVDjYEEIXOUjQOeHZFAJjQ7C7558EkCrsZ9Ky1S2Xio0qf26e5yfVsz6IlgJFG7S11BqqS4AQBnWmMG1aHDSZ/5ZdsHP7Ttx00w0YGtiGtmyrGrpkKoaOdipj6BVuORQkGnBoRAINa0TWD3xP/EWwn4DV0uoGPv2ZL2Ccqkc+c7wgJHNIcWSggcg19BKXk49nJnGgHAuNsSvTeE2kQoiaSuH7ABX8vNwTAlDB96JGNth8eK5XTKqmCiK1ijIqivkNy4xpmLqM9UEibrUSVZ/B+ql5o31mYfc0qCp4tpvKykATG6LxzDejMhuSy8rKw8GlsBTIEUNLMoHBgX7s3bNbg2RmaHDflB2fPLC1y9tww60hqPKcnZ1266egqGD4dH3T+mmL5QP3L85rqZbh+5GiolLRv/N84vM/PT2FNq93uRw52EulCYBkxKJcPHkB62sbsi+s12O4PD6FRiSu4TuVKSRr7Ng5jAbtdfp70dbRLm9w9hk8jKUeYz8UhQZpVBiHM1zAsPdJtk+adZmsgFjPOwM4EI/kJV5lMK8FuttA0wErH8zxfhRpQ+gkKMuyYM5aWed3c1jiQK1zsZp9AoeMfC9kvvPPAjicea59Qr785o8v3/5qEZkW5iTV0NfXjVJuRfZimWQMy/NzGBjoR7UelQqBhJe52VkM9A8o40FkrAgH7ARdI3j81JOy+5ucnUXerWlVD5bLGlIyW4DKt/5+KpssqFiKPhmc2XBXmRS0CVaWDM9DW4sa4LqSQgxRrotkHI3qBlKRMtIxJvaWNZAnwHD6yUvYvf9KPP7kOdlXsoZbK5Rke0nbKgLQPb19mJ2bxdWHD2tfoJWNrgtV3q6AMuCA5IdO3H33PbICNKKdDYwCQYefgWHdWijew7KP4dnJQb/OS1o/+towwMICnLnnmQiS/8f1QAWoV7oRvh8OIJO49babBCawbudrMC8vk20VeY+ALBVKJIdkUky2zyOTjCATbaBeWFfvK1JJNKksgafGZ3F+dAqtPX1YWluVukGKbQ+KZn01MrJde9PS4pJqLG3MrAvEfK6qHqMCkLkQvEokCvC8YaA29wqqI7cNDaKrt3tTNcI9qnlNjMzU7E/d9ljWV7TEqpodIZ8bqmwJLre3m40SX491lpjofC6DgtRnBnx/1p9zf6NyMS1wgh+BdSKfDT4Xa6urpjCNsv+xYXVQZxAQsXPHLJ9NjVQT2Ka1SNvlZFJrmraOGvj6muCzwX6bvTPPG80bIq7qoBVzIml2sZ4no9pe56m9Hgk5UkDTXqlo11X3fD2v/859jqWgWP5uYWVKElqcEtAL6gUnAAhgZb1p2VFSWBEkrxSRX1tGbnkF2VQU5UJJijeuq42CzW52jGxDR3tG6UfKbKIVViqObHur7L3m55eQL9WxtJLHWr6KWjSOslQn3GcNSFJN7caAfO8EZzhT4Jqh0oLXlfXPwNAA2jo7perQvMWH1uwTQnZWM9/DM7JY8xIQMaDCAQUHfgOZUAq3UC961iafR/69ATy0/LJBe6inwn7Dc1NDdT6nwZ7Rh9p6DpxQyc+oOZByNc1qVhbKbi8lmzG5hLh9k4bWVvNY5oMHbfschmsozHSCBVUYSnMexHqGYAZfh8+ggeB07dhKYtmcRgZQImSr2vUgUcxfN1gIOjjOn0fVSFBMNEl3IXND1pamhpUimrZ0JlM0O6Yt+ShBjShApvnfqAhxtUWwxOMM7v9j782DJc+v6s6b+TLz7Wu9pV7t1dVdvahX9aaWGi0GLYxgGGEwBiyBCduAsfCEsT0z9mAjazDW2OGJIRwBMWYGJINBRh4wCCS0otbaLbW6W71vVV171du3zJfry4nPuffmy5ZxhOdPK/oRorqqXuXL/P2+v+/33nPOPSesj5UNxv0YUApc7M179sJn53sf6uZ3rvbGDkQshpUb3yAyKOw35bKA60dMoKQTR9YmLgrwKQ8J9zQ96RP+vkF5EbVvw7V/XVN0ktif7xVOhma/lftT1tWeqejW9tozeD6iZ3NygUlg8E5s3lgHMQUSmVVexyG+ZmK5z8KXmjbEP45D+CTVa9ZP+/frtf/6DrkCx/HAHERl7yA30wU8pvK3lmrIH2jZxigQNvyNCyaSAgUFGzsFuhcVCR2ailZNV5QqKhJQMNaq7lWqFkuqMA9fU9ghDVo8cGw2BHxtbe2okaDgloJSG7wD02qOeXjD369fuUxjyucA7JPCOV63SYMVzLOre93LVwBNbBpscgo+DaA/m3K+l+Yjx7H4vAke8bPZNbgO+vvw8qdA1USG2HgfSWOj1Dhh+FjyewoQNq9eZkXYTGm6JUAl7kn+XvkaFcKV/JBMZR7fm16NCtSLEfZkytNqStck5Ck6XOPA8zF1JzcSvJIahhFqiioOeoKrdT56lgiHP2olhUEOePOM7Q9/x/fUdrG44Fq5vcGD3/+9ev1XERXkKgCkkDXQ9iAxbBpQP3OdUedk8ZHe2nxW1Dj8qpBgrDcadbvrzjsM1QXECfkMj34bUYEibGZu3hYOHdLamjkwqvs2OzffIyoARmkOqoTXjYz66HaQeHkgabqmRMhlRT+Pc4JwOxTWLz3zmO01d32iouzB5TrAaTM4VPGvV1i1X2c+r8iKsTErQtrEaDxKHP6nMU0VdCZS4tq1Zd17pkRownh2OOxqOzv28MMP29jIaPhYm64R47/yCUcNEEHeOVINYMZzRbGcRBZFGPeVtc+oOUQSTUt/cK8ItGwcAqBgDYv9bzWsxIhJoaCJCvylr1xZsrvvvttuv+MOAWrKaCgNKfByoDRk11132sbGJwQ4uVrVCyPtDajEdhs2UBmwwTH3rGbNadxY9mRuaUPxzoFO47G1talGanVlWZkL6yvLtrWxaktXLyhH5MjBBZshRBDAuVGzhYUFBQFPzy3a3NHr7MpG1a4urdpDn/kTu/jyi05UKAga5Qh95n7oq1umBYARSpwsRnJf0l4TiggVZgr5kjGFA44KZQ3wC1C4VBGYKRV9t2OjlaItzs9IAQmRMD45ZdeW12yzim/vhILVt3c2ZXEByAwBNDM7p2u1jTWdCs1931Ku6zAB1I2G/IZ/5Ed/1N7+zu+1UmVITfjy8pJ99StftC98/jP2ta9+Uc2vdRxkxq+d1Tw6MqigSt7T3NS43XHb62yrumvfeOIp+dcCBCU5RtPvZHSEiytXI0iLPksiFeDKMAHIhfhmcmsnnnOadJofgiXdGoO1KjunUL1R1GehnUSFg/kFK6AUxiOZ7JdaVTkTajoLZtNTc/Y3f/pv2o/95I9ZpTJuw4MTNrDXscvnXrBXnvq67TJhUBy2t7zrB6xpZTVoAMzYMaytrNiv/usP2Te//hWFjSuoEnC7hF0CpGPHSoVBn1QUcOXnzeDQuE+79eZ+nYgWTdfn69ojuMKjtEe6h8ctNzZBa66X26e5pQX3PYlVKZYDaPO/3w8FTJJE0DH3QyP4rur3qaR6TEQ6UCkAOkiOwQp2LKgDvXFlDb35LW+zn/iJn7T5I4CDPuE0XHELuoKuj/tyL6+t2dbalnXqHYX21rY37eKFl+xLX/y8Pf3E43ofmi5K72LO1iIey1PWHahat9S2d37ve+wHf/hv2NJy3c6dv2K33/k6ERUCNyAq6hAVZNpUrb0HUTH6KqKCsxWiYnl51SbGhu1f/+8fsGe/9TWzrtdFAnNDvyXQutC1W265xT7wT37RZmdnJVLAq1nXOeyxqEGk5CtXrAyJQJaEVHNY37llBWHaly+ctwMHZnT2fOELD9mHP/yRGKFHHf3qiQp+doKhCAZSrYftFI0OZwnNo4Cq3sy51xD9xG2GLP9FRAUEbJ792QBqIkL1EI2ST8hqbw6gXXVJWDv2ExU8t16buPq/936D2HUVuROVeRbmRGyes3sQEpVBgab33nOPXXfipOzmOM+GR1gH47L+STssiU8KRTvI+Q7QRl0a5wPZKBA1y+s79tHf/wO7eu2qTxDEiL3WPfWPtgSmKiF1YnKC+08jjfWT0EYHnvczKpx85zO5qAWwIpR7McXgG7ATH0lU5Hkir2kBS00rYouHYASyoo5QoaX7ioqbHCCBe4heekRPXzMdZ4hblro/vuxJwsYGgEFWFhUHYDNTo8uNpz6gHuDvNPTnZPv46Khdd/KEnTh2VHWc3mvRQ81d0BhERayJlZVVu3rtsqyjIEfJlUCRy7nHmstw9wTpBe4pi8YnKq5e8ikz7N/GxxywvHL1ihFcr6mhLsDTkI1NjAl4orbefeWK7Wzu2Mz0rCa5NreqNjI2pelE9l1lQIwyFYB6tSirIxcqIdjh/SuAyW1MvVDv2erl+gQ00vWJqWm3XfH6Xrl4MWWZwJfXuT7F3LvnAYIweEdugfzNY3dxgCv7FZ+4lgVt09XXbqcT4ErU8N5LeG+kni1DVdUXeFiriDeEEZ2WpipmD85bY2PValsbNlQu2ebaShAVZpWRUVvF+nFlxRbm530SjIlAADxDnLJnTz/zgs0cmLPLS0sSTSiHJ8RuPL/UUleuXtU11oQBgo2YdAeuSstT5RP2rETCLz7OFq45zy+fr17dtkqxZUOljk0MFawQ96G2U7eHH3nc7rznfnv40cdt4fARK1QG7cKVJT2jrHV6tonJKbtw8YLdduttdvDwwSCPvBfza48oi97Je83PfvZzEkhAKABAp3rb+0/AZQhsJyhld6I9kykqF7DlWSWipQBJPaS+SpYvqYAWwYfwLnIEKK/26trT3vSm+x342mvrGkCwMsnGc4IQQeug0/JpijLhxy2bGR20+ua697ciJiu2vLpjL527ZFfXdmz20GEp3wk7htxaWV0VUc77xvLMRWneT3E/pZwOkos9C9CZnk7TBiUXMLKX0n9gBXXyupO2sDivfAz3yffaj3N4a2tbf6bzSfuMizJEKmtKzPMTsTsrVXza3MOOvf8ilwpRStZzyqqIaTnuhyaVhAv489RvE6xaUPfBLbjIKcoJ8cy0SMsbAaCA6azLEtaIhGa7lY/yZABpIbIhn0Khz/meOIS+B9A38ueUUUNP3XRsBJU9zxOgs7I3ZDHE3oA9pk/vpOqbfT7XHfcBeyrvC53rh/jSvqv+3UWZvhdDktQlRmDtygJnr23dRtUOzk5bmUyZrS31PfybWr1uS0sbqkeGB8F4CBTHqtMxn4nJUZtdnBPJuba6aY12wWr1PVvfblqrW1CgdhO8peAEL9eOPU/T9QLiIVjqIoboZySeLJisi0fGx0Qo6jgVce8Eu6ywlD/igH/mWXHNWXNpL94vROKcY72kWp8+N89YrmMSGAnyS4gRWE2KOhML4R5IyCmMaT8XQrgJ11qCUPYnD612qyW34ObnQjxkhoU/x57Fp/otsi2EW8SX1+n7NkWy5Iw9k2/JczZxpbQD9Lv97V9uPynxJpMhgR8xje71Dc+Jfz5NjUQ+qr/W/qvldec65bnmn9+tv+VaEBZqqonj/asaCNzJBb/6rqiHnEDwPcp7+7SGAg+Q4AoxckyqPPfp/YmKW961LhwlCYD8GZ4D5b2IAsFDFJATNMI5ep/VxSF6/SBhUjzTIxIDn/zPLmv+geo+f41+8Vj+Pvf+7AX6Bpt757HWpa6BZ5goh0aTcxAmPpGWRJfea4TFqzboZadw1rsNJ9dEey6k4WsTFf/FW/faX/w3egVuxHc2AnYBiT3Uxw84V1w4kC+Gu0DRXZZ/NQFVGgUlpFTjqPgBu4WPmPhWUxYDUqQMUgg5qJ+HhFjhmFhQSxj2FTx0ehAFgLglUxmSQtZIvvEqlDGaPZT6YiQBBSJISw9t+o7q0OPhppD0nABXS+xZhWILJRuHLD6XHMwCjaJxlmuFB04roBhrpJrb8EhJZg4Ce5HjGQ5OGhQEOgKaayOTlRYgarD48lJ0oCeZUh1UUWlkU5Rj3fItjEOQ6+OAXEUAY6qqeC+phldDpOkEL46SaOG9iNkNgiY3W430he0D79NtGhwQYWIBgIcvwPTtzU0/3CWdYD24FcfOzrZU6fV6TQAj75Oi3IFjwrSZiPDAyAe/L62fKirMeF9aT3tdKV9zisMLZs+nENCv4Du/dlpHEBU5UYFKTeusbnfecYdUKmQ6YH30ja9+zYYGynby1A0KMqXsmJqZtYXFRRsaHLYD85OyTyKAE3XK1nbVFaHVqiYqcpogwR4/kDjozMpDZRsYJKS3YaW9AatY2y6dfc4unHnecGjPsVSK7vxvTSaE8gaVtj7/yIjG5Kemp61UdvsOVCpbO1uyfiqoAOdZ8meBsMqrV66qeL/uuuu8sFegdNMe/trDIpQo8ihuafbdA90bRtYDSkApCACPVLCVesp/n3La9+jkuUFtI1sqhR24dRSqaxFsYbWUo4qsVf43NIKlSd22t6q2urpmzz77vB09etQefPBBqboEckHUoDzrDNjJk6ftwOxB2+tk8CePtj9PUoDtVq0yPGSDw67q8rXhqiKphZmGalSlmN3e2rDNtVWROkxTMCqPAm1zc93WVq/ZQLdjxw4fsjHtQxBwVZudmZVVwNTcQZs/fr2t1dt2aWnFvviJP7ILL78Y1mx+vVL97vfU95P8ShLQwfGwUQk1RdoZZEOiZz68cl2B7d7rdBmsxQSP/ftoRvZs9sCEfhT3ABLp8qWrHp5MvgTNXdgIUdCzVubm5txqgyDwGDvlz3MMV41PsWA33XyT/cxP/4zddNMtWg80cV/8ylfsS1/5on3qU39q9Z2aDXSLhqA4p5i8sKUIH1A+yrGjR0W2Pfn002pOcyzeLXCcqOgpeAHCBrAV5AzCosf3AicZ/L7y73K839Xg2LK5OorPxGeA4GP/oeHjPJqcnupNk2VhLrIES7/QEItMq9dta3O7Z0k4VCrY9PSU/W+/8s/tvvvfZCOjk8r7oNE79/Q37fLLz9vG5pbNLhyyN7ztu20dP/w9s53tXasUSvaH/+/H7CMf+U2B7Y5Qcv99mgygDGJeCttG0xU0TIgM+kLM6N4AACAASURBVLRaNghuGeLNkArXaBwSENbVA1gNctGvpo83C5AMWyj2Wq1N7eXuae57EPaADlCmby37dAJJaVWRTYer3CAUnGyhcee549+k+l0gBuChyHjeMw2rj9O/5z3vsR9/3/tsZGw8wCCTCro4gApPrJ9Vqw1bXlqxnSqZH25vQtP+9JPfsn//kQ/byy8+axUYQsjuAh76jOK35a0+NcUETcluvf319lN/43+0dnvcnn/hor3+3tsUoJohppBa1V2ClLes3fYAcIKtUY/WqhCyJSlvsbCcmZqwf/Ovf8WeeOyrttfCDtJVsGnBpWtXLNhb3/oWe+973+v7L6CFCEo+kmdkyXNb53rRRseHtRdzfwFH2aMQKnBP+B5UvisrK/brv/7r9thjjwXp6UHQee+5n6mCVe0Q2Q9SkiqsOvIq8KRGXRZh2rkfa2KRc426jrOJuk6gQQTXBxGddUmq8bKGUL2QoH0QYc4SOwnF+Y/1I/eQ/QVSYHN9Q2tNjSy2J3H+yBM+lIr5c3IPTQIkf/W6c1Bn3V133SWCCMU2rzUxzrl5wMqcmXuo0esCyprNXVtcPCQgjpvSamCHApFf1STU1eV1++M/+aRdvnJZQErv+SqgJOXZ8TBiAJZ8NvQcqJn2BjMzd9L6SYQg9SPq8Mh86m8L1Kz3BSqqAe2N8TsAqv2PrI829l4NkanN3R2RFw6E+H4nYAXyCXA8ySImIhxCiXBvt1Z1pWfYAoSdoppo/ay0bAoPfiguyONBt4Pg/vJ/kJDkftxw+npNjZY0vdpRvczkjr+SjxxB5mDptnTtqs5X9nYIceozQFJquayleA8uCvJAT8QrAMVLV67p2o/L6sltUng+CJ2n5uRejI4NC8RkAhWL2PqZC9ao7tr8wYO2tcVUcNM2NmtWrTc0gcr3njx+lAQ1K5eLsnpUsK8IRm/0IU47e67U5fPp/O35gztgo0mSEK1oAjYz0yK4V9O+QTwk6IKNk0LqFUru+y/7EM9u/p0sZxqcaa7qpaZzMQkAZluT1yi3eXYEfJNfRpiyXtd7DwcxnJzIXousJGo1JhFbjV0prWcPHbTG2rLVtresMlC07c0NW1xYsAbK9rExERVkmy0eXPQJx+ERXUMyvGr1lj3zHESFT1S0qNvpRSJzjZ9LVgF7qdemTk5Tf8g6Fp0HoDV7prLn3LJQ5DeTB7KMcbtKXS/slxo1GwySolPf0kSFxDfFin3uc1+xu9/wRnvymedFVKxvV22n0ZJ6m/OI1yFfg3ro5tfdopwEzkfAK8Qu/nxjPRtByp2ufe6zn9O6UK6UXsNzEjXJNlBUDo5sXzWx53Yd7D+p/M/7I6VxBsCqF3XltIN/0tZ7DhNt4gBZPVgYley7vusB/0OBtW6jTD2oDBEm8wYKIpxq22s2Ply2gU7DRktme41dPWsQNOXysH3r6Rft4rU1q4xNWVvqd+9H6dO2d6oi8ZJshXyAmEVskGuRZ1eT/pq8d5CV9bWf50Jw96769ImJMeV/zMxMi0Dke6s1D8Tm7HMHA59WlzhrZER2Q1mn9CZXCj69z5FCz+kTbj6pyL/jHKDe0+QikxCqh7wmouagPlGdy/2VsM4FgtRcTM5Sh/VA4rBNAz9IRTK1AJ+J98zzK7KQe16taVooBZm8X4Bxn8Lzfp73x/k6PMqehbiDjIiK/q3qgHCVYAKM98c14pzxvYfJlSE9S/Ru7E38tyZWIZMgMSBcJGoKnCLCer2nD0FKy5915QilTSWTy/Uda9erspocKhVVr2sCqOPTG1zvo0cXrbFbtatXLsnWtFrbVv1LLasJ2B1IiYJ6NiYqrFRR/hZEBX0hlSzvnfqqUfMpGIQca2trmshhbQlvKJfs4OKijYyPa+3ofAoCNvctxzG8/8tnT7kwQTopBD1qV75XBKF1hV0lOJ8YR2YZ9vZKNqFw2OjHpXo1RxIA4cjh1ktuT60+t0sgfU31vIBlkRoQUez9YYkp0t4n9XqfLQgO5RP25XVpop6eS2u8or1QWFzgXN4X+hSF//x+w6dvIytiv2Gv4fPmWqeXcZLNuyBl3whLcRKFujV7EfantLDTnh0TqSliFZmnvdwJMhdBBGETglt/Jty6KgkjnwLxNeIYnZM1iVFpEt0hPX3e5z8z1yuhbnv3pixcZcUly3T/K71Xkap+Xju5yl7uNovCzuj9YlLGJ4Xd3ULi58ge8b26r2LbH0ju/aF/FhcU8+9yL+D6eT7MvvDOz+Oww6I3iEwb5auJVI1M2D6RGj+fmtyJChwifFLEpzIiuxaMLkgsWXIhOgkBDJ/3NaKiv+p+7b+/I67ADZWSioIExJzho+Cqa2yW4o3NNwFhmieKTgpqbzAGBATSyFD0oZZlg2MDlz87kxmVsoBVeYgzxig7j91ecefMrisPe8qVGA3mwZdiIcb8fHPyTRpVlUZpQ2Xi1inu4ZagXIb2eABTwYoBLKpRjtCpPMxSDeMbkYefaUJCHpJeiEu5oB7OQUWpq2KMjs+QExe8Bwpp3qiK2wjZzokHb1SwpnHFJP6unnHhFk8iSHJj6tlJ+b9xT8cIzYwmiddzj00/3Fx1FgdCbOypUOSA5H2mSsHJlTw03C5A4EewvT6x4oeHxrRpJGiSWy0RNdmMMcFAYco6gJzw4gaGGMLE8yuwf3rju936SdkhQaa4fdWe1Xa8ifUCdZ+oEKCjADyKebca4vOxLkUcUdDji9ps2J133q7X3dxal5L/G1/5mg2X9okKGqsDcwsKCkSJN784o4KQUXbW7CbgZYRZQ1RwLfPATzWr1POdopWGijZQ6aoZrnRLVmo37fxLT9rlcy8pdFghU1E4+DXFrqLSC+h2X08vqvksswdmbXB4zAoUPgVCezeszhRSKO/KMdnEv7ty5YoKQNRrR44cUaAhyquvfOUrel6wfOKwloXbtxEVHLT9hFiSKLyX/Ltskmm6eL7luQ/QUcKCZ8hzQxR+t68GcZDZ1eIQFYz7YsnGGD32TwDNb3/72+3Y8eOurmLdovrpDtjhwyft4AKKzZx5EpQTyt2ubW1tWaFctPHJaT2HKN64H3j8sga4JrX6tggmvL0ZnadRITSO5mF7e90uX7poK0tXrFWvacx5dnrKQQPCmFGrDg7b5OyCHThywqqFsl1dXrXP/Kf/YCuXL+r7+tUSCehxTVxVua9cz+LXQcB9ssKn0rzpSh92WSmFil4NCgBSKcDoAPZEWvo7UHiiWwgM2IkTJ6USX11Z86kxQukD0BJYSNMGacTzJSVQBDn2qV/8KjPpU7B3vv0d9mN/9UftwIF5Af5PPvec/fGfftw++ck/sY2VFSu2MR5wYpl9oLVHAe9FK5+ZJhK7B0AK7lfmcCRR4VqwUEwJyHfiLMkxrovUoWFHo20nwt/5Pu631JsKvPd9FeBO9z78iXnfaS/I9ySxyevw/Oj0wPcVZS/TNLu77g3a5Vp17cabbrZ//isfsuuuv0nEphSNG8v27GNft+2NDXvqmWftb77/71qtW7StZsd2sbjq7Cl8/AO/9E/s+WefdgW0POn7iGrsLwh6i/OV91gpu30Hny3VYbnO2M9EdMc18LUXXv8xiaLGKjzifcKB9dMRMazJvbi2uQcBoBMgnQ0Ze0ASPln8JpjMr1m8q8FQbpM/a3ntHRjzvBV+7U3shcUhWUfv/Yn32g//lR+xTqdolSGf9KoArpSwVuR1PbeKKTH2YRT7sprY3rEvffEL9ocf+6gtXXrFWrtVCRRokt3HlywmMpSG7aabbrWf/dlfsFJl1l46c8XuuOd27VMCoDp7tlPdFlFRrW1au+XWgtQ3w0OjIg76iYoDQVQ8/thXrduCiHXFrEDYIKlPnTqpbIqFgwftxtOnbX5hwesJ2Tl4/QEgQ53BhA8Kbs5JGu4mobRBYvD5s/mEoPjQhz7ktVEo7r2W8edB04l6r/68kHPTu2dMV0AwE5IdmVT9REXeMyd8awFmu3cxn021TFhJZQZXklW8lzy7sjv09cOzyx4e1kHFsH8KogJrCSbalGum9bFPVKQCNBWUueb5NX9u7qEuFvGpw9tvv91uv+N2TVQA1s1MT9mB6VnZjUnoUK+JqGi3G7oneJFDpDTrLRFSnA2bW9t24dI1+9NPfkpTNApg7XkVc5pBCLinfU6cUFvpnBBRwXPoYKO/f59WcObFSesUe2SToJUTdaP225xoDcJgr9tPVHhzTTYFytgG5BpZXzH1m8IJkbD8e4Va+96eNlW5Z+hcFwGVRIVP8+rzOqQSYZAFnN388/C9lX1VMqpyPj/X/Ojx43b48JwNU2uJLNwnKvQTuASlohMVV68qnBXlM+BpZcgtTFQf0lcoIwv7h4quDXYSZFYhTFq6uiTbOc+kIFC5bWtrq/q9gJqC18wIpAoDFSekLl2zzfVNO7iwaC+88LKNTkzZ+tq2nb98RYDw6etPiyRtNmt2+NghESIArqjaywNMeLp6mnpVYiC89MO+Iol93rDO3pie1jR4CI9U24XK2oVFoSYN8h2AQgrW8L1nb0DBrjoqwE4nKLw243P6/k+4piu9eYZU68gq1ms1KYmZbJUKmQl5F4vRH7mq2gU87WbDhrF+2uvYJNZPWIgyCVwwqcwPQl7ghT8yrAnBFYUsH5MIgmwCnp+h4XHb3KnZM8+9qEwxERUC1JwUk+J1YEDPHhMZR48dc0u6ChPxrmpn3ciesYu4pBGZAk7mU7/LglaiGD+7pdAuF63YrdvwQNuKnRqePiJx2b8/+/mv2j33P2DfePwpm5qdtflDh+35M+cUeM0Zgj3U/MEFTdXeeNNNyppiL/UazD3++R6ICSYDuS+f/tRnPHxeuRX7PvOAUbKTg4jWOJMTQ1mb8fl43ezzWAOpYJa9nMQr/t0+iKN5WhcaiPzbtcGhAXvzm98k8YeDzV0RllicVYaGRKgDeDOVWC7t2cRQyTrNmg0TG08unBV9+rhUsSeCqBgYHrdiZVihycUSxAfWmU3ljQhMFTpYVL8gm9DYHwT6yXLZvfuZaEqRDeQP0wESAQ5WbHsbW6lJO3X9Ke2fEjIMFAV2p8gQ8g0LV/YK1sXWxpb2dfZ81rAAP9kslYVLZG1Nj0OvjPVS9rGeE+lEInWuC/h8EsNzrKjrWGvuBkA2xPjEhFUiwyxFWjpDY4oCYZN6Hb1DFyQo4yimptxSxyeXfJLBxZo8d7rvAoGdqNYeu9eVTWFOAZDDoQnLSkXvh9whSAu3xKurB1TfFbbUft2cAKF38r2bE4qeIdaRRJj+HnSOYqVLPmYDW1IZbdpeu2nlLpPQLdtaW7Nuq2G7Vcjwjo2MlCWAgzA9uDBnc7PTRibM4sEZ29vzjJCp2QPaWy9dXrKr1zZtp4790661CyURFSxlzkatI1lvO8AKyehCF3/WyYNTRubAgM3Mzsj6SdkTmvbPsHoHr9kved7Y/7SXSnzZlBAqn6nMClUfGGSRLMxlbeY5HkmgZq6l8B715D5lrSysqLH5uQl0Axjz9+p1w+I7AWpZHxbIYyU70fMz0zaJ37N3s6aSlN8XQvjPy7wBPpdb9HktIZGOJnR879P9E/jOWvLr6OShYzh53XyQJu4/KzAEs/o8vckN71O1tkO81CMmIvRahGmA3t4m7dtz9sjwIJDZX3O6J89JnhPlKUU+C9fAs2p7AWVeR4VVnjI/IoBdeEDmviqEfM9e/Cy5lf51+nuWPfMksKkk4zXZEXUy+yPXXwKhsE3vYVt8NrmZRCZH5ND2JrB6188zwPqnS3pvQkRTTGOonvV8LXZxTd5EBkjiBLLawnJZ9XxkisUZkWdHirQ9o9a5Et67eqzAGT2c23EW7oPWR9x/SEvWU/bgrxEV/Xfrtf/+jrgCt2n0zvMMNA4muycHJFSQYN2RXnMqZhhL8hAnD7hyZX1+sXGzgWoz6qA0CS/ymL6QamVo0MOFIxgIIBRAU825vO4Y1YxiSYoSVDbun6cfRpPcU4j5RuzNOQV9gvzuV5lAisZCo6j0A4jj24FF+cGGGgaFQY5xyq9Wo8OMYzorK9CeMB958/ohojFEFBEoJJuunMcaBfWXACJZQbAJefHGVz8gR4GlxjasY3hh93N30FfsckyFZMCl+9c6saFDMdj4HoFS8gNQhbLIDd8sk/3n7/g999AVK+FZzmEZtLLG/gMMSTKjdwDKzziuX3lAa0ifqeP+gLLlEkFB40fwGM0YhUzL7n/X2x3IHkIV5ptzWktVdwiQ9mwTfmZOVHDYtVCaSLnkC46/5/u0TrGhwuO01bQ777hdGzdExYXz5zVRMVyq9CYqUJBg/XTo8GEV5nMHZzRRMXtgTk39+vpmLzBup0pgmwf08l6TWNF1bRVsYKhohVLHavWmDVrFiu26nXvhW7Z06awawgT9HdRx9aKU1COe+ZAFVl6P6ekZm5o6IECVCemtnW1NVCj4l+JeikIa2Y4U62Rw8J6YVCgPVWxjbc0eeeQRAaJ4qfI8Qg4yiZLgbxa+/YWdg5x+P5UPkiOWAqk8QBWFGqorMjn4DNje+GPoKvgEe7hOPBPlQVcAQyQwlXP27Hk7c+asvf71d9n9b3iD7p3Wqz5PyWZnD9mRIydl9eOAtu6yj2yXiraxuaHQUXIUqCloqj0kjLCxpq5TrUFjGiG0Hc+ogLTYkV3WJTt79oxduXTBqlsbdurEMTt65JAKlypNeBkv7WGbmJmz6cVjtjc0Zi9fuGSf//jHbGd9+T/b77lmqaZN0icBYQeCktB09Yi+PwtuiqkY/1TzGq4TKgY9Idyb/wAl/Wf5+ila7Efy2h2xmekDIoKY6gG40v6YtlSxhwBsdFqusOkHr/NDqRCyrsCfG07dYIcOH7Uf/fEfs7nFQ/YHf/yH9h8++u/t/JmzNsB+DwgdoLWGgCO7IBulHNEXSRLKmH2igj3Zp0hY3zlSzPsVcB9NhivN95UjUpUJlPE9OK18eP8ZOIj9ANcXi0HWFv8+Adq8HijPRfpEYUvTDFGB0q/biXCzUsXuuutu+1/+0T+262+4UaDKyGDBVq9esicefdReeuEl++/+h/fYxMxB22m1rVpvWku+4gP24d/6v+1jv/9RWbb4tJ8XzCJ1UAF13QqBBobPAzDCVxIVeQ35MwWuxxrK56v3OcKKR2tCYGME+kqx3bFm24ONkwRJ4AyF6MjIeM+2SYCoAEPfH/LXPFNyfegckqerv6ckfxJwVeMcREWeW0lYjk+O2M/87M/Y29/xbms19qyImrDsggb26xzBpqZYXl5x8Ft9TclWVtfsT/7oP9oXPv0JW126pJBhFMIIJPz6tMw6TVtYOGg//3f/Z1s4eINdvrZht9x+kxVlGQloZyLQAUx2atsCXMbHJ9Twjgy7HeV/PVHRVbDoD/3QX1beDmuca3XyuusEgvC+fMIL4M33RYAP9i8ecoGKIioy0JzpC8iuuv3Gb/xb+/jH/8Trh2iYAaPy3gO8cL1TFZiTUAlGo0bmGRKBoVXhopO8x/k8sG/n9ppAfD9R0U9U5frjZ0jRFQsiiQrPPQjkDaKi69MAOisbTYEbrHvZCEVjJzWbb1M9q4f+86OfqMhngz8D2Dp9ww129z33yBYUT++52QM2OTntwc4ivFD31qRc5nsI1ZZdR5PpFc4CLAG37fmXztofffwTInlFOIe9gQtfvKEV0NWX8eUWcfgoe86OkxQ8M26zpsZZgdVeF/Y/y7qO6fEcZ4PAwPgfREWPUJWgw7NsICtatS1lLMj2I0QNvb3QTeR6RAX+Sb09gp+p2tDPjlSQCjTofX0bUUFNzO0sey6Jf6+TMamOPX36pE1OjPk+rtwmLCAC2vs2omJ0eFD1B177SVSwt7PnsPZ4T7LMke0NWVUjAhKvXVmy3Wq1R1QAim5srNvoyHB4ODNR4XaZ7Cf8u9a5i7a+tKpnu9nqKjNnaXnNLl66qokbgpTLlQHb3F6zyalxTVRwfmprkw2TK4chFfncAOq6lmHdIXuqqAETSNdZEtk+sijCplPWFfv2EK5C92ckQU3dR3L3YrLON3r/f1nTU/OyR8pLO4QKCVxpvcUac+IjQtkDyPH6njtHH9WxEYKGZU/atZHRYRsdH7f62oqmCkFeqM8WDx1W3VyqYPGyYpcvX7JT151ya60ylit1G52YtvWNbXvq2Rdsbn7BLl6+qmwR9j0IKLe3K2mKk1xCJiqwxcsvn+LznlKglqu+fJ1B1vQseF2lK4JcrDSWVR0bGmjbSKlj1fV1mxwb13TUo998xu669z77+mNP2uzBResUi7a6sdMDRX0fLiqr66abbrID87M6m/26uoIV+yXWs0izwoB94k8/6URk0dXT7Lm8FwAi9vKtnapVKnjhe4aCwKNQO6c/eloAp3LWI4NcgaxnXZMlvD71iAvEmq2acnfe8pYHledHTcH/OkyQyGO/IbKCdYadz16bac6OTY4O2aB1bADbOPUanlX1lYcfs+36nnWw7trDipK+0tG2ja1t222hbh+UYIspP0j1BMRZYy6ac1CU8HqtNb1X/Omx36zJfpO9EoJzdm7Obr7lprguTvpCknE2Umc5+OYiPOp0AFgp1aO+UEiv7akO9wlQt+7iDFOfnFODYSOm9Rq2LpJsUFNoAsJFLXpOwwHBLdZM51OqkzUZKvuesNss0IsylYFtqU+/6IzXpI/nBElIE2I/sIy0gxLoLIs2V64rz6uOyHNCvYme+SC1mL7kdSB6NHnRCfsWkZP+d0yXOahNpplPSOz/fAeRNe0Tosu0zu4ptiFuyqHeZlJsd8cOLczYxOiI0WHRD3D+MSm1srYeOSFlCeNGhou2eHDSpqZG7ZWzr9iJ6066kLRttl3t2MpazVY2atbqDliT55nJMPb1AJiV3wBmIfLbgXnOX9Y79l4QSnMH57UPJbbQ/yvrm2eOXp/PI6I4yB+uAest92Cvgdm/XSDnIi4XYfRshEJlz2tmvZs1h0/I7xPLvu59T3VrOLdR8j3W3SqohV274niEMiwjx0h4SoQb5xmapEPu2VLaR93vdbKr89WjawqDOsRB9SQh5L4RRIDbkbl9kP99WCgl2C4Cjc/qE9HeN0VtwMFA8xXCCV+/kXcQz5CmqPostwSqxxm0L1Lat4pKYi8nQBJbUPi0HBeKmpjUNHjR8T2uIyA7z16PTNF4RrqgdO2lfqLiu5d6/YlIycDSfFLBz07ecwp99byyv4Y1dO+M7bPLzEooMaWcNteZ8xdMVPQVTj3Roq+B+P5kbgJ7TJuszLzhs7KekzDSWRD7ka/xmIwEA1QG2H6eBX+vfq7PIizrSp2dHe/vXyMq+u/Sa//9HXEFbsIvOjYOPlAGFgMaoNrwsCYP4ZEnPKN26sVC9bznFk3ZEI9hySELD9+IObR3YcX7POyycNA2F+EwbFRs1Onvy/ug4BiuEFTsygABtbKY8DwCbyIA5HlPaLvMPWcV0DYoZQF/TsPKwcbr4JNIcUBgr8iDsK3xJsSBZYELXBcRHxywDScvODQVzujKKzZn/g4FlL76pic0lcCGG96bFE0czmxSCeTwXnNkmE0mi6dsaPzgTsULyocRKTN4DakumPAIC4X0UQR82We0aS4rCjrzxsgbKBEvMVbmAKIX68qIaDS1iQosEXvrKlDdTzbkYKq5Hs0630ux5E0H39tskcXA5EdTCiFUIhAVAHbNNuBjU0RFEjwJ8PYTFRA+KEt4z9y3tH4ixLGnXQoARoHlMfIJUcHPxfoJkmx9Y83Onztvj35tn6iYwvppr2tTB+bs8JHDNgzQO+fWTwrTLpdtbX1DhYIsg2KiQsVwWGdwf1Qgts0GKoRronBr2lBx0AbaDXvlhSdEVNABS90WAcEq7iOTgubN/TF9ein/HJCXkfohJmx0/RyAb+2iQmyLwGAd8VqsvcuXL2uyAvBsZvaALS9dsycef1wkxRhKXo1dV9S09ls/pdIrAUkHp/yZTi/PBMwIHhSYMIAlVEXWS3y/JrFEHO6rYLmfCnnn/Q/wPNYM72uISIJiCYnl3n7f93+fQrXVwOu6VGxyas6OH7/eigW3k/PCwotO7B5QO9UadZuYmlYTi8pSz2bLfyYAHGHuKij32q5GrdettrNt6+srdunieXvl7Bm7dPGc7Wxu2KmTx+36k8f1jFCso/5BzTk2OWMHDp+w0tiMffOpZ+yRhz5pu9trfcoUL1B9CiWUMH0WLT3wNopG9s5UQvjI7F5PaaPPmMq8UA6pMFYAvQPYSVLkfxcKkK4d2QbRxI0qPNSbG8C6nqpDY9iuvuDZ5n6xp7ImuT/9X7SHUlZTnHfN5ucX7Rf+4T+wO+6+2x5/6gn7t//Xr9s3H/m6FbEOCDUHPxOfXMAPvhJUEFiaivBQ5+gzBAEVl0UkRp43+f18X/rP5pmQalauN/u/nqM9E/DAfQes4guFGq+DreDE5GRPpSrrvAx1i2wfAidF4KLibDSkMm83UVAz8o9qt2x/6S99t73//T9v111/vZUqTMUU7Mzzz9vjX/+m3XjjzXb6dXfYTrNluw3UW+zLBRFh//QX/5FdvXJZ90hEW3juttlblVngZDXvFUUo1zHXTBKGqSzi+/LP1JgkCRVEha8NwA4nGkS+Aw+IFHbAM7+8SfN1kwr5BABcWebgaq6znoo+J4mCmOf1koRIJbAHKbrCNxtAHYkKG9zVXvv+9/9du/e+N7rGrwCASh4WIISf++wtG1Lgd3VWG5YfbbML58/ax373I/bYI1+23e0N22tUdf42Ol0phAfLDua94YG32Nu++902MjJt19962ooCYPB1R9VZs9rujiYrOOPYgwA6R0cmpBTmOeZnX7t21WYmJ+z//Fe/bE8+8bB1W4D6aVPk1/jBB99k733vX9MkG+uPySGyuo4dPyGbEx+hp9FgvaLmpImAnGiJkGDCDLBGoZmRe3XmzBn7xV/8RdtYX49nwhtuVyUWQwgATS45MgAAIABJREFUYOEWARIJsO/m9GMpsoSGsNUi9B7MdX/CS5OaES7vIbZee2lCUArR/YkKNUOydupT4cc+1E++JjnmoH3B9gqojNsCKETAN1u2tYkXdk3Np0/45OtGXk4Q+LlWEtzn9WR3F+udNcm5d+jQIbvnnnsEhBKsvDA/q8mYgrl1gRMVTKT4FBl2jlxDahXuO8QkQNy3nn7O/ujjn3SALcABnzHwcXzWJWdXPpf53Em4EUTZgHzgnahI4Qzuy/m9+Yzn85ekbP++2yP35fIV1k9dBBEADGGB06jKsod9KsEJwDR5cBsh1K7sFlgQZ0kUtj7xGyGfbtHgmRppV+rAAmpWzkzqVTamru0RUdEjx71u5N4hvrn++hN2+NCi2xTizx/WT1otKjQKRpj20pUrNqqJikEbZSoT0JDnNnLHJDAJRbKEPgrehaioiKggb4sJCrzSuXfs7/ze4REXs/C/8uCwssbK1zZta23DNrd2bGHhkKzkOnsFO3f+glUGh/W8Mh0FEIwt6N133+MBr0UUzW4vBqhK1orI5RBTcU5Qr6E4zhwCnyLytSJwJLzl/fn0SQq/Vw6e6j6HgjdrLxcaeXC0A05OWipMs8v5ti3/fu6zfN7D9ol7zWsIPA9wLteUW4b4vo99WRexWLdj46Mjtkfd30LYVFDmSIdnBWuc0oAtLy/LM94nkyvKp7p88aImENhLUPNvb1dteGzKNmt1e+pbT9vho8fs5VfOa6KF+45afGp6SgHEPKcrK8sicFmrej/xntNmx62gHERTr6Wzap9o897AgUHsaMZHSzYxXLRCq2qNnS0RFZsb2/bcC+fs+HXX2/Mvn7fZgwet1mrbxSvLqqGxy2ICYXxiUvXCLbe8zsYnIerJ1aA3aWlf2a1hIVRWP4Al0hf+/CEHlGIPZeqK73d7vZKmsrBDzfNZKuzIC3TiwkUsTIjkhD6TfZmD4vtc9HZh/YSKnomKymDJ3vTgG1RPcJqrLA/nAGUBxFk/OlSx3dqW8immsEErmrV2NlULqN+rDNsjjz5hu+2CVZt7NjA4amQ0yi1hbFTgdLP37DrxxT4ASJ8T1limIvyAZAD4VI8nezK3LSarg/NI1ljlkk1OTtgtt94irIBzk3oAmyYmJLPXY28DW+D5p+aWSI4+mf1E3KcDcp6R56BeCvd80skBWE0Xayrfw4npA7EZunr1am9aP0V61FwCAeVO4FmcPrFR0BSiQHSyJHjWw86H/8aSGPEhzyTnptT1Ef6ctZWflwN6Pepqrm9lyCcU6Cd4vnieNUWpCQ9e022RAe657pqIIi9UWY0RuB55eFxb6kQPEvc6e3CIAPq29hfyESGYWGfs79QaTNE3EKDSWWnSadcq1rLq9oZtrVdtuGQ2NjIsa1OejfWtLU2eHDmyaKUittgFKxUQmrZFWpJDwppfW9uxZqdsaxvYJ25a20rW6ppVEZBof/ceQlbZYdfN3uXCzLZnlXE/ybFZPGhDYEzce8LOt7Y8O0RCVcdDhKkwqRFWPqr7wipK10616H6N69NNDuLLBSEmPKo7O3reWDtJiCR5zDrjnmQtm1gVP1c9GBPVkTGkiWHtU75fsa6SKNYEXO774UahIzHyJXn9nDpMrEcEQQhoNTUXolnuMwLJtGL3TCjPfcnzI6fvsq5jj3KLVg8n700chADJIRyvw+id1ZMGjpAkBO9XWZZhgZ77sn5235SBeqrAMrg3boHn+4LOuRBD8N6UaQrGFEC6zsVwxGCyQuI02YQjggbDAV/zrxc/sx+mfePbV3riY32O+Ka0DcvaMa+Z2zRG/mqQE+qR+siTxClzNESETpBaOmdj4sNrOc8K6YnrVDz1icwiWyrPYr1H1nJgof34oguPHSPlfWfv5USW1w655ymTt69+SJVPTpJ4jp0Hg79GVPRX16/993fMFbh13BXaFI0A7n7QudrEDxcIBA+UFFjb9fAWiiUOYTHBERQlv3E1N/5QZ0aDVA7xMCnTIlhoTWPEZoJqlQMdpcHGBlZSbgPFIYs6nAOBoo+NrxbBxDDz/Ds2e4qUiTEP2hN72/BcA5pVNUP4lYZX5TZByzQEGnNn44pNqC9DwhtuV/6wAbBhiSQI0obfa+yP0VyN7PnEBV80FNqI4tDqgYKR+yBlSHgSpkLKN0QvQnxsjlwQGHYHKjnAFdwaG7tAfI3UhVI7PB4prnWYRkAPmxzekGyS/DkEDEUMr0lDwetkgHpaPFFw9jbsCCjLSQIX4/hnRfnG9RDIJ39hD5/CegGCQl67hEK28DRHVYZVQdvufftf0nvRphpKfAoFDrzaDg25e4kmGC6iAqAFD8CwGkkGXlMZHQ8Y47NR8BGmTQOytr5mr7zyij328CM2xETFdaeUTUHzMT0LUXHEBitDNjM3oXDiAzOzriZjoqLdNoqb2q4fpKn0lgowbbbIUqiY7RVbCjKGqLBGzV58+hu2evW8ACaurYqVfrVy3If8s1SPcz1Yz+PjUzYxMxU2PjRpNJR1a3K/yyWthVSTLC0t2aVLl1R8zM7P2erysj3//PM2PTnlI9VAOCpa3F4qAfM8wLnP+edOVoRfcEyt+CQA67+iiQoOT/zmuQ46THtK2f0gMNYURRYqIZF6BK7VG3bp0mXZP1GQvu1tb7PX33232zhozxi0sfEDduzY9QIXv52oQD3L816t4xM7peKPwh+gAZIBVbSel4EAmva4btg/1W1zfU0AJATFhQvnNFGxs7VhJ44cstM3nNIUgQpRgFgbsMHhcZs/etKGpxfsC19+2J765pesXtvUfUyA1n2G2RuceOwvTnpERYRqJ3Al0iiePRo/Cm7tEzQmUeBLB00OSxpzhHoiwWMKbUAaXzteUNIIeNaN79v9YN+r31dHvqo+LeNK754yNyYqnKgo2PHjJ+2XPvjP7MDCgp27dN4+/OH/xz73Z5+2Ij9DHtKudMyJCk1OBWjSU19TXIXHqque/P065QzQuj/9IRVTgD0CDmPElV/TSkHngaYQBvWZReLJHsQ92wGytJ8NDwmIZn/uTVVEDkQvOD7sTwqdfcX51o6rv0XGForKjPnBH/zL9r73vc9mDx9yQLfbtUe/+ojOhgfe/FZb28JqBhsF1IL4EZfsg//sl+yhP/98j6DlHgi4AkRCpRtnqUgZWU24YrB/nxDwG6BNNlTfTlQoV0bnEWvQwUQRP1rIfj/6J7Z8gqstokLncJw3+brZPAkkjuuff6b7l2PhUVznv8smxEEEFy2oKYu9HXKa/ef4ieP2937hH9gdd9yNuY6UzLKZkUUWzb43lgBisnLAl5rM0HbbHn3kq/b7H/1tu3LuZWvXtnS9a03U3Hs2OkyYLgDSsN151332lre93e64/14bGMTyDpuokpSDnEs5UcE+Cyk8IqLCJyqYSgLkmBgdsn/5y79kL77whHXbDnorf8DMZqan7Sd/8n321re+Nawg9wRoQ6wcXDxks3PzcWZTHwzpOrrNE7VUU6GgIkVL5bCYQADSsA9/+LfsYx/7WE95nddPUNWeh5sm0NwDwmPiEfC0WB4QWItAg8kKZZ0I1PL1nWdMTnLyGHK/etZGkVGVoGH+mmshBRMCs3JaS6AAwLefKxAVCvhURllbJDEkO3WT2xY5wd+v7M8aLInK3LtyD0jAl9qN9Ys14t333C2rQ/JkFlFljo7bQJFn3YmKVgtA0S1wZmYOaE02ak2BbZxHu7tNe+yJp+wTn/qsctQcYEAxGERdCQVoU0CZN6j7hI2mIko+8q/PLUW4ky9a90gp4jjIz5Z7sL++T5bkM5LPPgPEeW4UuY4il32qYq9ZU7A2Z5mU2IA2Q8MC6ZAStpKowMZFJXWcASKy3CLMCc2cmnIbMbeA8M+iPQZVuWrhrrWLHQkTXNEZOTfy5EctP2M333zaxkbHNVGhobqYqJBa0rq2vLYqooKMCa4/kxUowQH/WXO5p/N5ZKeRHu3DoyIqlq4uW3V7yzMuBn2Cm/2d4HSuCWcHRJVI6rAmGt1o2fLlK3qusHLa2tnVhMuLL56xgfKAvfFND9jK8jUrFF00w4QF4yNDAgF9r5RKueLXiudJop1yRdls2NgpQUTnlHuMU4uxV7GfiNjiHM0g1gCgZAsZQElONCJS8r3b1wvPC4COLOME6FR6k8OAvsoJiTBtnvFeLkIE1iZoKjB1eEgZZLu7VStAArP/0g806wrOHqqU7PzZMyIr6Jno+5hkO3L8hH8ufn/lsmxTb7n5Fp17leFRq21jPzRmGztVe+qp5+zEdafslfOXrKapbiZsfQIEsgKbsIuXLtoNp08rDD3DZiU6K7iAyoEct3vRxDyAbYBdCchlZcUx0WltW6FdtaEiUxVef21tVe3FF87ZLXfebQ996Wt206232sWrS7a8vmnDY+N69MhBAGhdWV2x++673yanJ5Wjh2rb+xJ+LiRwWfkPS0vL9vDXHtGZQC3KPkAtzX1hv5ANsqY/8Knn8/hemiBp1tZ8vrQL5n6JgJK3ik+cu9QXYot77f11o0HGX8EeeOA+Gx8ndLkmsoLzjT6OqQoU+jwLcmhjUrrTsPHhik0MlqxV21Hf0WriVV62rzz8TdustWxgaEzBx0Mjo+ISqZtW19etUBnWn5ElxJQfzw51pBTxshVGXOZKXfZWCAfWO8A42w7gs8iCEDAiELnldTcrE86lNnsiOtICh2y69dV1rTnVzzag6+ukm58Zo+Nu+5tkCK+VEysuDHKrJ/YC1ZEBVrP2uUYQkuTZQFL1i7p4PvmZEJJek0GMDnu+2a5jBU5g1CJ3cUfvU0rmUHkrQ4IJi7Bo5e/yvWZPqol3nqOwhCH3g38HlsE+A7bBrxKHRAamel9NpfgUUdYNAsI1/QsF0NX75XNw7DA1CAmofpw8TyaYEXNCDm1v25B87t26e2JsxLbXr9qRhVlNlFQ3N211acW2txCEkCnmVlKsZW794cVpu+H6ozY+7mLIuaNHjZiwlaUtq7eKdvnqhr145qINjk7aLgIpdSUEc2MVFRa5Du/0ro8m4Nm7NYFV7CMqfM/kS4A3hLzEfY4R8HcSQUUANH1l1pmahsGZQ/Z51DluH8Y1Zj+S+j/EHPu9kGM6rDvWlYilsEJ2gNhxnGaIfBA+afo9lP88X1qHWv+tyG1xDIg1lXubSNicQM76PmymBEbHue21lts+eb3hEx1erzd757ms9cKKnHUABkMvDZndA7OVJeP7TL/7gy6v8tMcaHfLTuy1HF9yoizuWzh7pNWkiEip+V24mvUQ1k/8N8IDsBeJZ+N+KOQZAoPeNELp662m54fEJJ2TBm5nxLOrrAnlnyII9kD7pz/h1sx83fSOlZ59sa+xCM4OJxaf9IhsjeghZZEFoZdEeISM5/eJZArCgdeUVVOQAv4Mu9OJrllio0Ew9EQ00aMm2dPf/ziZ4NO0SZCILI16U/e7bwpDPyscVNJRIZ+nrCHkvKLP7s+RV19+PdQ3vBam3Vszr/3Hd8gVOKZQMQ/tlJcfav3YoGnuFcBDMHKwvfhsSq2JkgpvV8BLxhIpWCplHcZMW1EAijUV77ofQCcLJhRIfUpPfITZ3BUWpdR7AvcAhLs6dCke+BmufK4bsLQrZGNigYM/fl6OlA3jM0ljXBywtfV1rwm7ZosHD9rV5eUe0CeQOw6ntHbS5ttw71SF/AURI18/Dj2plH3z80yICH1SNgfASAALFBM6KF0ZoAyJANrz8PXixoMmfYTcm1Q1z33fy/sBWOGgygM2QzsdTGB8jn/bVrA4B7UUX6HAjOpBP4PDQsAQo5SAGIyfl8q6f6kUczWuWzflexEQGRuiiBWNBkYAU+SF7DZQKLqqF7ICwADliCt8Ycr37J7veVuPqNBhJWDbCaXqtk9QpG8pRdl/iajIf5fWTzSSFNaEAgOur62v2vlz5+yxR75hw2UnKrANYoufmz+oMO0kKhqtlmG7RGAdyhHAJYiKnVpDI68i8wLYyYKq2xl4FVFR7pastrFiLz39qDV21qysojiJCldPpYIH5W0y6glWeIE1JPXf9OwBTf5A3NEYt+sNq27vWKfQVUHNWuAL4Auygus0Njlu66urdv78eZsYGxchJVBUQARsu4PqOUWRo6YJLCdRkffEf+//Exge1k/Do4QXE5JHoRHKlz5ARwAsXrEtQu04/GnAmrICOHv2FU2AkA/y7ne/W2AwY8NMVIyPH7DDR07Y8CAK+WhRQ83M2kTZBFGhZkuj0Khe8R2HrPAAvTLe2mr8G8YEDu9zdXnJVleWbX192c6fP2cXzp2xzbU1O7QwZzffeL0C8pjEEODSwkJsxBaPX29DU3P26c89ZC8++5jCHHsFQ9+kgwexhvVJAtJBeApkC8BW910e8hGihyVVve4AdtjcCdgKxYtTb6GACcVWkkh0DOmN7kQlxCJgW4wAC6jan3JxYTJ7hN6gCE6uixRjIyhWh6XaVGMZNlSswZ/4yZ+0H/ihH7KltWX7zd/8DfvsJ//MmtW68hhy/6ZpAFLvJypYx7mG0r7IL96+n7uTHF7AJWGXR2o/cK/rFhMI/VN3PJNcO9YwwAFrmGdBI/ODTOd4TsX+v/Hr2SnQPABAuPoJqxS+eC0IV8BAnT0xgXbsyFH7qZ/6Kfue7/8BGxmfsGGsAHaq9srZc3bzrbcrtHOnVrW9lvvJo/79/Gc/bb/8wQ+IlNUJmCFtkP89gq/oe1zBR32TqEgQWM2Az5a/igjLNQFDmOsBgCUJIBWqkIflfSsQzg4B0rL+ozlxD/BsyAR+xjrNNa6zA+FBAMv6WQESJAHR/29QQ0udnxMfPSUxZ2BbPskda9tNt9xsP/d33i+yotnaC2uwCB8sOkFOEw94rympumeSsFd++YsP2R/8/u/YztqSAJyt2q51EQrgMx6Th2MTU3b3fffbf/9XftiOnbzBKpVR2+ugdiS/BtCcEGsP+u4nKliDW1s7dm3pmu01G/Z/fOiDdunCC1bYY0LLp5RYY/fde4+mKbA08Sk7txRiYgOC4MiRYzY+Pqm1x33hGsm3WgGhO1L3AjoAlgDycIYzFffBD37QlpeWes1iXltZP8Sa8Z/nzaHWQai3tQcROlv2Gkn7NM1vKjJjWjVJCr1GEBVp8aeAwbBFS5Iq9zUnSLxBzYBFJxsisygmKviMHTcicqKitisgj73GmygaUMQweRZ6U+6/931Az2ivYffPKcUlgG6xKNDrzjvvFIA6cwCiYkE+/05UII7BrgkFrCshAUmZLKzt1FzJ3yS3p2mPPPqYffbzDzn4R+hieIvrs5dpnOtSBfcIo3wOea96K05U+Hr3X7WTxLXI5zQ/E7/vESGh2staz2vefbsDJyq8Lk2iooX6XRPNPvnqdjxl5bBITyrQI5retJSKNZJezU5WZHh2nC1q0uPPIVk0pgNi5KSLT9U4uZz2laOjQ3b8+FE7eeIkfOiriAoBeoWurayt2dLlywJbAdsQLkjx2fVpm36iwglXREpYRvL9FVuGqGCiYHRIgBv7FuDsyAgTSyhyC9r3AeULpYoNMVVxdUfTO/Ua9eOkDY2O2+Pfesq2t6oiJt70wP0iKbAnbbYatjC/YEPDo9bdK8pSh7VJLgDPO/tPWm7s18wmMDHPFSl2NblQ1tnB8+8qfA+B7g++T8sRB95cxKUaPKxgAHpTra26doha1kUxXFNZ72CRE4HC1Du5ttwmxuv9JPy8Vqd/YiLLlO221wRgLVhrt2bry0s2OjqsDBf6vc2tLVs8ftzqtV0bHB229dU1u3blivIGmLSBZAJsLw+N2fLKuj3z7Is2v3hQnvWNdle2XhITtVp+9g4NigC+7tQpn/whaJxchfDnZn+Q3UrsK26JgYUsEy5haVt2goraZqjMFOWujZS71txZsUHqBk0PDdgXv/wNu+ve++3RJ561mblZK1QG7fLyqnI1XBTm9lzUiuTbUD+z/+l54HowaQJprgDqQTt//qI9/vi3IrfHPfV5n9x3hSxDFGkaxPtYB/Vf3YNxv3K/dAAzrVPoF/uICqnHfaqJNQOZjdjmgTfeF9ku7GtNK0sR5OsAAl99qK5B2wb2Wvp1lI/ZZi2UFY7c3jN75vmXrdrsWgVCvukAoCxbrSsVfQuiRKQYqz3qfFlNeQ4hPYPnr6UAJq1Yy5o8kcgpREMQnNMHZuy221+nPsxJUF/raT3spJSLMjhXxkbGdHaylhFUeV/vPXEGk/N9flayhrCE8jpDYCi1c/S/EHluF+XrLWvQ/voKLKFHzkMcaLIh6i9NDpEBsi6Sg15MwLAySVo9u85+QFJ1m/oOf/5EtMnu2olv/g77J/4OLIW922tnFz86jrCfdaFw68ht5Fe+120Z3f5IpBp5eiJMavq5PL9pt53kH+cGwk/VAZy7vJXWjo0OlmyUzCAszpTzC0i9Z8urK+6eUDbb2V7XvlEeYCKmYBub23b48KJVBkfslVeuWrVuNj45by+fu2y7rT0R5dQfZNXsqc/x+l/3U+IBJkhxsKA68Hqba0gmjsRvEHR1t1jOCaoEsb0XSBwjn+Naj8DI2j33whQUskaY/mPaRAA71l1hJcu/US5E0Z85rbmwWtK6jJojsQ329axLfIrCSWQEtAD8vK5PwnQCS/G6SPkyWRf0WSepxxJek4KzsEIKvIfakH3Un5GwISRfaNjXY+LavtY9t4g1rEzTEB+58MCfWX8O/JNpAoXpJ0LQIxuJfZlzTfVfgvHKQHG7SBEZQSDz93KwiGsmIZMINH9v+axlRqCmWcmciTxSriVCMN6oaosQVngQtpMUCmQvee7hM5+cybbQmKjw6ROvEzPXUaLczHHNOjKmLUQQhO25LN81ZhLWnLzzIDeED8YkSNbXbmHuXxIfZOZUby/0uov3zb7N3pqkhoi38Df1CcKYgOyz2RVh8RcQFbwXJ/Z9SsJrrz7tpmrkIJxUzzlJkV+vERW9S/Haf3ynXIFTJS8Ke+NQUlI6KOsbnW9wvTElMioGmXAABPJAVW1/ZFDIxxPVK2pJNmlsNfzgzoc9g2M4hDlsKeYBbDhwBSrJ43HYR8hCacwDjZ8sBbDGPCuD9szzzwtjItSM/+PnQowAQPH0D8mfekCTFRS/OX52YGZGaq+cVFChIC9nnxKgkRXQGaxvKns4+KRmoCEpFPV66aEqVbiZCkAFWtI8ht+tM+A+5ZDNikDFKGqy0PNN3osuP6D2AaoeG2ym5uzUqVMqpi5dvOwFWXgsezEZmyrFZoyQ+tHrGzzv+dixo7q+TBu4OsM9HsXgy98fOyeYdvcoTYBEB6vel2+aHPRSBqAUJjCLkcMy6wk1LH57TFRQ0GNJ46Oue9223feO79am3g9ocrBxTXa2HVBIoiJBNu4jExU0X3yOPJhybJD3g1cqStsTJ06ood3YXBdR8cQ3HrWRyqCdOHm9TUxPG37QC4uHbG5+XkTF1IExfe7JKYiKkgpwn6ioWq3e6hEVUk9E8whQYHsQFQXrFJn4aFmxZXb1/Bm7dPZZG9hrWAW7ij7lcoIxrHXAVF4v2XfuOdeZImVwaNSmZ2dsZHzM1UKttg0OlKSS2abJALAJcJb7h+f2+vqalSolgV2rq6siKgBgeCZENghoc7Cpd2jGwc3PzffWD2YInIwRUggcwn1RHzJ1gkpWtgfhrZrrlfXon6NitXpVDR7qDa7PysqaVHrkanAQv+td77LbbrvNOrL5GLTxsRk7uHjMxkax7YkdNogKGibuOUQF4ds8QxS+gGBVmrK2k3vgqlKSA+ygoNbfk/OxozDtc+fO2tmXX7Srly5KZfS6m07b9MyUtQEkARWbEIuDdvDIKSuPTdmffvqzduncywqjS4A2r2Eqvv7/EhW5D0BU8F65v1KWqNn1cbS2m7v2fmZOVIg8AoSWWst9/tmv1fBLfe3Pfyp398FGXtuNgXR9mk09++nxy7OjkDbNtypxwGYOHLBf/MAH7PCxI/bbv/1b9vE/+mOrbm5Zt4Wq1y2/+Pcyoo3XVYPSZ23kUwFBwBBAK7WSnwcqrcKOpEdsRIGdZEUqrZKw4PtQQqblBXsVewXErOd0+F6PFRoEDM+YrG5iT2Vgmf2SaTAV21gIxFrjvdJUEbgrP2CdJ2W77bZb7ad//u/ZHffcZ+NM7O0xNVe3yuiY7TLVU6tap1G3VqshIGh7a9P+9s/+tF27dkU+0wIpQj0KKZX2HLxvwp7TH9WJolBwJ1GRj0FfhoTuUajxeC6c7MhzGg/9gvYCilyuDwQfz59I7JZ7RHNt9keLXYmzDxQ7GJp7kiYlef7DtseJd7c36gGxEfLaaxhiP2Md7hHAroK7ZZgj33XXnfYzP/Nzdv0NN6u5ZVU6Oe9Eucc/uiKM67y1XfWQ4k7HPvNnf2If+73fFnFYbzaswbQgQcOyRdiTenzxyFH7+//4f7Xrb77VKuUxY4k2Gu0eUcF62CcqxjXBwedjH8WuZOnKZfv1X/1Xtrp0zgrGVKNP2MwtzNtf/ZEfsbe+9c1Scid4wJ4HsMnaQ7m7uHjIw30F/Dois7vLHr0eAdtO7nM+c18++clP2L/7d7/dUx6msl77DbYH0ehwPzLXRvttkFVS5ImoQGxQ0f5cAiSBh0srmJZPT+SZI4Aurq/XBam6LzrQIKu2fUIkz4f0XHaQFdsK33cEkBaoxLxG4D3XqxAVvgd70B81FtNf+1MZ3ojvN4LCvfsszvrXJZ8fQODmm262e++91+YXuNYQFaM2UKgIFKFhbLXrqj1YSqxZrD/rkNnsGy23t/zSVx+xh778tcgU8IwyEd1lriPTptVX7Ru9ekyjbzlR4QC/rNeCWO/q87j4op980aMdXgX9wo99smJ/yoJoUoFVClDsKNC906rr/VBPuwoxJiHZa2M6zIkK30N0BuRUXo/U9Hyi3jkW9kXs9axvzxpxa4jiIKaOMVk1wHrw6RHuz8BA1yYnx2WjMzMT6ItxAAAgAElEQVQxKfs8t0J1T2/EFKtrq3btylWbGBsWqTIyVBFwTD2d6zDVyIBI1N7sT1iccJ4tX1uRUGR0hDwsPzMI0tXULiHCFbeZ4d8iLJDC9MqWXbt8xSbGp6zewPpj2F65cNFW1zekSL/u5DErl5lMKNl2dduOHT0uRf7oyLisjQheZiKInwfQylrlLAB0Zz0LqIa8Yk+tN2xsYkxh8ceOHVNPRA0JEMM9SiVwTlhIuAGwhIqrj6DvJx65N5zJ6gl0DroPve5NZLPJ1lWZc/HnIp9doZnEc9bV5Jt0yTnAQoiJLqZRsbS1PdvZWFUwx9TUtLiprZ0dm11c1H47NDpmK0vXbPnaNTt58qTXFwS8IkYbntDE8Ysvv2Jj45N26co1kwFNwW1KAXip/TXBsLxsN91yiyZWRUxFILHnvTmIJ8VrWP0kGaoeMcQfPM/sk5Njo9ZubtsQRXaramPUzwg9OmZPfOt5u/F1t9uTz75gw+MT1h0o2eXlNRsdnwi7SyyB5gTG3njjjTa/MK9nUb0PQJx6RohCzvuKvfjiy/bccy9o3UKAcj0hKDT5o+wSsvggIlzh7P3IvmAnn30H+DwwfnAQ4qkVJEWSFS7e6ErA4aI46mmEbm980/02PT1pO9ubVikjKGvrTJc6Vx72Plk1VGbKs23D5QEbZhJqt6a6H1JvZWNLFlh7xUHrlgat1sD2jAmRmg2VSnbp2lVrF8j+GVX9rByaciWCe0OCHXULGU+A/JAIWmecabVdGx518kmKdjObnZuxW297ndsURRg1PTOEMf2hQPZBn0Jy0tQnZn2qzSc6EB3y/PFnaSmj4OA+Cx25HMQUINebehAlfuZlpEJez1KoqffPPscFAFeTBJQffBD64Az0fkmqYRFJnSu3A3qxIX+WsyYXaRIB93IGQIwZOUPgEBJYMm2UmVFp0xdK8DzvWW+JxVDP+pnE2vEMD/Yc1ayyNXKSTYRYb0Kv4O4IMcEFJoIDgc6hLiZNddvdWrcGwppm27pt8guHrTw0ILtUCKWDB2dtsGw2OlJRyPbo6KDcBkamZ6yxXbPnn3vFqruITip25vwVq7d4aAas3mpp2qeh0UAHt0uhJs+9Ka2fVNMXCiIqIIfpK9lfWR+sGWpzZdVwoqTwRdZDHSnueW4lBAmbIbl1hJ2P3CRiekFTQArudsU+6y0J3VwLujaaYPCpIeFU9DbYt/HcZbh2ZKRAFqs3YRIwpgewjebLs7d8jijBbmFo8Xup9SVKcHwle+WsBam7EEfwa4qFdY7o32T+Bg4Yg9r/k7ji/Qj30nQDtQ+Eub/+q7+cGOcdMT2VfUf2mbymk+8hXIopgJws0PMaILlsx6I+9Ofczyt+TcyItaxcE7JigmShXhQ/ERkfwhZl7YWoz3szzzV0gv65Tx3ofYSb3r4SlkhuL5XWpE6yhhAkvtsncPz1srfkOmlqI0aH/HM6XqHaOrJ19blw0YzskJyGyNdhf46i1fumyNtJfM1F0UFUyDrMJ8VZr9oHQpiTH+zbJyp4bQl7+kgzfT49C17X9kRimhBxrNYHZJn4PXhfwifftgBe++1rV+C/zStwhMKIQKuw0KGYEgg9MKCRMsYgBeyEjYZjTPhOO4s5VBnSxklTJeVkkdeimfCCX+OJFUaR3ZIJ9cTE+JjCtfKL8TX8TRWqXW/Y2tqGNkQeaixsOLQZwwYcqO427MD8vD37wkvyx0RRRnPBoYxywdXjRRsdHpa/5A6qEYXI+kbO5q2R/r6gUuVedE1qDdkEMHoY2RKoIGVR1S3Y5PS0Nhv571vBlpaXpMqUoh9FboyWAhhoGiEmKlJFxU7Sa9J6wU8etu3diysNVPhobNDDgXSdGWdHsaURXFdi0xh6s+cjh67aCRDgVeNqHtbEQUqTXtvFRqJrU5MTKk4pUPyA9+K0H7BSsxvqWikJNF7J91d60xW+QbuFR72x66PsbffcpMDlZyEca+8BlDTsje94pz6nlEg0tl0vUJ2o8LBTFFqlAsSRq7S4JyjkhRNQsMZEjhQAQfBQpPLzjx49Ii9jiApA8Se/+U0bKQ3aieuCqNgr2IH5BTu4uKj7PTaFT2bHZmZmpWxiksgnKrAaYlyRZtvD9BL0FOPfMSuNVqzdbQgsG9it25lnnrTNtSX59ssfOiZG+lXL+HKiMNCz1lPBhUqyUrGRsTGBK/IwD69uPjPFcEOhZB7Eyz1V9spuTU08IMWFC+fVcDOpkASTlPzhrStlT6j6+wGhBCUTyOgBV+FFK2CkXNYzmE2BfJxVsLw6o8Kfp661OjRxkB1cu45tbGzJpor/7WxV7fjxE/ZDP/yX3UO7AHkzZocOH7fJSey5YncI2xV5i3b3bItAyMqg++K22gIKFDrJELmmAgD2PIS03WJqgRBSrtmura5e1kTH2ZfP2LkzZ22wVNREBc0VuQ8eqojCzuzg4lGphb7wxS+J+PH71CstXDEUFivppZ4EWoKDWbQm2J4TFVkscx9lI0HToDCzVOU6WOeFhxeHPcuVAKhT2cyvkFu97BvVpuG9F4XOPsgmGDDGLlxVRHNHE857Zv/l/uK9LmCx07V77r3X/t7f/wX78y8/ZP/uIx+xFVTfUeR6LSZvnrADdK9Zb0DDXx4Qr3fh9kO+E4hIH1HedYI7/LfGbzWC6yC6vGbDUkOqvO6eQFDOLmwmAN63t7Yc6KmUQy3vGUs0vfmcNUL54jkRRSkHfQSb39IQYD/QkGWNGqM4F97+znfY3/6599vs/CEbGp0QkYOlGU01FmMtvM3bTa294aFB+ze/+qv20d/791YeLPtYNQUtKjop5Fv6Pq4L56DndAQBvM/QBczoly/vYTb3uv9Yy7GHKv028wj8fKahU1GuZ5TGygmLWm1Hz5FP0biS0tcnr6cuTd+rfxOeugIMIOZDFQSoCNnh4Xx+r/N+ZdPNXpkNAIpcb2qwk6ERrdgDb3yj/a2/9dO2cOSwNUNhJTWdJrAAQmjqvHmtYXuH9QH+zM2m/ac//AP76O/+jrVbNattb4ok6nLeULAXzA4dO2z/6AP/wo6ePG3DQ+PWbhc0mcG5hfVTo47abkxKfNUUO4CDZdve2rG15RX75te/av/hd3/LtreuWWmAoHtUqiV78LsetB//8b9mhxYX9XNyxF+ig1ZLGTqcY8ePn9JrN9sOuNFIr64u+3MM9dEIv+au1zj/5Jf+qabgeBalBg3PWs5TAB/PdkAUwHPhEws9YjmsIZOo0HScJt+ijuBeYicT4dZq4HRfnSTh+mpN9VkTShkeE51Jyr6KqND30+B7AG0SXkxUMCdF4yUydJc8Dp+ocN9hry38tX1dOzjp+5wTI77JOpjh5wqf2eMyINsrtnDwoL3lzW/R+TG/SFbFuJWKeEeHfY8AUZTz2LkM2MLCvO1W6wre5dlmPT30xS/bw19/dF/VGGIOJ4DIVnKxgsCwJCLi7WH9pIabWi32ZqkPo4ZLso0PyV5KncY9cJ9Ev3eqq5Rl4jZZLix0ZaeCfnuTqljtcYa5bZWmK1tMKPl+IZFKhsH2hEVOIjpx52SDT8wkARU2cX2eymkDlaGYe7C07FdMOUm0gtc6Fk1MPRVkpUQOwc033qg9TZ7ifC5ZgBVsbW3Nrly6ZGMjQ6pjRocGlakGwJs2ZNQOvE8BRCwaWbEwUTFo166u2Nbmpo2ODSsDza3ZNtVTcH3IpgEUBDQsDY54RsXlDU3OcPsnZ2Ztu9q0l14+Z1eXlqxc6Nob3nCvNVo1GxpyG1lsiQZKTDZ19e+mZw4EodaxysiQMlaK9DbY2FZrNjQ2bn/+6T/TmgZ8hySBkJycnNQax66TGpQvAKcEWvX5mKIQ+IpC3p9H2etqatn3Ep+yArT1HAByb6SqDlsoJhSkmtWktE+gcO4nkeIkUEN7DPsFz1yl0LVBgtGZgqy7FZS1myItWLJTB2a1F6ysr9vcwoL2rMGxcVu6fMlWV1bs+PHjAtmxEZL108i4ra5t2tnzl2xkdMyWVtZtjwnFmDh2QobJwhHtEfMLC33Te/vviwdaE+s5MSZ7G6YTmJr3afZUxXNvhgfLVrSGDRZbVu42bIhJd2qXWtOee/6snb7lNnvksW/ZnXffY+cuXbGqJh13PRelDUFasqXlZXvjG9+os1GglcjMrnoibMywf+KzPv3UM/byy2fdZ79DX+hWRALkE/iEgFDYqdu7SGkd1yC/14n8DGN3LMmnKfJ/XqtR+vF8ObBIv9e0B7/rATt8+JCtLF9Vzgv5IoMjg66YDoEglrDkCVizYWNDFRsrDdjO+qo6v2qtbps7Vdus1q3ZLVm3OGg1bIcqQ3pOsUNtEPorEozAaHpCf86aDQ9tpmfnPbGmhkdQTGPxUtFkCsWC1PKs8+hL2W9m52ft9I2nJVbjA0OAMQXHwZ7XhX5ANXuEE/PfmoZQaDVT5d6Lqu6TuAKLoyH1EFxjnjWyKLa3t/Q9YAr8e2EYTByF80KeIwKltc848UEf6z021rEeyqzJApEtTL36FA/rl7OF/Bb+XJZfUbfxczjrqZ0zEzJJFZ7HnV23jfJy259XroFPsbvVj9Zg2Scl+Lusf3mGEILJXjumkVga9ECe2cF0JnjJoPInJycmNHnP1Ch7Ub1WDeEhP5O6ec+Gy0Xb3Vm2U0cP2RD2SrW6ra+t285mzTZ3dnwSs1S0yxeXjMGGTqtgR46Pav9lnz11ww2cvra0tGmNdtGuXNuw7VrbGntdq3F9i11rIAJotgX46oyXSGJPFuFca9YY79OfvZIdOnI4ilvTBFmSE9w37oVsg4RneG2QhER1d5/MZZ/rn5jJ+iZBdfUKYXeU19dFMTEFGeds1jeZj5GWRAn1ixgAh2GdKtcHq24X+Q7q2cA20Htr9S+hls9CxwkRz7VwZb/XARK7hP1Q2or5lBl1z74tEtMhrNXcZyQQjilfYRIBmIsYwKq9T3ik9yNiIIVwTCj5s8T3sdZwo+B7dN9c6dAD4+UugpA4gHxhaap19kOweR404RtEiAgL8ik0CQRBCq7W1D2WSKxnheXkDb9vEmyPq0ecCcVyyZ771GwPJ2SiQvclwHrJb2OfyBqZa5ukSWZJCPMohzA08Kx9Igms0wUYrIv8EvkZOSmcsUmyu3ib3MH9iRWeSQlzo45OgU+0db39Wtgc2Co9cnxGHQnJSER/oF4qamX1VtH7OhboE1iOzzgxJvv5cDrRun+NqOjdx9f+4zvkCpws+gPKA8+GOS6/74HISdhXmrGp8ZDIt49nNPAu2SBpRLFl7WbDZuembWyU4LyyHTtySKqnDmr4dtu2t7ft4sVLOlgPHVp070eKps1NBVnOz8+pWGdDYzx/t1q1zY2NaFxNoaUUyWMTEyqw2oBQ+FhrisMzHmSforCsQal7AAIyhJBNeHxywlU/YiH9JrKxr66sOsgW1k78lZMQKPS4PvukAe85ixIOKD6HrHhCASXGWhMFDhbwP5EY4YXso58OPgqMC3BKPp+hbMxx7mTF+fO0o+LvKGaY/pDCLVhiB/M8XCoD+fQz+2w9/HxxFQGNkwf87INQvK4Ye0CiUAnh4enqo4LGHSm+AQEEvKlxcvKCAGuCl9sdL/j8NVrW3mMSIWygOm178J3v0muh7pGipeujkyIqADVo1gBbWIf4WqJgklWOh6pzH3M8tsdyY2k1PNQjKrAcIEz7ooiKx2y4PCjrp4mpGU3iHJhbEOCBEm9kkgaga7MH5nQIoKylwALAghjje3wU0a1meJ8qMFpdKwyX0D9aoVmzztqqvfTUt+Qzy+mTahAvFJy553oRRi2/5r5R1CyeAB5o7MnoSNVIvwoSUD+D3Vl7/A/iimKjvrNjzz//nJ4h1qNAnvi5jP57mLordNTIcg8jM4B76mF5rw4bkzqj7N/Pmoeky5/rYLSXclkwcm0obDV5goKfsdsBD7+DqMADHquqrdUtWUT84A/+oB0/cUI2E6XSsB0+ctKmZ+YFBPtD4l6vSVRsMslBUR37DhZOGr9nXarg8JFJt85wZThBcisrS3bx0st25sxZu3z+il26cMFKha7deMN12rNojpz8KuqeT0/P2srqhn3zsccFbBEC1//lRIWD8gn0yY8yCvHeREAAUFozMWGjEVGmlVBoYUeCUkoTCk5U7PHRNQ31atuf/D2gZP5cvY8KHv3hSy81+v6+sg9w+1RV3q9eAYS/K2HS1ao3pKy90TE9ZxSUPIs/8qM/ajfd/jr7tV/7NZE8ORXg+xboMc+3q4oySFs/V016xScn4jr0GoJvmxbJZ4rvS6K0jxnqA+7IuXH1jUjMdsfGRjw0k/NFOULlkjyUAaH5eTmSzGvzbxMshZTkHEvlWrcA0N0VqCjLubp75VKAHpiesJ/7O3/Hvvf73mMjU7NWKo/IEqPd2LV6fUdWIoTscV6gHn72mWftf/qHf9/WN9b3x7xjr+b6CYDqtG18clJkrT53NCf9xXLu13nd8vfZaLEGeb5oah3cTBF/2uk4kJyBzhDHVZpobBqZuEL1rzPBc2wIoXfSe3+vU3OPUq9gYV3mDTN/wL/LfSbPMT/TvEF35a/7+fLO3OuZPWLY3vGOd9iP/8R7bXJuVq+F2t3VxE5uca7kXiMFGK8XuYkf+fBv2X/8/d+xenXbalubVuhgk4LPe8m+/z0/YD/xt37eukUEEgBQgFFtWRHuVLcExIioGB2z0ZExAS/se1ub27Z69ar9/u/9jj381c9bo7VllZKLIE4cPWp//a+/z+697341q71zNAB+aicydLgPx49dZyP49wPglSu2sr4qEg2cut2ERGVf2rOBQsm+8Y1H7UP/8l/os6U6N59Z7WXkd4QCax+8DpUkjW4QFQPs3bEfJdFAHousJpoesJiEheqB7p7ODU189nnlq/7Q2nBrtf7nVXsOZ0haNSkXxcEtTRFAEkMqhP0AqlWylXgutR+HRkwq5hBk5ESF1PipnszmLBS5es0gMwD0AEFfd+ut9sADbxJRATgjKzdNxLHvuyLQ7QSKNj8/r7BcRDfca4QIf/6Fh2TvkhOzgCIJDEBWQlT4+/EMjpwC4xlgKqhfqbf/vl0FyPd6ODWnmpN6Uj9itRnHmh6PIGETtE7Axf2H3YfYc86cqCB4Usp0iAq9Eed1UoHfX0tqraihhmzwaRmunU9GONDgDXHO27piL6cwVJuqqc+mmElhty3EqhFQixrj9Okb7ODsbIiUeE0ma4ox8XvRxoYHBYKM4NEuL3ts3XySMMU1TlTsyVKQMONyZUhEBSKEsfERESN8DypxSAsp1IfI83KiYmAQgdGQVa5u2JVLV63d7tqBA/PWaJm9cvGybHB2q5v23W97syzYtrc3VK+eOHFS5/zAANM4AMD+niiJnDRiwjvCgjsdAfcXLl2SHa2Azs6eepZDhw/r2btw5bItry7LspOJVlTK/YCHsmSiJhMAKQs2zwQUYUiWXwShApZSz6baXIBxg2cVwQrAu0/BeC0MKewTNqk65/sl/NrasGK3o1pnWEEPTIbu2eqVSzoDRsfHtACq9YbNzM8JbGSignyRrY0NO3rkiNt+Vph+b9jI2ITqIiYqmFhYWdu0nd26auSV1VWbnpoycgqoYddWV+3osWN+DoeFhSbzw7YnJ/KyhueaykIEYr83IQLIW7Z6bccGrGHDA20bLJIHV9A05PZ2zS5cvGaHjp+yx598xhaPHrNqo2nX1jY14+Nn15AU/xubm3bX618vsN3fD2pXbGHK1mk50Mt58PgTT9qZl8/Y8DC2gb5XZV2i+1H2EGkn0z30VIRykJU9pW/0dU4w+8TRX0RUcIayBl0hTf/Wsu/6rjdp7SP8Yzq4u9fSRMU2054tRFUzqvQqHCqtXQNeHOSspQcrl215ddWWVtZsZaNqdXrXQsUKJXdBYBmsLC9ZaRDyApGdEyUpqOP1uRd8btn3hrUSNV5liIxJfz4gdZTXwCQ+Ybidjs3OH7BTp67ziVQITuUYQoSQ4zIiko/+0u+5CyIh+bkb7MueLbBrBw7MqAZT1pLqAJ+6AJyjP2PPR6CF+4J6jXhPqr8BSEXWh0I+/OV51hC38FreS0PGYAPmdQzvgWeXHpTPIvIxhIgSf0QundcL2L0wIeP2zxCUvD9NYkCAFQEk/dlu0kNi5yPg1kVbub+yJ/BeqP95DURmesZlu8U0mbsz8MyrX2i7RbHbPiEypO52Bh2Rh3oRH6v2ek42rS0rdls2WGjYwdkpKzKRATHT6LjIZ2TUXj5z1sbGR218DHKlZRvrS5rc5uyu11s2PjFqjWbHlle2bXOrpRDtXYabKP+p+0cgoflZpn1ehCoCysjNk4U25xaCu8i4XDx8WN8rgDiA/MyFop/j37Dnqb+DkKbmjMndtHjKPib7oSSlmu2m10aR19lPUuSznFMxibVIXAMRH3kRbkPEHuH3wycKA/APGyWduajvvcPxcyMEVnpugljOetHJN8/ryrpB1mM8l/G9nnfqBBbXUc+s9nsXBLk40zMKMjuDtce14888FyfyCgJQd7DbiQrVf5G9wJmXLidug94ndg07PvVHfXZHOUGbIiitUe4t91giQUK1XeDAecpZxrOYFoBlbJs7LV20npgy8pnUn8U5SL30zJ/tT1Sc/p5l1VTeb4ekIvbYrNUUTu53InAuMip8GktEC/cqyA7Pp3WcJr+8P0kMgfrRySSRS73v8uvnU+U+teHTGk6q5c/3Z5A939dNTnS4ld7+119EVHiv5PkYSZK4VsexO/Vazk74pDLuFjH18xpR8arL+9pvvhOuwNFORwU1G15aDKTCAaXCiOyOdlVkaAxXzasr4UQKME6nsbOuLFaGhytqWBXeO1CyU4xbF4sKbQOcoFDBu1A2I3jS7TFS7RZQbPaohlC+sEEzruvWHmMqRq4trcobdGV9w3ZQxxFMKl9Lb8gAgAQeAoJz0HGIRog3HRmA/vikh6xWyiWBc2JSZd9Rk7UUDTUgMjYOtfquT1ZofM1BXTYPmm81nV2UAN5MOIPsFig6DArRKIYHs4BoKQuceXWFFb7hPsolkEIWPR6kxPtmYxezHjYROW7mh7RbVuU0Qf+Gps2cQ0IjjD4S56BReNiqMPAulwZf5ERYL2n8Up+ZUKum+wtic6SQcC9KeftSvkLYcMB02lLwT08RMoeSacc2N9ZsZW1Vb5mCDVUkhBKKXogKvihSOORRWdCUcVEAE2QhBUBOMVXHUsUVyPXdmj5HTjdkweEfErsTV8odOXLYJibGfKLi/HmfqKgM9ayfaGTnFg5KQUZhOjzOmnWigntKIcy5LtuK2j5RkU1nKr0grzrUwqgP61XbXbpiLz35LeuQdwAYEyB2FlHpC4+ykEkgb3L8kBNxQwPM5yhXVDz+f+y9eZDs+VXldzOrcqms5VW92t6+9L6o1S11Cy1IQhJiEMYYxsCMJxwzjG0WOYDBRLAY7PEQwzgYexaYMXZIQohFGgYYYxCrgBaLJARob7V6Vb/ut1e92iuzsjIrMyvT8Tn33qzslmD+huiKePHeq6rM/P2+v+9y77nnnEsgLbl5WKdFtjQMNmDzCPBEdtxq2er1695Iew7gnYbDzhpxGa4nBXxxHVloy/fO4pszeNImzEEorpX34lrSR9kD5IGz0gJcznEB7Obn4Fij1k9Y82xsbIptuXlr03YbdXvooVcabHUz1m3FTp+9aIuLpwTy6QsAg0IF1k/9Q2vAmI8CF/OzWa/rHkkEFG/IFcmZHp2wfqKB5uXLz9ulF54UkLGztWu7W9uSy9999+12+tSyklfWY6E4bju7ewJ0rl9fscuXr8jrd7RQkeCde3q6nZGCpwh4XOXkYK+KhwHSq6igwo8XKvjqtTvW2W+5qmqkUEH/l3y/PGeGAGYwrPPn+Wz8eZcM+5EsmAwLKVFUYl8evc5kTqtYsd8Uq40kAXABX3hePzk1Zf/FN36DPfvss/bxP/sz7ZdiDIW8lf4Mnqh788jhWOigIIV2ED3nyehY8b0scnkc5vNVYxrz9aUAJkFjq4OVCwn8wCYnajZZq6mxHHsUezT/R63A+2ShQus3wMtkD4oVLnCfU8t78nBuUNxWA3uYUuzdxYHdffc99i//1U/aiTMXbHIadR2qnq7t7zdUiEVRqCRZlmiH9sEP/rq95z3vVkFYRXmdQXj3elLB91FPsVf7mPhzy4A4FQ3JLM8kY7RIpn1DNoxHNo2+bo7C6mSn8i2Ah536djT9q1hpnHVzlKj3D7GqcnUeZ2E+H9+bimE35EUxxi7ZgaNzNZPHYbKkBRDLOe2ECgUVPb/lv/l79k1/71tVHIMpmskLwAlAvffHcssqxqfT7ulcJF742ff83/br/+9/sg4N4vfrKlRMTJTsu//J99qbv+YbbLwypWbanQPUJACkLWvs7SqpgiVLLwkANs4cQFj2/UvPPGXve9f/ZVeufdGsT/PNntUmKvbWN7/F/vF//212bNZVlQk45lzmWUE0gGRxfG5Rfs7F8bJUerfWVvXZJISAzfLoFtGjYO9+13vsDz78+9bptodnMCPlY2dWqjrYkmrHLAIpOeH8HfNmhVLHsPcRQ2ST9ZDxJwsf0CLVXoAZmoMBfr5ISSeLPycOZLFCcyTUEMNChWyffA5I0VNAhXMYcVdPjHT2aNYl68Ktj7wAJXBa09T3QWf7OeCSY+vnCe/rjT6Z08wLALJjx+bs9a9/vT3w0CvEPCdGEV+NeYs1jhRpnhxSqKA4hcUXIBPWjn/0R39sTz39rH6Pa/FinseP6lPThfEbPShUeskEFMdHT+bz7My/GS/OQxXv1O2US2CEnAXfDyew3M9zT5SiIsY6ixVaQ9HXo3/Ysp7sn15aqPBkNvfw0eeVc0jnYTAdBThTrIjnBSgw+pVrWPoq9jCpPvw+/bWhtBEAQxFuzE6cWLZX3nevx8YF8QD1nDZ3KBpcV9GWIjKKYByu4MsAACAASURBVEBO4kYp+DhDwhv+pYUKgOWVlXUVKiajUIHlxs7OthJyHjPEgkkabQNglaoqXpVWdmxzfctqtWnrHnqvqc889nk1eKXY8dAr73ed8QAblbadOnlahUXWo/ZI9n3FAEPHNgHuxE38nLNcIFBYxDBeqQJg/bX7PVtdu+VF+8GhzR0/LlU361xruVRRg2tIOeqL0OuqP1aSmHh/5jBnGmcw+54shVCPSrGOva6TdEQAAYgtosqCDW++BlDQoaTg92D70jevPG4H+w0rF/vW3ttVzL67vu7WWRFzotSdmpnWOVKqTtjm2pptbW3KHqtcm0QMJ5b+5MysyGJfvPSCTc8cs7XNbamOZ+eOi4QyPz+vNTczA7N7385duKCm58p11LvOBB46e97Ztrl+6EmAip/vuXKMWJgzti9rv1rFrGIdKxe6Bj0IElO9sW/Xb27YqbMX7dnnnlch5bAwbtdW19SDbhvFbQ+gdcbWNjbsoVe/SnGsA5+uOmH/5/yBHEeh4hOf+JRdu3YjCD2QQNxChv3bgePuUC2XLFw1RRYISy8+LzSKzBQWJMpTxWp20M/dB1zxSMGaB8heiQIKAP7NX/VGm5ubsX6fHJH5gCVLl2BJ61Cqf1jnBYqhh1YdGxidMlAXkqDdWL1lDXLkHohoybZ2G1at0XzaFX6o/1oouqOxueL1sOZUbhl5K9+fnT0WLgOcSYeaP7qXIWAWJJiiaS++cPG8DnxyfGdnQ4bpqGDJ+qJ/JLGPznSKAzW3BoNxz1whhmMOEIORF/K8soivuTU9o54qsgyUwsRjA65Vcw2lcvQIUVE8+oswv1wJ7/NLbGwMKYMNzzWgZM9nKvVjkALZC2nOLLuoUFM29vaEcXBt4COQZCi0qOAJBhIe/GkFxwajAoV6jAQAHYoAV0GhkG/rbzAR9hcKBb7/ui0wewXKjr29+lBxqL0+cYqDA7+GDgWoQ+/tZH01Xe/ubdiFMyet0D+09ZVVu/LCKtNJuebZc2dl1cZ1zB2bsMnauB2bm7bxivdzq83O2e7Wju3utmxrp2X1Zteu3NiwA2JqegRYX/Z5nK9cOzkO+Ar7H/frObyfN+xlkCkWlpbcOgxXBRVxGDt6QOAagfrMD0zunz1VeSl7Ico7LMK6rmLwfM+tu1HcuqJ0XH12eH++VEwLUob27SCLJukxCxk6A8UW84KqgOGIS5izHob45/E7eiYH3gxeThoU/uKaXnK46nWZE6b95Sj5RKRRWUK7ElTFvuhhxEwlx2XtOl4Qvb3AiwIvSXVnKry8IOGEJdZDNiP3mM5zDf5onUZ8nj1e2JdkpyxCoxczEvz3dc/ryobtFfNDDbVVdEpLqCPbrsxjlC5m75hgVGk9QKYMFxI/J12Bw9g//qGjZtp3ve3WMLdk/N3JwPP9xMayGb0/I4/nvD8aWKCrLTxmd9FIxmARhDpZI1QaOU5OKnD7LX7f4ydParzh+FHur7gzvjKe4lpVkMFOPgqvGQe/aI4MX3fU81KfojjNFbT5uuxJozM13B7SourlQsWXG9WXv/c3egRedXxeGxngYQYDqs4NBgomYcdIGhZNnnTAStrnMiY2TsB6mPQkKiRT9fqO5J4cTtNIofs9MaoIjCcqKB1orOcMA4oVfMFygFnRaOy5rUKpZBubW7axtmnnzp+TLBvLoltrG0o0CQVhcbC/sskRCHFQ4dHIRoSSgn8LMFQDMmyqymJIcN2wSgDBZaXUctDLmT9FKwOaF4u2Xd91NQWHRGXCmwgderMvEqMsIHiQ5B7ZkgYSLCAvV8DnAQjjyfWwOw5BzJDSOTDnRRApU5CcKeGlEDCuA14+iFiNqAmdB3/ufeeWGF7NDzZyspWjqu4Al7OQtfmyWYux6n6HAiVL4wJq1G83vs8BSBCX7KMMJAj08KNkzI4fnzMCNlmgHBDIFa3VhglTsGoNsONQDa3oHcGmTiHjTV/7dR48cIgQaA4OvcFdKE/y4B1DWhmsTz6TxIf7HC1UiO0UAC92BLBf6WeCvyuKChUqPv0Zq1WiUDE7J+bH4vJJ9ahAuVCd8oD6SwsVLRXEUlHBeKXNl4MpRRuUC1YsDay3t2v169fs6rNPubSbBCIOxVEgWaCBmrTTtNFZ+Xm4Sf2ixlQTKh6yECQVVfDjyU+l5jZUBGoETsw1ACdUSZeeeUbrGLZRFiocvC4abQ2SdZqFivTt1PEXMtQEiYeAsdiTzqRUo+8y6ghnJClgUjdNB5sZH/+98HAtBcgx5sEXzWq5PrzaN29tCLDAGuebv+VbbXYW5kTJzpy9aEvLZ6045sUxFSqkYPIkcA/Zb3XC94z2geaHWHPqOUB3OE88sGyjgfaN69ft5s3rdmvlhu3U12xrc9u2N3etRVG1XLLbL5618xfOCPSgsSrMtt1GUxLmK1eu2ebWtlil/RFBRYKTOVYJXGbCnUWCBAXd2se/2NfExoVRrAaXXcmwBeQFnouiIoY1igoepAwDn2G/mSMvdJ6pM6phpwYwFkFTAv2w85LVzvfEwBnpfUCQqb0w1FOzM8cUqMpKaXZWPSuefvLJIfBPMYX3oxeIVFzFosvoR6yfSKNd/e4FklFA1IMw99bOn+f1CNIcYVjn9/X6YsEOul3b3toUUDQ1NS2rPxhwYmQVCsMeBMwNJUlROOLMGBZCKIbJm9r3zr65Egwmltgpna72ODGEwrLlm7/179sP/vCPyjKkXAWEGrNWa8/a7ab3nqDADOur63Y/v/Zrv2a/8cFfd+ZbsHcA7mDeqTHnxIT8zZO1ORroZhD90nEYLUBq/NS0OUFfB5Q1XuFtnsmYg589azR3lfCyz7CnexDsCW1fPTUc0M7noz0r1jWFHk+S6FvBWetA9WjBk9dlIqgiVFhP5T6T98r/Zxfm7H/4ru+SlQ8KO56nAFHNZUBql9G3WmGfRQLXHQjUWVm5bj/x4z9uT37+c1K2UGQB8/nar3uHffv/+L1WGJ+QogLiI0QDxtsLFZzfEzYzM6v5CoDNZ7b22/aRR3/PfvU//Lzt1tcpzatQsbiwYP/T936PPfzII2J7p71iFpiHILO8f0miJ6Uk4sw+deqsra6tiiWrhIozmv3ksK+96Md+7Mfs6o0rGvtMaBhLVwzSpLY6ZLPx/PKztOeyr4efPTL5ZPmrd0U0OXWQwIsGTrB0azyqc19eUUG/i6LGh68sPuf6+3KKCrFePW1TuY/IUMVaqUe8UCHwNq2cokCf+5lbDB2pT0cLFVl89gIroB4NpMdtZvqYzu53fP3Xyl5mSj12ylIacH9SCavQ1VOhoteFSb8nAgpKyT989I/suUuXtPZF0ggmIfsFqiPvsebFQ+/dkH11BtanZ0kUq3I/y7WiRvZF7+dQ4NDo82q3mOlpfI6+cn2LdRrKWl33SFNkxWyHqahwdinxrCsqKIy4nQmvy9gk9wsBEfTkCUUF69UtTVAfY/gzejVH54vAZIguKjFnIR42s88xsToBkczs2MyU3XHbbXbm9KlI3Lnlgm3v7NjqzRsCJb2RNhZFzGWa5AJSul1qFopeqqhYXdlQ361UVBBvb29v+tpTjFRWjCR1UxFLymkbu75je7sN7SNsBIeDgj3+1FPW7dNTommve91r3bapVrPtrS1bnF+M3jR1FeM9inbVmMAzw6IEprnHPlL16Pohz6DeIncg9qprv2q0AYn92pYW53wPNpjXh1YuYaPjBXFUHVJTeAlfChV8/A9poo1yYa+peKY8xlnupKdu39VmFRUq6PsGkBNkMYGdrv7gs2mIjZ2FCEWA2YigBl2pzibKYyqQXHnueTt1+owA/Ha3YzuNXVs6ueQKoPKEbd9atfpu3U6eOm3t3qHNzC9Yq7FvE7VpW9/csucvXbGZ2TmRxnb3m7JOIrYjv6J46jFgxy5evKBeHmKNi83K/QdLtdtVsRo1PWOsc0WFlmwwHMxTmMCDvkH2Hu+3rLu/Y7NTE9ovUXdcv7luJ06fs6eeetbuf+BB263v23NXrtvE1LTV6WFUGNjC8pJduvyCveYrvsLmF+Z1zvDsiNEpjngPJwpBFfvox/7MNta3BGofwCbH8ifIRGJXo4iETIY0O3qHZGyTOZbHxC+2URHIJYWWExnyPcWUDsIcwDzKvIcfebUtLB2z1v6elbE+U0zhynOKjW61NrBxcifsCftdG+PMAEwrjtnK5paKSJubu2osT8PkIvOJ3JiiQLdnrQOIaIcCk5M1zXpMYD2t2bgmt30ZyAIKZRPkQYpIYAM6EwpuezM5PWm33XZRcTv7EuSy6ekZNcYmlxborl4sLY2rxwr+3g4mc+45tpDqIOWJEUNDHuP3srh8AEkG1QKWTxSUUN1HnEm8lQB1sptZ1xBJIGywpyRbmX2VMw9yJuuP+aszkHxd+11J+RbXoabysi1zADxBdeY476mG6HId6KqQwX2y7/B7zpx3y07yenIWxg/sBUyEe+Za9P/qhN4n9xs+j7FKG2vwBPpHcL+p6JE9VDAJwRIqFDMpYhQH1t3bsjMnF212esqqNFyv16U+29tryRKXe5udnrZup2n7jR2bnJkQroMd3OLSvAqVB+2+HfTG7LBQsYN+0faJkTmTCC4gkhy4GwIFZOJxKSMGBdlAujriUIrx8UrZTp89q/wvlYV8vudMrrwAc2Icckxkl6NY0NU5GT/I1ofCbxQIeY/sAenEA4pwXnRKAgbjn31SMubO+Ir3yyKBSKFh+czc8ibRPo9VuMTuTf1Io8eUHAxK+nxZEEfzZMURoQJgrUs1Fna3IqnF/FZBQVbY3l/S1Wdugcr78pwz3x7NC9RcOQggiiVS3RGOCh43uqrf1QEUv6KR+EjjeQoOLD7hEpED5DhnAUbrHQhKDcFdvUTe6CpcJzmJfBAFG9amTm3ZqXvT+XTEUNQYNutpOeXzgGLWmD0x0qPiFV9LLu4WXCJJBwE3oxg1REc0SLFLNnycmV5oUTErlBSu9HDllZQRoa7TPYXdbapXpIoNwpwsxEbIO9nXRrlOqE/4uSzfFGv7ZwgXiT1McyzeZ0SiMRIVvvifacnpsfhRL6rEg6QkU3+Wo1ju5ULFXzmcL//gb+oILItt5A121EgrEp4EHhIYOkqS3dbIPb4dMABMJ5BiE4HJyvfFBKIpIf7P0eSnWiUhPLSDljd4Sy/mw74HOckEZhMn5qqUx21+fk4HU7dzqCCLZgcKIHV4eHGCz8uDWr01JmHluEe2GOfdnoIAJYH9vnpkcFDLO3JszHa369oEAMth+bMR42UOE0s9FLhmVY6dSZKWVVyHNiasV0p4zDqgCwjEGKm5XjDvYORgDcJ5pKqzucw5GfFsZO7BCDOBBlze54LvO7vVkzr2JLxBAao7h974Or9SMZGb7eicFFAXxQoADgFIMBuCra9NXmx7b0Arz9wSPSIIzhxE4bqkwiiX7TgKirk5u7V2y164fNkWFxckFaUvAGCFQKFGXQGhNx/CigHA/dDe/I6vc4ASJU7YSDH2XBNAYx7usEEAoyV5BRxvt4Z2Sgk85pin9zyKFYony8uLtrHpQPXjn/6sTVUn7MJtt9v0MRonm80vLIlxRYJarjkLcHFhaURRMZC6xxUVLutN4DnHlSDPykU11O41d+z6k0/a5vWrNhi4zzCvyT+pRhCYIimhy3+HQUDYbHDcMBaj48F8IqjiC0CKIG04t3s9W1lZsZs3b1qrgaJpQvOfv5M94IoKwCCXwrsqxsGw/Hxn6Pk1J3jMv1NRwevyPaVW6NDkkMbTDmZ5wcXVUQlUjpej4WfBmXMUKgCtSGh3NralvOE1X/mmN9q99z5gY2NVW1w6bcsnz9nYGHON2NfVHWPjzrTdbe5ZSUCEA1IAcexFgDdcDx70eK+ukWjvbNtunR4WjN++7eyu2s0bq3bj2k15TrMHXTh/2i5cOKueJgqoiiWr4+27u2dXr90Q2+6QhocjhYohaBdM1fQK9eTFA0sFl8zbAMgTfBLwD4MXRZYGqi9FBTYpYrgSeIxRWErWhs+2TNQUsKQsNIoMjEvuQYBQ6oYQIL83u3ZWhgQO+IuHmmO08OY/Q66NEsWLXxQiAB4oVMAI5IsGpwIVA1jrwD7WGnfWiCeQ0ZtFVlOlLylUeOH0SNmRQNrofiVWr8bA5dQ5T30uYKFSEGNrv9myaoVmrRPRr8VVcOytsoSJ3jLJ7sey7qhwQ9M5b+Cs/QQRO4BoxHzMLRJj7dE0Vx1DBTBl/+J//wl729veIdl7Ydx79WBNwV7JfifH0z4MvKZ65Pzyr/xH++hHP6o5yv4OM4r7oMCLmoJCRTK6EqjU3B9RH+S/c+1msYXfI+HNhr6MWfaLyIIRf2difdBt225925uBl7H5o7DE8wIkwIKARMjPOCXRqRhCBUnyFUx/Z1A7u5NzcDRekPVaKFfEAIo1kM89703/Lwzswu0X7Xu+53vsFa94wMaKqNu84M68E5gqTBZ/cE90+VwadG9sbdv73/c++93f/E1Zu3QO9q1chQl4zP7tv/9pm5w5rkLF4WFRbFkK5s19eiChqKjZ1NSMzm1ZOYyNq0/WL3/gZ+3DH/qg9XpNs8GB1SbK9obXvda+93u+26anZ72fTqyfIdAUeylzi4ut1bDdK9vW9o7Nzs3b1s6WzvNKgAgch6hRfvs3f9t+8f3vt/re1lC5kIo24g3O+CIoY8yD9D3O9ZDqHBWuiDPGHTxhrxJYw34UAJjA+/CP9ibrbm/G3M71mgkZ1nKpjMo5lGvGN5G0FSNhdTBf8YR5cYD1o+IgvTE6kE8a7pscZIpc03rG6k/kNiAJ+mdxRNujQAtYsQ7r8nnMt9rEpIo4y6eW7a1vfYviEZ5pFfVnfL57CRdExGCN0KMCkBeg6Xd/7/ftyaee1pbjSTXECbfO2WuiqHTGsxcqOHtC2cIeTY+KiOuyaDgsMIjwH77a2KrBolWVG+C7P7R+yr1O+7oaInp8l3GabODUw4J1iFqrPbTu4j3pE0ToBiifoItY1iOMPjG3w+rOC4uupnCbN/dlPkqW81xwBqkDTxQ7PVZQ8SUKUtx7noFSVSwu2v333+vkI+LR4phtbm3ZzevXbXpyQgQdihVcK2ccYIhsJg7JJYg1ibmFwokQVK5M2PraliwisRzB1pV7pFeUN9HF5pP3pBBZlXKCfaxwddPW1zakXACkbrba9swXL1mTM6p9YF/1lje66lrNkwfqFcN+7s0/S7KeUb87nQUUCWHeO3NX/uqAoVJjA6557iCrjWrFFpdO2BjK5Co5QU+MZyx7AGZousz1YaFCcQNSD/cBPiKglP13fExFtLmZY7a1sSk18XjRY85x+gK03UufIoMrbYiNnJUtgD2sefGthyym3KZYsAr5EUW3fsd6B03RBrALunn9hh2fX1SBB5uUvf2mLSwvakzYE9fWbulsPXvhgnI8Gi7XG02bOTZn6xs7dumFy+rZt7XTsO1Gw44fn7dbq7cEemPty/WgiLn9jtsVy/KcFXMy1iVX+wpIjd4EIlnFvsq0hCRHfgFwDHEAO5oaqoFi11q7m1YrezyytV1Xn4xTF++yT/3lp+zue+61y1dXbHfvwOboY7DftP3ugS2dOGHPX70sFRbFGYFZ2O602+pHRU8hdwsYsz/5kz+1+i72iBXZvjHviYf8XHUyGuA1wG2ufzGRS17UGmXLKl8EzCOuhhxHziqw3lnIHp/42JDJsVYAY++6+w47c3bZyjR/R1kdYKD3buP1aoBoxd6BFQ7pUVGyKZSGe3t2fXXVdiG/qO8CheqBNfb2rVye0J4JsL/dqFujCajv+XQydNkDM950qzEvtjg50fsJCQSlNYYsl+ltEM9yomKzc8fs9jvukP0tr+UXHSDGPpfcAiWf96fwNb2lMUCBQ8zh5Kkj5Tfg8Gjsmz7+ERS4KiMsocjz5XgAeYk+Lx0vhLEnqmCBFSH2piI6HRWHiWvYW2bmZl0hJXKLq2O5RtQbYmT3+4opneGMVZXHwvLdZ67IztCGfS+Y8xDIRICUYgJL0knZTPPejMkRuBtqrSASEmdnz0liRlQnvDfrRcWhIBox9uoNEFayKpzQQyEsmWXT2ju0yYmyderrUlRt3qrbVM374swfX1AujEIONQoKOPaIg1bDylVij77tNnaFzWDHt7q6YxtbXcW+KJcoVPTYyGS766QZEbPCIYDnWStPRB8j4gNE1uPWHRzaxTtuFzYAcK68OBQ6XgyCoe/4SIKxOp+L4964PawyeQ7qh5MNjHHlkGXYkeIx4xs9z2pVzy2LFiocyh3D1aMqBpdRvu37eaDefRNB/PMzlM8nb5X6LgDzjI+4P5RAytdDYa78VFaqHlNnP7FYaH72B1lB6qEorCRZiJ95XuV2wXk/HjNwDnm/E+Xj6b4wYoWWcZ3UCmL2O0Ofe1G/pLBGSsJYWoxrj+p4E3Kdd0FOSBISz+2IqOFF2Ow9wbpwRYIrQym8E78L5+vT24a+F45FKI6WeskVMq468Lj/yUePelTc93c2tW/6szpSfYvwGTmIu754UT+Lglxnjpt6iwyLFhChjtT+ue/JmCHGUaSeJNqFSk5OMCP9LFIxwt/8vtZ02H8NXxufM0oi+c8VKrJfWMaKHhuC06alnStUFPONiDBeLlSMIgkv//tvxQicC+Bc6ZU823zzS/BLqohgPgjsIInBD1M+8d7g11movlnCZOb3SE4VdKlZnCc/Yqoim1UzYA8G+AIsAiRMLzc2MDYrWWZ0vOmPGK/kiCELw6dRvsywKFpNbXJ8LsExoRSHjZL98JOWOqDrVgSwjgTKFr1JOEw7B17wqJzSxioFQ1hbcR0EMynrI6jiS6ywQ/eW5rOzeu+M0DGBe7CcSHKQY6ZsnISEJD7tllQlj2RfSaISEWcXcDircXWxaDvbuyG5de/k7LOhTVWyQmcgZfFCm6Kq+LEZY0cVkrshKBGScfUtiAZISnjF/KAZpNsv0KzQm2hXnKVXIHjvWLVWkbKF31cChr1IWMF4U0hvUEuRggIGGvKv/Jqv9eo6ChMVKmAKOXjHWHoA4PMF//5hoUIM8JReOvPQAdqStTlQdZD2leDgHby59eJCxfmLFCqOGQSeheUTYmJi/1GadDYyhQrmvls/DcSCaTSx5PAgO4GEBA0PewMbUKgombXr2/bMJ/7COvVt3SPFO28G5qCtQH8FQe7Z3wk1TR6IGo9YX+UIYNUkNLwnCU4VyPeQSAMMO1sI4P/SpUsKjqdJ3OPPKLOd3yM5VYI0UjzJgtsRcOuA0yjAKfVNMOQIsrNA5M8IIMmbQfprKHThy+yAC4UK3ZN50gAgCPCPomJrbUMBMEHFhYsX7E1veqtVKlN2bG7Rzp69w0pll+xmoYIpjsqo3ty3YnhEez8aZ2cARNAPYLe+42z1Fgx32KcAUy2xM9c3rtnVK9fs2uUb1m42Vag4d+aEFBUE6c4kLSshX721bteu3bSWGCZjX2L9lNLbUZBPgFewkEeBJ3mQBotC1k+Ac2GXN+j27YDCZjRW1wICvP5rChWE+6NsGv6tApSCWTyEj9jJYvto73TvbcCLVEhlcJsgGwGv/FkJqtm38NsloaxWjAbwzrY7iEKFB0nsCd2e24BloSKTBDFkRgoVjI2KZtx7fCkY5/rDX1vPPIBZvp//Hk1WBaCNuz/vHudMyRurkqCxDtKig6TSE8Eo8gIEpqpMDBjOD1cUqLA0YC470Crvz7CRYX7RuJMml+XxMbvv3gfsp/79T9vs4ikbFMNuo9uyfZRjWpt4gkubpsbxV69dsfe973126YvPOcvI3PYIBQ9qMorjXuhzBnh+vbRQ4XPN1XcvGktZi2Qlzf1rE0TPtal1L/u0rgoVJGsANdik+B6EKrAlQEgswgA8vSDi4Lz3gPEvPk9c8SAOZJLjwIaPn2eYrlahsJV+vZ7AsGe4dJtGjK97/evtu7/7u21p8YSAPa1FVAJqeOr3RoHBCxXYI2J50rc//vCH7T/8/Pvs6gvP6flYAeBvYN/+znfa137dN1ilDFABg/NATPmXFiqYHygqGIubN1fsfe/6SfvMJz+CXtMKg54dn5uyd37Hd9hbv+qruCAVSd2S7IjBxPixzkiImFO1yRmdjQBBnC+AsMRBFCrYs2jgDoHjXe96j/3RH33YDrpNVzrFfeYeK1UczLpYkyldHxYq1P8nvOmjz5T2GYY1VDCyhAwLmX7Xk1klkwOA+/0XJb4eEwA6uIXbsOAYhUKB06M9KsTM90buIrII3Hb7mixUUIB9caHCx417yHNRoHnEnLn+h8QYFRvYWyiKUGDxgirnDKBDZaJsd951p73qoYfs+Nxxm6bJ8Ugyy+1koYJiFef6wUHXfuu3ftsef+LJIyUQxBGYwxS7mw1NueF4DLyJt2yqmK84tQA0jxAN8pnxrNWThbOJkWCd/BWFiixSJEiSf+sZhhe2W5SguMP6yRNuhHGA/FKtBojCa4gFjpiKvk4B3r2ogDWNg66sL821sE4IXGlECYfFW8SOYu07mJkAIkXifE4oq49NTYlFfebUSSmdAVO3sH66fl2NgL1Qgb1oVT9P6ydX94RdK5+H6jkKFRtr27a+sWY0EcWLnXXqhQpYzBRNxxXbU7DCckSx5NUN2QTRP4DvdTQmTWs0vVnswjyFS2986tYah5ob5CLV2pRyCBV3ovjA2AnM4ewMhjxzBEtAKSwo2ISdRbPVFJOdeAiwr9v1hqvM2TZqMBtX0RLyxNTMpPIkCPn04ZuExQxwTsPRVluqCjosp1UKYEqnHyxu2Qa5dkl9gsQUxls8bURh1RNLjuksP8TuZGxghwf7NjVRtu7Bvlbs9vqmzc3Ny/oJwLlziH3TnHIsxmptdU0ALf03JqdmlJ/gnz8zt6DY6IvPXVJ/APp5YTFET4ErV67YqROn5ElOs+N6fVdqeB6a+nNVaRYOmOyKK/YoAB+8+d2u4qKDAAAAIABJREFUh1jFSQY5j0U6wPIEe5VB22Ynxq3Qg2SiyW2buw27cvWmXbj9bnvs80/YK17xSlvfqtvK2pZsklh6pWrV9g/aIsY8/BWvkd2r+ud1espbnREvD1ftQx/+oz8WM5xchxhfxYTwIGeNCrjHJizuhbXkHu1+Rg73LshlI3kc9+vqTI+LIUFQ2PH+PV6oIQ/m/e+/7z67cNspO+zRMLwplSZzkSIexYVDWPvyqGxbddxseqJiveaeihc7zX2Ny87evpQU3l+Rs5s9uqgsbK/VsvZBl0wuelw5+Jd9FHN9uwWMkzvcrspJMTxHigg807TqYh3NLy7YbbdflMqUfRqlMrkLr+G8ESNdPVU8n6JA5NaczpRnXNxyMvrSRUNyfkcFmiiWSNGEdRgAb/RK5Jq9x2Vb700hiGtyHAAHAApSk07SUNN2Pg+yXBJnTAAq8429H6wAYqXGm/UVtri+b3s8w56RasDMwTPeTFtc7esQ/SpeZOA5qsekSJRhtQxbnqa4I8p28n7IfmoSHioLvsfrwBP0OdqXPB4UeQwwHja53BzoMzeueY49WLHXsJOLWDhtqqE2xbidHfpHObDLOqBctjg/a9OTVVs+MWcTUxWpqacWFqy907TNrYatre/ZrU3m14G1aKB9yJ+0u/X9U8UbnnWnZxP0vMTVgjkD9sP92MDOX7yg2Mh7WXo+P1RWBm6ReQ6FA793sATmjeeHsmAKtjl/+7wKomwoVZizrpyFyEfPI3/eXtR3gm3+X+d4z/EIn/P+/tkAWwC8+q55nK0YKdZtjqPbQ4WLRfSwcWWkn8XsSZnvO2Go7HiXMCfXEzl25vshD9IVFYD6rsjh9aOqZR+LkWbQI82YuX/lej3v1cD7OZ7m9klObnLHBqkNIK1Gb6th4TDSC8UNocz1whRrAKtBwHkvuPDmXpT0fJPPlk1uWFal2kP7pWJ5J+4O8x71iSBfHXuR9dM9b18f9udQ/hN9tFznGA3DZbnu5I9U+Us14VGqz5Xo4aKc5ctYQI1wEvUshHlqL/fnrrGL8RriN3HxPCeRBqJBeMaIaRvF+ZKkNF3Hl/kaVVEMfxyKG7cN9NflOaNYMezJlEe83Ez7y47ry9/8GzwCp+Xn6xuLpEWRf4upTtOwVlvBPJuikgFkyDBAopKspJm0Hj9UDqSozlJ1porKYmT7VODQwiOSpNQlTMnu5jOb+y0PWDksS96ISU15YaAQLHW9girVxuSUgDMWJ4f/5OSEPfHE45L4w9ZWxTQDx2A7cm9ihKlq7kCDEh4Ov457Afp9jelzBUoHG0becni91iYcrMOuJYoTur5xrHgcUOD65CFKZVdsJw/IJblLplNYnXBwvIi1GuwM7wtBUShYCgEgYF+RoJq23TE/BPIwUzKF1C085LWZhU9m7NRuARXBn1iXgB3hFQvz1Vlzzgg+NlOz+bkpJRwwHGZQIxweSuqOnB56IKqZLDjJw1FJiPtjSuIeDbUB79Vss9+1N3z11+hAVjNXihORpCngD7mkgPhopp2FCgLNbHyUh7KUHzRgk/rFwS88VZeXmQvrdh1FxWdQVNTswsXbbHL6mBhFyydO2cLSsjxJxyd8019cXNYz4/4A4gA98cAdLVTwDBOIRVGB9VNhfGCtnU37wp99zMa7bbH/vX9BWEdEcYV7kiQeYF0ezc6GSOaBWBPj45rbfAYN82C08zoBPwSEva7mOGoPniWy+Rs3b2g9YWVEIIZyiYJFAl9aZ+HlmIUKFRmDgZHBYILImhfZJwDAPDxeJ6fcP5j5lvO/TeIbgT5zTGyzYFCjsIEVzFTxBna+bmT/tLGpwgJWNBQH3/Tmt9jpUxesWpuxc+fvsmrVZeFZqAAjYr02mAMlL5Kyv8Ag29necXb9PpZwrgxyK4QDAcfNxo6trN609Y0bKlTcuHpD9giV8YKdPLFoF86fsZlj0wqMYI42mvt29eoNu3FzVdJ4t184Cl/yfvl7tBA1CsArcAR4VtPkAAgVwPmeo74E7AME7ySUClKjiPBlChVD8F5WaRnguCVUAn5eDKu8uFCRSabAYQKaBApdZZEBr88FLw4q+ML6bx8Pe5dNY4eXhdaB9hcH/1E5HQ48KSKRSOa+xkgPcHyoqOC/fD9VF1n4U9AZBbIM7BIGzv/nHOV3lVREXx+YZ/R8QMmXNmgqfJbLsh9k/uk8iGdAoSIDfDUrlBTZg/zRHhUR0epsYz8j+e112ipUwHT9+//gv7Xv+f4fMhvzZoyAQYBO7JUUKspqMGy2sbFugFj09viVX/5lzVXGj/XJWq83GzpXxUgfsVwavd/R9ZlzLgNV/T+a/TogGU2FozCWBe/cs1jO3cMDNXfmfKtNTLmiEnk+/tYDT5wTDB/O8VDUJJteYJkSEW+WmSBmFus82PZz332BjiTUud9l/wEiBM6gb/nmb7V/9I/+sUAF9WTg3Kxgf+KMdOacS+NpkDewdrtgG6tr9kvv/zn7vd/6Tet093VvAAR33Xu3/fi/+JdSNwwGJWs228NCBbEE+xSKCv5G6QVQ9dhnP2vvf99P2+XnHrdigZ5Uh3bx/Fn7Z//0R20JxjS9espV7e0J/vr5HcUh1DLyZ67ays1bNgazuzZp1RqN3nd1postdjiwyy9csZ/6yX9nzzzztPX6MEzTS9jBaBWX2SciDlCCFWOZLPm0fhKrTX0q3AJIJSKAdIpT9F7oYgvU8b0IcoiKcABDrUgifc0nMA+bXlZyobzLucBz0O/oWj3JVFodhI5s/k3vDJ6TeiocdMQqPVJUfGmhIpO/YaI6std6Esb+4ISLft8/G+KEQIfymOKyBx94wO6//36bmZxSHCpAoO+xl1iwfWJU4hInIvzO7/yeChXDApvIJd4UFyCdz9OchsAShQr//8AGHKYjVnyjBQb3nvaxUQ8Xxqfv3vwqPyTzLWwGcq1lITv/7zEYYRhxQsv6PbcHVKGO53eIjUNRoA9rjhids3V9bX3YW0ZzhrgrLEFTFZE9NDKBT+/pTLoVx3JOjCgqiNWyWEGhwhV6zJmCwLCF48ftnnvvUgNi1ib9p1BUANqPKioAEdRMm/kRhQqPlbD38Qa9/Nnc2LH1jXXF9oDuzEXiBj7vpYUKivPEga0vouCY1ryuTExZVwrighiwYpCK0VzTZ3MNxO5333OPg/46B7zIx7kNWSptYRJAE9gw9NjO2C2acRYKDsLJqpVcCIu6jjcgL1bsyrXrUlUAVNK0lrUi6x2IUzVX0BITENNg08Y5zPrhjIAIxFp2BbT3hwOgVYNSFVK8MO3qaD+XUTlSwKeiS7pTKhCL7FsJwLtQtGtXr9nS0knZpxEzrW2s2+zxWavA3MbeqtW2q1ev2h133KnPYy5Q6ENVdmt9w26urnmT+P7Art1YUV+4Gzdv2ixEoE5HuRjFcF7PyyFVue2YF9oTREorm5z/AtGCiZvnNDE/hYmxXssmxg/tsNWQlQ378frGtt3a2LETp87aM89eslc++Cp79rkXbLve0t7Z5swmbzPTWfvIa16jPFOFgua+5ib3ihJVbO2Drv3hH35Y+xrrncJZqujTHgjVJP0RHS+KGIxCPuBlNgaOGEr2LjDIAXK9GZZyGM6BZI0niU6gfzga3H3PXXb77Wd1BlFUplAhpRiN1MP6qTxesO7+nlWKfZubmYTKrX4wz1++as2DrrUPD219bVtzu3twaFV6jfC5h33b3N6yNnnvOIUGV/KSuzsbWFGWzttsgOsNft2CKns1qIk44Hq4DjD3Tp0+ZecunNO98fsJsFNEZj5A0EjLWbf1Gdf5wPfZszOv4Drk2NABlKc5sBc02bsXFubV6461LFb3uNssA3qnpQ1jyjNESU0xCFyBvRQiAeuZXJVCt4oV6dFfcPKhx7+A/KWwyKxqvbF3cT/u2HDkZsC+wHWq72b0IaAvI4U9PsMLF96zUzYtASqrCTdqI6zEuh3let5M2tVtGbvxO7JRquC04E3X1ccABwJcBlSoIAalUBrne/Y9ZN9gzmA82Nqy08vz6veyvLigXJdYaLe+Z9euXbdTJ09ZCTLYzqbsumfnUCk3ZLGH6qLdxjaUHpR926q3rdXBBrGkhuzkJMQf4DjEs6nqVcGEo0wKlb6ul1yCeAWVE2c7RQEwGL54xqwPFGRiv6uY6SCxj+1Rb5QkL43GYoy1iItten14jpv5Rdo7jhbzeda8hrFNoqn4VfEctd9H02UH+B2D8kJFNgGHNBqfE6B/xnCcW5kDau2zjikCBKFHNtcitHqRSrl39DLkPOE1aQvOuGTRMIkebkMVRJEEs9WP1ONSL8aEIj/2ceVh7N1ReFR+pHXkuUM28Na6iP6oXIOa3kchjesWGQb8RsQAt88ctaDKjFlFRsZUNrBOUlKvGL23WyP52eB5mgB4qQQKL7J+uu9rNrQn+++44j6LHv7ZODz4OvCY7CiPyRjW7aU80lShYIQMN4w/4x+JbcomPV6neREibz2v6BHBffucYY/xoowDGD4KjjtSWEVd54XvVGbl547+ncUKN/j0/CkLE6O4jUjN0ftmeP0vFyq+3JC+/L2/ySNwWwQb3AOHeYJtKkyEb2hW/90PFsi5rwPfmwy5IkKHLw2PUQ9IATHQAdlhA4ymWkih6U/B4dXtHtikkhqX/hFsuE8mjPyOmpuJ4d+hwdmkqxmigq1+GFa06iQsCbwmq3bp+eeC6RHet/Ip9D4YyCBJBFwpAChCYAMjJX0FvTrL+1fLSNRdnsbmw6HGht1qN21iErDOPdid/erBE9kNB7ArRSreJNpJF/Ib5TPl7RugoRJt+eR55T/9xXXAK6hxVi3MMH5OU770USeQzmY/XqjInhW++ybAfNSIFYDHGxcG3uOZTnwlKM3vUGyRxDUamM7PTdvdd56TrUK90bCV1TVbvXXLxssVgfnyAo6xcDUDTdPaYlY6qx6QFoCdvhuwyiiK9ez1X/N2ByyDGU8iJuknh56aQwOW2TBZg4XEnKHQlYCtN0JzRQXjzfiTZDKu9EJBUbGzvWlXLl+xLzz2mHyJz5+/TVJ3Gi0unThlSydP2NTMMVk/cTAsLy3rme6iqBiYmsg36kimAQP88OGgIcngWhWkU5QoDWx39YY9/YlPyDMW8MTtSo4se/K6KSKoSJEJzrC5Ewm4KzC0xg57duzYrC0tLun73CvBEQkP1kbYmBDUbm5s2MqqN5mqwXyv4gdddZsA9S/BFxKAzBMq3p/1zFcmgh7oudoiq/05L8TgLgHilK02hVoCNqf7nAOkwcbLAzTfOy2lmBOADgwE+4IDY30pKna2NocAFq974P4H7cEHX6UmtOcv3mu1qeNDX3Bnc7ttkQJYgsox2DpdW1tbt/1mwxmF9HVRI+OeAHQKW1gw7O5s2tr6mm1srNqtlVXb2ty0na1t9alZXDxu58+ettnZqWBKj6svyaXnL9vKypqAMTGuRqTFR4COj1uC74xzIFjDZ9XpHUTjUO8lw1hJPSBVxZhAa3pCqJGiWHXRRDr8sEcBsQR/j1avIphIbGDpwe7nGpyFns9FwXU0iSZryH0vWfMAN66McbBDIFuwHQkyVayA5YMlHcwZfj/ktKxN2SVFoYLE1gNuRWlq1phAmMdt7k/toOiXro8M1pWECAgLNkxcUxB6wu6vZ829hq7NEz7OHxQe7pvKWpddGYx0kkwYyQMHgo+uw69X+30Ubvw5+dAKHGUv6x4IyJclDHvF8kn75//iJ+zVj7xWDHQ1n+352hSrjebG/b7tt5q2Xd9S0vr+X/hF+7OPfUxFdO5L7L6OS8Tzc5zlFAXqkCnn3jEsNowUBrV2xeB2NjznaD5vBf9RpPG54EkLQ89ahNXLXuEsymh4GAqp0fNBAGUwRTPw9rPLg3LmrMB7KSf9uSYImmOYrHvFCWKFsYdGa1FY38WCzc3O2jvf+U57+9e83T2xYeyjFAjFh2IKNbXj7O3bQXdgzfqB/f7vfsj+4wd+zjY2rlt/4KxoFG0/9VP/zi5cvNMKBVid2MI1rdna1b6B13athnXMlDV2922sMGaP/v5v26/+0ntte/sm5SkxVt/+1W+27/qO7xRzm7HF6suVS2774gl02DMVvIk7xdHLl6/Y7PF5sZGxZNreXFePLN6D8+NjH/uYvfdn3mu3bt1S8V5+waGo8cQtbPOIs6KRtaZkgEieJHlxweMN7hlAx61g2K+wzlJShD0D1k9Slbr9AMpWVx/5M8xCodQb2MOEUlH3OUzmJNXQfphFeD4oG0trLCQ6+NIeFRSNUVvo/Aj7MJ1HgNTBDFcBZURR5VsInxnBVDAV02oKRjde17zHwvy8vebhR+y2CxcETIl92Hem7uLikpjRrRbWSGb1xp79wR88ao99/vGIJ5w0w5yh8En8iZInG0+zvmg678XXvhVKDiIlUJKAkpJ8inbqpeGqCj84gvGnkX3J7h19figaZjLs1irO+HRFRccGvY7Y2ENiCvERTZ5RH5fKUoOyNxPvUCx1pioM6CQfMV9cHcEfqYWDUTi6X+e+7UGptNAOnqh5NmNUVjxf4JkJzPW9Y6JSFpP6zOmT+n1s7egPNqlmuBX1pgO0Q10LAONWphSzDkW4yfWEYok9e2uLxtibNolqBpvW8YL6SlBsh00MEAjgzLOmUMG/Nz7zVOQIJVtYWLYDAEA16uQaCzY7PaOxoXCRoOdDD79aMSfKAs6NbIrc6bo9Fdee+yZPkdeJlKV+Ot4zhPsVw1vkjoI193btxIlFG5TLtn1jxTY3dxRHTFSdgFLfq1t1gsa4bTs+vyALpZ36ruIyyBaLc8fdgrHVVn4EgA1o06LAc+j2Jd7bzwtgWGowV9y2xK2pdnZ3FPON0yWDMx+Vr1ygDpRPba1v2cL8gixIS5MTdtBqyi++MFayq9evG4p1il86c1Adwk7eB/SftO4B7Gk/L9oHPfvYx/9c/751c8UuXjwvdSr7IDnCnXfdpTMB2xz14JEUAuINvaUmZa+SZIuMo8g1mH9J0qHn4VStahPFntXGQetb6rnG/a+ubbiqsVyzT37yU/bww6+xnUbLLl2+bmfPX7AbKzdlrUhT3bXNDXvNa79C+6UUHICEKEbL9GCQpkHX8wd/+KhVysStruDieXMtzA/ODEBjrJ9QI2Qc48UHChUUiTyPJuZQXjXhtpRYeEl5zucqDnTrE2IW2SBHo3hA79vvuGgPPniP7dV3o5dJ3yqliisiokjZJ6c62Lf9xradXlq0g709NRjf2WtYo92xbt9se7ehM44iE8UYngPKH/JSChbMS8Y94yfmEcW0tExilHPOswdwbhL/MRaycAqlpQgg3QM7f+GinTh1QrEkX1OTk7axgR2bg/jOtD7q0wh2wGexJ7C/cS0o8nNcKSiKxAFJK5T2NGxXsSPIkuTJrFsUtWkDxD5J020+m7yWMWcdk8uxtdFMnM9l8jE36Lsh25mxMZuZnratjS2brE1IVc/MODbrtlAeD6PIwDazEj0UPL4UIYx1gvqhCxbgRQWdFZAeu4fCHdQjMBqiZ6JIrsnnMrcgSjpo7lY5nCk8k3wW2fOO+wX8VQyg/NnjWPaQ6alJ75HQ9jGdqo7b3tZ1m66WrL69ae3mvtV3wRambHF5UT2FZqam7cTyop1cXrCxYt9qE+O2t7fjNsTEMFt1u7W+a9v1ju3Uu1bf61gTdShFIfJ5VCpReAW4Z36r8GRjUg8Fc8kGYwUbFIu2eGJJ55sIrpwFajLuhQnOdFfju/W251b009j3/n4xlxiTBMJ5je/NTlRgrmUOxPPl/djPxTpnrcazSaWqvxfKV8ci2JdEEESJEOSUVAUksUhnI9hHNugOpwjmAc4Zun/y6rAFJ6ZRnw0pr8HR/D7Jj9Ujhb0lLJWYN1lAYa3xNSTcBlHASbcvtgbW70WsP8zFY2/SfekV0Q8olBaJ5bkq2Ps6kBto7MMpQPceCoMkTQjrU/EoLZS8NyfjMbRNwtqdJuHKG8HCvLfaaFGaf6O4cpszxxmIlUabad/79o0gdHlMk/Ey1y5VyhhFIfaCnENBvu47sVJ7VTS+FkEFRCoIXZlj+aniX7JaDaWvfq5cy9UoPJvRPDIJdUNCXBR9VXwh5pbay60GydO9wPDlFRVejPNc2S06Pf4V3yt+piJNEhaFwY1gei8XKjJ9ffnvvy0jcCrsl1i48mplsROwBwANoMLmrv4JaizlTW44XPiSlDfySA5Q+apKKk0ASENJB64FQnfaAowJ0thgObwAHZDxY5EgxhQyW9jQbDj4PU9MiJXH32LWIL+MoIDrwT6DRnS1qUkVCggC2PDYXNUEvFZzX8jNDfmvwg4gKHAvTm9+6YkoyXpRTDVVq5GeRkDLhliueiKb9kguB/PfdV89T+QYO5IY7KQqakIWcsdkU8qzs6d7FxiBmkHWDN4cj/uT/VNU673JnwfRBwSfPffDVAAUBQEl0C9qUOQbqQPQHBguqxRTSb2D3MJACX/I4sRAiQ2YDVWAYI9GfCQMU7a0fMI2NrYE4vOM9ukbombK6U/th4GsU4puCeTN2NikKZS49RNs40fe9hbdex6AXhQLuy+Sv/CRxz6F4FWSVoLEYBiMArC8jsO8deABJeOHR+7S4rySUuxWnvzC45oD589ftCmYdn2zpRMnbfnMaZuYnLKJKffyXlpYVtIKkEGYDSi+V99XgiA5n4pq3iDNAUAADVQ9ZleefNxuPP2M+9OXYZH3pQrK55BFAMBet3EOO5UoEAjADo9bgCsCZO5rfn5R88kDIz+MmNdcCwkOtk9Xr11TcgrDiOtkbWJxoOKUChU+pyQrDRnsKLjCe2aBK61yEhQVgAVbl/eFjUhgA5uCpJM9Y4SxQaA1TGpImrGwqpAYuOeos4VMNkzbmxu2t9dQsk5gSmPL17/uDUqQz992n03N0i+EcXYGb5EEtYBtR3g1dwvW2j+wxm7DrAjA7hEGcxJQDCZVs9mwvd0d29ndsq2tDf1pNhoKBm9cv6agZm5u1i6cO2PTUxW3mimUrNnq2NNPP2dra1vuix6WNwlMjRYqFPKFSoBGjO7/7YAtoHj30MEleVry/NLyJCXnI30QgD4TMKQ+4u/jQH3Oo9GAKr+fwKYKFWqmTeM2B5iSUeNv4kinv6cXYhPI7vUObECBdORzc51pnw4Gl+8NDkSyLnNMePtR66c8H2HfHgGd/t28RwWFL2mYnf8P9a5+n7PCi7kjqhY1TaPvSV2/46y7vpJZgnPmJoUKbB54JsR0uuZDwEr3cuVPznsPTFnTav0d6rgM/tjnKa53ZAFFMD9Vm7S3ftVb7If/5x+2Y/PHJWXnDGg3W7bXwKoBX22YpF3b3F3XGfmJv/xL+/lf+AVbW1nVfsN4sWZkIThiTzVMggTiHjWq9mCY6z7yVdV90LPBFdch46ZhqQMMOWbDf/M77CH7e7a7u6P+Hq6o84QsWVZDhms0gM/mzPlc1Qx0pCkyjF9PYlyNw3t6DMEK8uvIAF/na3oIhwxbhchi0c6dO2M//uP/3JaXlwWG9uSR/+J+Lb4PU3Qa2H59YB/7yF/YL33gvXb5yhN22KPoB0utYN/3/f/Evv6//K/s8HDSWq0xa+w1rdneUTwxOV216kTJatUZa2y1rddu26/96vvtd377V6zbZU65Muvbv/0f2tvf9narVmqhVqJ3BgxuL6CkAlW9s8pV+Ylvrq/Kkowzc7xSE3O6vrU1TDp53a//+v9nv/qr/0l2BJyRvm/6mZlrXgqlMR+7TJSSWaWkSUoKtzVQ8Ud9FHwOiyUeoKWAJeaYEkX/jN5hRz7MSf7IeZafnedzFir8b+KGUBlEwje6R/GZmqORxMmqqNvTPXYpyNGcA6h/RO2j9Rc9NnIvSbvKvG8VX9KKbKRxu5p26swZV3y4vLRkj7zqYTt16pQSY0B6zsiTJ09a58BZra7E6diHPvQH9pnPfHZYCFH/kPExWQeSpON7jt2Tgx2owKrO1AuFhxeEIq4aKVoAVqtQEWoM3XKkvoPC0e/n3pf3LKuAkaRC702xgjdQLzKPf4aEE6k8xtSzijh1afGklcerAvdXbl7T87UCpAonfaRVG7ZPHgt4X5OcR0dWZs7cHoxY0OUZBxDAvC9P1awsi0fspLwnFS/Cn/6uOy/a8WPTIrZcvXLFJifoH1GWL7yYs9gMiYDjPdMy13A2p4mEUFHD3l3ZQ07SgwOAttSX9SnIMTZSFGKI+bFiGh+fEIC8/pmn1GQdEHNqcsbAnr2fEyomEzgohm7/0Jvmttv2qle/WrZAqLSbbVSqfpbImzuOG7439IWOvSsLghBjpDRi3vcB4CFqwZBtCeDDQ//mtRWbrE0rJ5BtkMAfn1cw2m9trNnc/HFbXFqMpvdiCymGc3WIq3ApPGYhz4HyYGtKEeg2Hsx3iFsoprRXYI8qBcOBzc5M28H+nuZIs7FvJ06fscZOXYq/foE1dmgT09N218OPWGtjU8USgPvFxUWdn3ymbHoB7koV2eymNejMsWN2/cplnZHra2vaf+lxcZHGyoBiYkcn09WBP5FoArxReVO5ijN7ibGJGR1cLlll3Ky1u2G1cbOS9axELCu7vlu2sr5lF++425544imrTtSsVJ2yazfX7NTZM/bcc5dsfmlB10mh+v4HXiEgTGf45JT2QCwFUVdiUbq1tW1/8qcfUWFaOWy1JitR9liehXokKKfFzs8BVcXSjAlzIBjgyYjngYkRv9+EeeXxllRRHtdkXwWKbzw7L+gc2p133W6vfvUrrL6zZcUiIHdXdqDEt+xFPF8KFSfmZ62+vW618rjRLWv15oq1uj2rtyh+mLXagOYEB16oVAg6VpCKkEIF+4EKdWGZo2uK/F9Ac7ej6yfW81yZPdRZ6xlzAbryOgoMNE9fWl6UksvJhT7fKVwN8zYxgD3f2drclqpdllcq9BYF9DOz1XAaRX7sRezOpK8OAAAgAElEQVSrxBXMK3Idcn/eQ0qnsIJJj3tenyoH2OpOjnFr4f3WgR2bOSZsgmtSThdgMs+YPVyCzrD+kXWjHB1wc5iMZtkOiguoHnP7MClSsEwcH3NGfwDnqZSQVaYY2SjiPPb2eNgxE9n7hKKAPUz3H2cMa1oqxbBf9bEfqMibjYy5D53TLkZV7lwqem5b7HesWmzbuVNLNomNdadjm+sbUtugkKLgsbXZsMKgY2dPL9ng8MBmZiDoFW1+ackmKdTsH9j6xp7tHxRsp96x7fqBNegbNjA1aCfm9B5FBc0bYm8RSUtVxc3ktDqDIfNVynbu4gUVrh08dza9F/hoQnzUVDtJAR7/ekycALxY6lFwEBCsHiceJ7N3KBcIZWgC2xnTCLuJAq+TTohffF8SHhLN0qU86bn1nvqiikTi+bjjP+wDHu8moOyFMS98jeZgw2bWoUrlmZGfpzJCQHSA2swN7k3kpZG+fsIiQpGYOV6O0VGs6PnSqAOErMwC7BamBXARQQfxkuM3TjTJhtTCXiL2UiEu+jtx5vE8IV5KMSNihRcnU7mSfU+dSufnh8f9qCJc7cqadtKwEyV9zOifCQG3b099eHEYFdFMW71fo4Dna89JoYop5VDhymuuW7lq2DYd5ZWO1wWPTrefvV3zg8AnVWgJtxK/51A0R+FMSuUI/tn33eIe8ojfgxC7yJO9X4e7lXB2gM8Ib43X5PjIQSXIWHoOkTtrToWFbvZxUhElMD7mnkML/jBftn4aCaRf/uffjhE4Fz0N3AbkCAySxyDS4cizxGCn4IANkwBoAkgvVgDuq0oo1oDbEymJVgCNzQ3VYkB7/Fvx2XHZOsAORQXY2i75xLZE+I4WHU2tSEDx/pZlgpjoHpDzewKoCQj0ej/khwmQArqjJp98Dr/DS1UJjaByaM8Tj1OSPoB9VUQd7AVcBzxGUaGqbVgzJENajMDwaVbzKBQgIWHjM1V8gGnRPlCQQ6Bc3627XydMx7AlGe1TQTLJe7C5kTS57N6LIVLFqbG4KzI4lHkPVY1hUcGq5ZciEMqD0i23PCEesmujgZUzFo6klwIjSboIHPFBrdQcBIbpCiAsRm1q4Lzqi7yboJrxgnXCmY+SwpmNMEs4fF5cqEjQM4E0FAPDSjWB+QFM5o4zalrem0HV8ABDBMyrUNH2QsV4Ueyn5aUFAeHPPv2MPf3kE2KHnTt3wVU8/YItnzhpSypUYM3hINvc7HHdH30U+jTrzUKFms560MihOvQkVVdU1oHZYx//iLXWNxTI97E3i8PQgxpnrDIvxICQl60zCrJAwdhzHyQsrBkCX+YVYCuFCt6DIJr34W/GCJbI008/rQKf96aAvehWC7JcEuMZWwVAJk8OslCRwOjwcB5h5uQB6EG091pRw198cDm8SYpJtPCXjKo+r3G5tjO35SM+wf16EK6AJ6ymAEgb9V31kdhr7LuX7HjFHnn1w7LnOn3+LpudPynLFpp5at8ZJ9BhbtDgr2R2CGuiIAunQQGP5q5/DgWt7kGoKXZVqKg3dm13d9ta+95DAEXF85eeE0Me9t9tF87ZZA1mKmzEqjWaB/aFJ562ne2GFypCUaGtcAQsz3/nMySJh4XrAATBgzP4s1ChwlUEnT6uzvzIhs34Jada568rVIwWB/L5cQ0KyEd6VGSxeXhSBbMrwci8HymFpPwA3PK9N4Fk/ibRYx06SOafI7A4pMBHBRyYXaEKyg9VT4z0CI2SaxRRcp69qCgWAHaq6xIITVa5rytPML5coUIJddgPelP5yaFFDXvlQc8LFXxlgSkTl0MKFVHUHX3OXrgg4e5qD8pmd6eWT9i3f8d32Df+199kh9HzAquXtdV1X9fFkuZsY39HLDfOxp95z3vsYx/5qNYma5gknXvJxCaTEhXRY69zENkVCLJtGRYq4jlJTZGeMi5DV+IezDMF0NkbhfnbR1GxJ2WTGtXKU90LMflMcnxzXxJgm4364nxW8U1qEAcYBdhxzgGqxOfJZrDAmvA9exhMZ4HKMxvfn+TwNLC/+3e/Sc21YY/2i9hNHhW7eGYqOGGtaAU7aI7Zk194xn7xF95tn/vsR2VvIivCQt+++qvfYj/wQz9ivd6kdTrlKFRsK0mfmKzYJArJ8rTtbbVtfeWG/eIv/D/2qU/8KRzlYaHiB3/o++z+e+4XU7NUmpAajxgomW4aY8USY1bBb7vVtOtXL0s5evrMOSuMV2x7t27N3V3t0Zxz7N8///M/b48++mic2b7m0pIgk1KdHQANf0UxjyIFACDv65J67/3CuQyhhJ+JABAFf2fBUaRAYUHhGAabnwsqvsf5kPt+JqZHhUbWvrN6c304KOCAy1GhwmMs9js+E59tFG42OGpMmMUKFQt1JgLwu8LmpYWKnDcCEqKXl+IXsTi9MS+gLvHq2dOn7b5775XdU6nsyeb58+fVWEKWnAeoSg7VTPtTn/r0sFAB+M17UqiQmWkUKhyAwK7PyQL6XOyYwvpOyWwoiJQ4DxVp4QUtVxWPB4gVRtdAbpEOdnhym1+5/pzV10WuPCxo+h4Y9pIlWM41W5hftrFCWcXwjY1btrJy3QoqjAD2ep8Y+eUpTiV2RI3hKhHGn7MzvY/FJA/wZ/TM0/2Nj9nEzJQsNIvFihUNtZWvbUCC2y6ekV0a8TbWQcT7xC8TqDxhVaLkgUEub3mfH7JG1XlZUE+W6mRFhQps3bDsLGPXgmp1Z0d7BWsL8HBiqqZiwPiYq5h3Hv+iVcsTApkB8TkH6CdHQWIMQLYNeFZTXMcetdto2EOvfpX2S0gVOs/CThaQRPt8sJQTVJA6VSC7z/HhHssz7B5KpUlvN9UvbKDm3l94/Ck9H+xJmeOQF9hDIDb0B0U76HVsfnHezpw5o3OW/hSltECiDwksdvVF8DmPokLAVqkslZDii/SjoKBAHB77Ml70nYOWes1NTU5oDF/44vP21JNfVP+I17/xjSqAFJjTxYFUKGPVmrNaYf6qf5+D3Kh+vOmrWX2/pViaa4G8hH2Vynj0QNrdtcsvvKDz7o477xxaanLNWJV57uFnV46hrDBkQXwEAGcPgPExt36yTtOmsdTapy8V87dqV6+v2Mrapp277Q779Gc+Z/fcc6/Vmy27sbph84tLtrK6YrWpKc2Tre1Ne+jVr/b+AJF3EStLvVfwNX7t+g375Cc/HU3QXVWVdj2sSQoVqBEK6ikQuW7sW5z9zBNib84nrRd5sLti8DAtYAP4Yw2nJQjrTKBlGfucfTtz9pQ99Kr7rdPeU7FJKg2BYDBzq27TSD+Uyrj1D1o2Xato/NvNtl29uUIzR9vbb1kHe1pANsJ2EGWAcmyw9ptuXSXF69FXNmdVQQUQN843NdjVWVO1VrPlFrUTVRUkE1xmzZw+c1L2T2m7JxeBVM+OkDEoUHmvpLRmc1cDggnW48zMtOYR8xDlp8drR+xxXVfY74BHYBfJuer20RTFvY/i0VlK4Ysm2xAh2T9R9Jcip8WqjWdGj4ZQDUZjXK6JM2Mc8llYOHnI4gC1FxwjjxsvD5vGk4+iIqPXpdT4PV83/JtcEuveVFFmAYc9k7Nc53eQRrOBO/sr40x8Czic1k9ihGN3VCl5w/PID5l3AL6T1ZqD9dgu729YrVK0QQfniKIrPMXuLtrlK1ftjjvvsGqlZBOVcSsOUKU3bK+5K7st8mfUU7du7dphoWrN1sC6/ZK1DwdWKJetSQ+JsDVOVTh4jOy+C+Tx9PsIxSTPrjRu5y6c13h5kSz6GmqsnFAhNduIBZlUKaHG9T4EaVnur/XYx4sdo8qdZO6/2LbZ1XJeHPJnmLiDLM/impLZ7jbNnns7ScXPPNZlxqfKt9I21Q9O7Z2uwvBzVzbVEPbSEih+X64XgVlp7ekavGio/D2q5nxmkgEzN8rrzjmSeJKUhBFbeNHN55XyrbAnSjxIe0v0xcqeTCrigKlpr/TeGMRQHk94T4scW+FSYevkZBov2njMFv1vVXhxVR3rIXEpkWVCUcx7ML4qAo4VX2T99MA7dtwuMnAN9lXhVpDWov8G2JP21ZFcYxijhepDJGW5mwsJ036oNT1i66UCUMypYWEFC+QSa/zITkt53rg3Hdc9a2/w+ePkY1VR/G8HWL1gG3th5lQ8E825PMvjmvS7Olddkci+K5Kh7tcVfIIowh5e8/VlRcXIifbyP/9WjMBxmmoiSxPY7r5uicVJuhjNFwEHZckjwMYXoAIyNXAigJsQ61b2Uaq8+sYlCWiRzXVcySr7rVjv0zNKmvDhx8f5iSeeEOtLR1mwFJBssvRhQlGwWF/fEHOKBFuAGe9JgaNctca+HyAJYCtBD8Aepkd+sbDFcCBpGDY+85/qMOEagp0kZqJ8HA+sNEEjMy+oAMIDXGTgktVVBQw0p+vAiN93uV/2owgpGFJYNiUKFXfeeaetrKwIxAKQ1iEc1VnGiGAXdj9sLrZUMXhIMLGgUMDpwVIGkzAouH8v1rjXoDa2TISDZeXWUb7ZKvEfH7P54/MCnDa3NsM/leCt5Oz5sJlwj2Zsrtqyf8rkmmsjOQLoKhQB3ZApwqpFjtsUaIT6QMqKQc8eedtbg5XgLASuNxmd2EDlwasgH4Y0zdYO6XGC9D18VMMm46XWTxTAkNAuLy+qwPXMk0/ZM089JUD6LIWK6qT1BkeFiurkpJWrzgKdnjqm+Y98VYUKGvDtNt1KCRlkKCrcm5vzh/XAwdi1T3/kw1bcP4A0Zb1g96uBYBRSuE+CbrdJ8Qo4f4sREF8EqSRCqAYc/HYJK0ULZMMEjDwCFBUkDswdrENIvHhvihz5eVjPSN0jhg5g0osLFcnUyCA7iympqEjAVIcnViowhQiGAdq5dvHPCtaNwEGNPSlCBkDK61Gr5GaSwDY/p8Cy19gV+3C/2dZagcx/24WL9uBDr7JzF++1+eUz8Epk2SBriBIJvoPMrMvyWFV2HO19WGgH6h9AoYw10um2Vaho7tVtnz/7e9bYq2tc6yTqzz+vRBpCKcwsFBU0zSWhIlndqe/bY499wfb3XS6vPsXJbkiv+JeoAcTIks91NC5l/yM5KNDQ24MrGJcJ9mu+AxD1DtXbQOB6NMdVwPvXKCpGGToZrGotC9Bmr8jmgEeKDI+gRhUVRyoNFSq63iw6PT/1fqEUUbArINvXZhY6RudQFjdcFeRFT+2pwdp9Kdjq6+dI+jo6D4eMqADYHdx2H1NnXxEMegM+2Npcf7L7hoUKrbdJnS1eqHNv0wO83sMXVSBdFBI9eARocOZcFk+cC+SgmgqtPS+6kQxP1ybtgVc+YN//Az9gF2+/3VV1YzS4b9rWJsXDmoD3zmHL6ru7KiD++cc/bj/7M++1jfV1jU8yE3Msc+/T9eBlGwXEo/FzRUU+A43NgCCXs89jYQXgASoOi0ixzytxUlPerhRnslKpevNFzptM8JKhxDWqsTKJxFA+4M92WACXjy4m4mM2gbVdWDjkc6RQQSElr8VBTU/0pPDRXA+AujCQyulHfuRH7OHXfIV1+s76zj4YWXwDCABf6rbH7frVW/aBX3y3ffzjf2B7jS0l8RSML148Z//Hv/m3VirNW69XtcbevjXb22Itc8/Tx2pWHp+2vZ2WXXrmCXvPu/61XXnhKSsUAKCcr/yDP/h9duftd9jU1DEx7DtK9lyR43uuA+VszLDMaZZ789oVsb5PnTljk1NzVkf1WW8MLR3W19ft3e9+t/3FX/xFsEjdr1yWICPngfbkKD7k88+fC8yPAipgIXMPUC0VFRT8mT/EDgCiOkOjUMH873RpPH9UqMi1kPOKz1EM9ZLeMcazjGJBFigSaJH3chBUXlqoIA7Abip/NwvlDpR7ESzvUc51QfxQnDPiTy2CTMY/kBWsL3CK++TM48+999yr2Gr2uBcpaew7VoSBCsu2ZwedrqyfPvXpz4TYYaBeCMxbeolwDowWKqRsGfezWMln34k6/BmSKuIsz+aULtkHIHRQzIOtLy1UDIswwx3zaG15AdmLFADJqbxyph97x5iYqZPTMzZ/fNGKg3GpD5iOn/vsp619QHNdtF4OkmkA2HIFCMJmHNfrc00d7ccArKHiyaJk3C+/W52ZtJnZeRXuBofx/Dx9thPL83bP3XfqnKYPAtcDuEmDaIBBgClsXlSAkaLZz5MvLVTUbWPllk1h7wVLoexxA6NKoYIQDMsW+pOgqCDn2H3iki3NL9pOvW6zx+YUY8nqE0BZDYUd5EFRDeni2tXr9spXPai5xzmBMpv8Rf0UivQ+wfqirz09gbShfUTYm3mTd1dmV8YgaxGvtjTEFGa2t3bshUtXrdv1nh6A0fwhjyEOZz7Kmmhqwu66607dH2pVwPWizilXOlDcuL6yarfW1u222++wFy5f0Tym39orXvGAwFfiTTUYr1WtQfEARnbHz3VICCdPLNmN69etvl23z3/uCZ2Pb37r29SfCwUOapex6oRtbO/aqRNYeGEHTBN3QECISx2NKfneC1euyrbqxMmTdvXqNTt96qTVpDZo6jWPPfaY8pSLt98WMVFJ1+sMVieRMbayaRmxIU1QKUlmxDQ0lO609myqMmZliB9tYnLvLbi+sWvNTtemjh23+l5T+eBeq2N7+x2bnp0z+kkw9+nFsXprxb7ita/TOqZgBSEpCVIwpVnjWPZ9+jOflfWT4mYcAogJwgucPb/V3lehgjyBG3JbGLd+JE8BwAeYTeBJoDK9S0R4COMVwLtQv5E3SkVOkWyiqnl4+vRJu+/+O63dogcXa9FtpACx6ZvGmUmxhuh8AnkJuV2vZ88/94L1iduqVdtrtsV0V7qu89ftXiCc1fechIN9FfeQ4K5iJCyMieM49+WEADmrqHU7tKgkRw6fffWQhM0/PmbLJ5ZsYXFBsb3OkAB8pSQibsfpAKJVt2v0vCMNZczIlQXOq5+Hq8CYwzRpJ59mvfBz1rLIfzozYO47050cnOvWWczOMhiI8S2AvdWyqekp4QfYQUF8ow/dzLEZj3nkrhDEwACX1YBbykniGQqWR70Y2aHJM/lsKZl07qECcmte5g3qrHQr4HyW8wS9X9qotyY15klMEMErYiv1s1M/UCc8EWcmKz/Vt1JZqfeax3qsIa6F62Qs3J7VLaRRZPJ+NcDfxqo9dP89tr2+LqLYC8/dNNqTlCeK1qh7D9LZ2ZLNzkzYwvEZNdUmn59bWFC+X9+q2+b2vu3U27a53bbtRtvWd+rWi1hVih2pPPzsE5u911exRLGH4s5D6/R7smw8f9tF7QXOOPdigxMxfV8gz9XZUMKCas/7msqW6ahglftEgvOZh/A8M6ZKFbiem+YHdnmOCTGmsoulQTnvTVwatqauxkA16GS7BOvVfDp6YWRB0gtibrmkgkGQhHR+hL1bNlgWWI0NUSjoU/0h++JQYKjvQ8WJwlJPSFnmjdTBrxibzCWzyJL3l7Fcm3kbaR8Xl0UGx1x8LRJ7Mcdkexh2WNwf8w+1OnOVsc2+QQm4u/0me0P0ZgELEFbkLisa2yRYtp1YSeHQ+736fpkFf/Zs4iZfh/6MvPfrmH3+Q7PDyOi+v7M5tMXlfqT0CHK1SFwcunJzcSeB4VwIFRvvz5zQPIrebxrDsPVSA2/2/BjzJLTpAkaqueKchPWr4rdQnWdBKmNC4VpBauBdU7GSz1GxdjibqJAkq88oAAW+4DmUx8AZb7Jesmip/B8cgX1HqvaXm2m/JJR++b9/G0bgXDQSHd30VLCQnZH7iSpQCXae+xB7wkYgyuZOAAr44QCPS/O8mRXsj5JseQisVJFFKRDeoM6g8Ooui/fkqVO2unpLwaUKEXhpNvesVnG2nDc9I6CAMel+jDCp5C8r72Uafbt0ONkZvC8bi2SY3a5sX7yK6RsDQZsfLN5MUeyaAUlGRVZRCiZhm8ncwwsDzmpxmaGq5GGHAqCsPh5ea9brMnEVQxZf/3JZvrr8fHV1JbwlvXLuMmr3TvQE3ntrsAlxsFBc6fcoAJSG7C+vRhMkORDnVXDf8FVZjuprbtrhAOSgUzAU2fT4fMAMAgSCOwIDxkCbdxxsXhTx5n5SU+T+LbcAb7JeqdBgjUQU6SS+0Iw3947aw60MXvWWNw+VBJorqVCRPPCo0g6wK59NPLajMafuLySCOWcJNvCVllZk0FdDPxQVMPdfuPS8Pfv00/IbRVFRq05KDbJ88rSsnyoUB2o4+Rbs2LE5gZ8twO+CWbPdstZeW3OPQgVjSOXc1wXESnpUmB10GvapP/2wTfQG7gMM0zUaYmUCMD09HewGb/dMwpeHaQK7zJ0MOvg3QTLvg+UBknR5EQ8I1A8EMmLFxe/j9UsCxfrKhmuAOWKojXkjd2/IdaTgyENT+Ekchu5z6qDBaFAnGxHAZ6TrzFEOas84nb0dDPzsfaH3KxZtcmo6rGgAWXx/4FmjdFERYb9p7VZHBShsnI7PztnDDz9i97ziETtx+qIVx6oqh6T1E/MK1hOfV6tOW2kMdte+tQ72rH/I2NATByDZCxV7jR1rqZdHU4WKRn3Hbt64YVcuX7a1W/T1MJs9NmMLx+fs1MnjsprBomFjq26Pff4J63ZJeLz5WRYqhmDVS9QVCr4Mr18Kkc6A7xdo0Izaw5NMsVRHGnxhNcUX9yC2D++Qdk9RRH0pwJ+gUp49CmLYA/jMLFREIU1zNOWg2dwh5KLD1w0LqfSBOfD9Ivrm8Hrui4B2tC9FggkJsuWYaM+mCXDsh/qModemF3Cy8Zv2p7j2vKfhHjUM+p0xldeRr5EfdPSuYJ9CTssa5f3Yk7Pp2zQ9KihUwBY3D+Z6A++Bk2vvRYBsgX31CITMYoUz/dlb3b5LSXBzX8VNQNBv+MZvtH/4bd9mfB7nQa83kOc4bFesDKzAudNUsE+S+W/+z39lj3/+87rWLFTwnqzJ3N8EaMQ9spN7wSIYWxGgk0yIudPj3HW2payhggXpQbAzxZIdLwZ9MMF2drYFgMBO5kvnYdhQJaCs5x/9CuS5ncWlkX+r8BB9qUhs8jk6mAscEhZuMWkTrPEzymXYXIefIpAeKvaWt7zFfvhHftS6lEMlC09ViYO+gI0w/LoHJVu9uSnbpkcf/Q1rNjdl/dQfdG1pecH+l//1f7MLFx9UoQLLh8b+porftcmqTc/M2JjVbGttxz77yY/az/zMv7b9vS0x/zmz+KTv/d532sXzF2xudt5m5xZU5GbfSlCEfZfEkRimUpu2tdUb9vxzz9rxuVk7Njtn52+7S2SDzbU1/R7j+cwzz9h73/tee+qpp7TfompxCyhPVLOIw7Mtsv/FWhkWKdIygsRE88v9zisV7Hh4Rib7DPWpSP9qNchthYUH6rau4qxkNHty67L8vA73/fXP9+tCBQjz7qg3T57B+r04Xzwp62qecX6T8AK4OZfXv3L9hZeNbPd0305EHH6m34/HlXylmlcAmJog46s/5j0QkNRbwThr3/zmN9odd10cntXT03M2LiCZudO2D37wtwRI8sX8B/TnOgHYiCeH1k8qvGKq4pZ+kuEfdhWTjCbDKurAOjdXwfrepnBErGEBGTTGHfka3T9lo/mSvkIJvqiKT3Ek4rssVOj5YPkyMaG5WSp4bDkxAVmmZX/58Y/pXPQvj40cQHJmZLEIOBjrLuLBVJCkdU2OfybhPKPK9KTVpmasLDDXYxQvPMCEprH5K/Q9zloKFOnJDvACCMnazWJxFv0EUKGoID6ertnObt3Wb65arVxR7HXQd6uywaFbIjEdJumFMDUlJZF6VHzuGT0DmP6ofrCRRG3K+ENAcO/zcSkqiqUxW721Zm9805ts/6A1bLIrAD1sqQ5RGYRNi2KbgkkpQv8RvgCkmar0H2J/qoxRJHJL0PGig1Vbmzt2+YWr1ul43kBMTV+i+fk5WQ5tbmzJUnZm7pjdeeftAvnp61HsHdqNG9e0ho7Nz3kugH1OqaKGtR//8z/X3IeY8bo3vMEmpqbV02JtbU092hgjCBpcabk0JlXF8bljdv3GTTUc//if/aVVyjV74xvfqLFwQubAWr2+NZotO336tPaDxu6OKxLVc9D7BGDXiX0aYz+/uGhXrlyxEyeWdVxREIEQwt7Gay5cuCibKFQu7Q5qLlSEc24Pc3Cg50YRn+eiXnQ92PFOClKjY6niB1Kqle3QaqWCjfU7trO5JcXr7h6WSmUrVSftkF6BBy2bm1+2J595zm6/8y7ttfML9AqaErHnDW94g9aA7A5DyS5CT2VC+89zX7xkn3/8C2qi7cV1Z+dm3yjmIooKBgyFiYrFxARBbhDoXhpXoUJAFLkn6xp2NNSVUI6Qnzpg53sKZxz9rHjOrJF/cHzR3jF33M402jbb87Po5a+XR+CvGgGOmc1i354d69snCj17tOQNh8tFJ6FMVss2ftiw++64aIedjuKT3e0d29zasY3tHVtZ2bC549PCPGSVVRjYwjyKmT1bWJy18+cvWLcHic+svtezta096w1K1rWCtYgZsQSTdWjfff/DjodCBaq6FkVEyKEoEWh4XCnbwtKSEskkWmqtyHYLlXlLxUQVc7EfC1xFxcEh+91VWYkh8P1UQiQZZjQ3UW4Q/Yn4PX5G3MU5mnsOZ7o7iXhhzWMxj4v9/Z2ExXnn7HYvTrg9kpv4KC4I9Tk/l8onFEmMkRwp2OfKZZ0njiFhK+XFvezxxfeI68BVOIeyr1Nea+ZN3AfXBw7CfWWDeIoZucfILj16hmj8sqdBqAyIp9TbDIJpkFNEAg5saGjxnYSF6A+TFkuyswvRQLnENRx48TJiIZ5H5iZ8fo6nsA/1t3aLarfe9R565DdPPrownPIPfX1d45x7qNxRgjQkTAh8AaxSz8xdQxRDo/KO5+6KwMSuQnk8bL5NoazsCuSwZcpiYyoopQok1wlrJ8bVXVRckennhMfdWbAgZ8x5OarqGZ2bIvsOe9hGAMhyeoQAACAASURBVBzYzFFxyHM5MEK3Rox7pYiN/diYu6+8rKh4+Zz4WzcCZ7Rw3dLD5UNewWUDYUGzKFkQ/BsAQZYCUXnVphLsSN/Q0t/bvUYlmUemCENCG7n79sOqSmkyQAaya5JMkn1dC0FsB7A7ZI1qktMTaI/3s7z1Cu6DKPBEfvkuSZMMTLZU0Zw5iizeL8HZBygC3LMzpGtONA6ZoQN1AnoBnsPnGR98sSVGfalD/u2WQ7DFnBWdSg15Roa8WYBRt2vT0zMCvPx+SHRGJIdsrCTsvAabEhgSITHmgORwa9RJiii+uL2O1C1ZlEi5W5bR02M3NspwtI281SvBYsaTJHTd0y/VGkogAf5QowQQ4g0fQ2bJeIU82N1xvHkjrKtSheZnWFLhB70vRQVsLbVhH/Tsoa96s64hwbPRQkUC3zrYAPNHChXyaA5ZZibQCgSiUOHSxYGACnpUAIg//9wle+6ZZ8TeOXv2vAoV+FQvnTpty6dPW7lGIu32SMdmZhVo0bgKIm+z3VahgjEhQeFLDIoAanrdtnpUHA7a9peP/r5VWTfYPgV45AWCoz+6T3qsAOQEIJqJegZcCQTyvGFkwwDCkxZAlkQd5tv169fs5s0VHdgckAQuHqR4o2w9x1gPavBI8ZBrCkYXDEcCifzKYCZB4WSZDYExCg9U7eHq45sPcMgoEESGDVwy6RPkYm6idEpZbd4XewnPpbXfVAGBQgUA2j4FofGS3XvvffbQI2+087ffY6USPsFZqIDBBRBNQ+O+TU0cw2zXmo09L1TIYow1eqSoQE1BQYQixc7OpgqDG2trAlBozEkiPjc7Y7MzU3bu7LJAEliiK6sb9uSTz1ifSUCKSAYeLHYPLpxFlV/DYoLhF1/TahSwVuxbHxZtJLIk+uktqWIObAua3zWbw0KFW9E5m1578gjTOIHzIVgcAKYHgb5/e4+KF3v6a39IkC0anyUQ7fsZYCDFR9/nxYYeAoTexwbwke9nMTSDvbwWBxOzIbv7b8u+btgrh6Tci2KjYGy+LsHtIVgXe3IWJRPcdts/L8HyRTCuoDZs/rJHBb9PwZXCkfeU8UKu7MPwfI+AN4srrJtB/wgUzjHgM7y44haAWWhCBaO9vli0Bx98yL79O7/TXvngQ7oO7IF4/U69IYsd9bsbDFQk5/o/9Lu/az/3vp9TQuFAdfb9cCbhsEAS/tdcI2Mm4COStGReKSEbYdPDatNYjfQGyf1V6zuAE/Z7LHna7ZZAeSVckYQMk4qRwqaK2eHZ6gfOkZSZ/8pjPvbinI8OxHLBXPfRnMz7iJtxFrFuLYsmA9n1/NN/9mN2+sLtWk/cbyaX/Ga707F2+1CFipvX1uy3Pvgr9oeP/obtbt/yBoiDjs3OTtsP/OAP20MPvdk6XQC+tjX2N9RcujY5YZOTM1Yaq9nayoZ9+EP0jHiPelyIlcWSN7Pveud/ZxfOXtTZQIPe6uS0zgASTOYezxubIVjtgIVXX3jBnn7icTFiT54+Y8snz4qNuL2+pkIzc/CTn/ykfeADHxBw5t7nTYF2qbBLANubXEfvj5gDWRiQTRPFG3n0ut0jYKzPD3y3ezrDWLvlcY+FSOLYf4mtmJd/VaFCTLARRQXXwF7p9gCcX76f5N7ha8gl+ErgYq8Aqf/PFSo0P1jS0VzdbTS9wJoggeZXFCrEbByxJKFZchZTVfTjOgZmFy5csDe+6bVS7HJty0unwiKTPWPffuODv2mf/NRn9Dmoa7AtQuU0ViqqKE8DdKyRZOfHOmQwY08chOqT10KmcasLt+2jUOEWANGTBUVgqEP+ukIF4E7ufbkOE/CQKmKkUOHfjwbglZKVJ2s2O7sgi7Xp2pRVqmP24AP324d+77ft+eeec6a34kTiY7chUGPc6ozOstzXNc4jNnMuwnDiSM47ESim6DcxaUWA+SJqK4/bie+rlTG7/7571ET32rVrVqt4fKIYCrVV98BasPSjMJN/y2Kib2LMVqcmVDTaWFmTIpRiR6/Yk10KhQrAfvYsChWAQNlMe/OxL0rBQrEUCyiuC2BL+94hgNGk7oNCBQW+zc0te83rXhtELO8vJ0WzLKCKRqFieLaPWj76VhWMTgep6cEByFfWPogllIt16OOANZ1bCKEMpSC2axdvu2Dd9oHVd+r6nJnZY3bf/fdYu7kni6bttTVrNuqKA2ioTHGjWK5YqVLTPblly8D2W/RJG7e1tXX1kkDhx7ni7FzIXr6Pcb4TF29urKuXzac++TkpCF73hq9Ukc57mgyswxShsCArtZLtbm9bFWV1WMvKquegY5977DF77eter7xtbX1NzHfZck1WbX1t1a5cuaxYfX5hwebmFmyv2VK/h89//nGpcIltiVc5+7D4uefeewVGEue6/Y2PPWuMfAyrGuv8/+y9d6zl6Xke9pzeb2/T23K2zPbOJZdkKHaKVSJFkJItUVSzolBKYMmOAwSxHQsJjABBYFty8keKBUiWJVEiRXFJc9nEsuTWWW6Zfue2uf3e0/s5wfO833vOmSHFwLBICcpcYDDt3nPOr33f+75PqyMTA+K9NtZX1wQUVBsdlOtNTM3MY2efwb9ZZdCtXNvEsePHpZCY1BpgisDJyUksLCzYNRd724hYqlujcbz66jm88uo5ZNI5W5hoqCTrDrvmCrylbVJQuOv+ENgZRSJqwyPVz8IFrZdVcDL7hvAZCD5pCw3EFAuJZj/Vx3vTOfx8IoeFEJZ+HZV3UHHe/MPNM/CDz8BmpIv/O1rHV1USRJDnHKa8i/FMAvVKReS2Rq2NhQPzqFRrKJYrOHjoAMYLOYHi/BUB1TU1KXioPikWq1KbV2o9bO1U0KUtJ4FT2h+FeoTKf/bQVJGIONZoIUHrJ6qxlRWSQLvfRSafw8z8XMgctTnPIPMsECyV3zJSZ/AZU9bSSHaf1/FWp9tz7CQ87x34794f8P+134XBuhQFIpxaZopmXYEYYWV0UIeEtch6AQva1s85UBJUB14TGeHCLH48g0RqIQ2zrT/k+XEVrVtE8Tg4S/P+S5mxXSMacW7lbHzv2QWy0pY6EAZtvexqbuU5J/xeDfcDKZmfkUQSt5RSvRdyFLzG5ppk7g5m+eZqau9fed48u8JIuF2t33wtXjfuo6oZNOex8GizK7KAa92VofdU3RRmYvx3qiQJWvP/X3xicnCjn3n7rvUpAczw0GxTmFvGLu0KfX7h9koCM8I1s17KMvlkHadMVXfIsBrM6iUjNdjqHoS3oSfV93i2CeeQzMMINu5OJjHihdlecS/wHkxzwGAZydd10p/uFYFEdu1H53pWboQeLQTO+0nh98tKMm69Nz/LTaDi5u7wd+4MEKhwtI8NOBlZZIlySL6/tz8o1D3YSYGiBAh6PQ1ROYjkoEhsWUmsghrA2SIs4IIEjIP6JoetRCuD/x0XOLG0OAgObFB6AHPxMbkkQ6FsUeX3svBjocz3ZHHPHYNWDgUubly00ynUatYIJdImXeUmy8ECh7NaTHs9hclxKO6LrdqsMFRjJ06liHIxgjdfP9oVE88KWhtQscnTYIpsf9pNhGPme7Ah47/zfHJBZSNTKu6boiJHKSSzEMjMbOl8q8nn+7MxKZe0WJuk0+TFDOTkBsAAMVo5aDELXsW+kppU2Rj0GtYEGZwG+M7cCRuolt8gm+PnZRPjg2n+Oxe8Iu15ggyXWDuHKVyQJSkPg0k2EWIEUWWjhtqCAg2MYphbVQM+NkL0eOf3UFGhDTmEM/Fa+ZCc12TAVJS3KsORTVFBRobLI0eBChZFPE9WHNAaIIMFWj/Vqrh4/gKuXLyIfCGHw4ePIZPKqiGeO3AQc4cOyQIgnTFFRS5rVkX0JCXro8YAsEpDm8cgPJ4bXBg8UJJORUWrVcGzX/0SMl3zJu7FzN9VbU4YMJqyh8HkY2qQCKlwA2VTyeP3YSXva2d1c0OlhcHMDIOl+wpjpJ3DxYsXsby8IiYuGb0m92dYndm0OFDB6+IZFcaatrAwAypoz2VfXvT4Bi8pcvCEdS9wsu7YYLqiwvQDFpDFz8/P4MocDRV5bRMM6g02ZWEQw+/Vs1ivSC3ligpaQPFZO3ToMO5+4HW48+4HkcmOCYyQpUiCQ4yYQoAJOBay42r86Zdba5TF5OO9NaqoqFfLkjgXS3sK0t7YuKbGm/YHxf09PccTE2NiMBKoIKjKYc/a+jYuXVpEJMoBcsxC60dAAx/E+hBjcCL7tL8iUKGzB8Q4FRYCagGzVH0FSaqeRxbeHJyUK1IBSAocgAmBQuHPQ2b/9wZTe2HshR+HNqNAhQMK9vxbpTU6fLGhqMnEHaiwonZoU6D7PQzpvh9Q4YNVbwg4FBgAFWrybb0cZUqPNhuDdWd0dzUZw2AYKnAjKHVkxiSZLtntNbGixGgO657sCvs2sMqkGYLMkHQbpllmyFDdw9fwe5eZJz6k5+t7WJ4aFoENQ6BCwaVUVUQi8kH/0Ic+hPd/8IOywyAQSiUJFRVitUatUC6XStq3yK7/F//jv8Dq6qp+XrYBwaPVARtd8+Axq+sVLK90nW/IbJCkmhYzkmObJQLvVz9fg6I2ABW8ljwXfP5K8uQfeq468MR1wlQMfu1CMPuoJYwPV6UEDANzBdLbz9gXvV552w05odddb0mdzW7SsjfYsHY0YP77P/dxvPt9P2HD76Ds8ePnXl+td9BpJLGxvoP/+Lk/w+ee+A/YWDdLlE67jmwhg1/7tU/ijW98D5oten/XUa7tWkZFNoNclkBFDktXlvD7/+538Zd/+WcKk7T9zAZ8H//5n8atr7lNHtb8/pmFAwO7AFrRuCpmcmoa2bEJXDp/Di889zRuu/U07r7nPqSzY7J+inQ7sp7gsf/lX34Nf/AH/173Lc8TwVQNvUfCz+0+oJopGSxIqLZyT3cLi+TgS+F6ASjgoM2eOzYvHQOWlZ0SN/vIEDLIe5IKx78KqNB6FWycpAgkUBEULfSzVkLCyLDAAUrVYlSROqswZFT8IEWF1g6JDkwl5Y2yA96+DjlLTmrfkLOlek3qoYh8sHm/pgmO817sA7fedlIM6skpDicPi5xCCx7uo3/yqT/Dc8+/YAScDJUWXexsbyOdTWnwG6eKV4pGUc2115idVRcEKqwJ53CDIEe4HiRrRMzix23Y+J6c4Ws5C4CgP4++NvPvDv54XTMADSXL4ODIQG6vjYywEUMinUQqn8ekAxVSMfbw2kcfQXl/B3/4+3+A/b1dGw4QpNCHYXNOm7aJQbAlBxfKkwlNv9YQB2aCYpLXRsrNNBUnZJYy/8RsXrW/gCzTPm45eQIL8wtYXV1BOpHS0CqTTGl/ZV1McNSBD2/UBbxSP0RgIp/RNdpZ3xTwRDuvXqwnQL/HDADu07EI8mN59Q0MpCZgsXP2kvLypianTAUgGxcqqTvotXvIM0yaIB2HIr0eypUK7rrnbquZNWQ2hTQHarLvoU97CO5UjgctpAKQzHOhzLCwNvN9lTmhmpv1HG1b6tjfLWJleR1VBQDn9Xyw7j99+hbsb++iTTVgJo10Nomjx48iQi/7bgsbq2vY2ljDHXfcYfYoyRgabVoX9nF1aQXZXAEra9eChahdA4bIM9Saoebyc6dVL9UdwoiZ7ZFBrdVWvsjWygb2dos4fuy4+hHEenZu+Iz0InpmuG9W9nZV0/Pc08qD4dqsVZauLuOuu+/W+25sbgiYpZI1JXVYUTU/1yGqPgjW0BZvdeUazr74ktR3sodRLWR9z1ve8hbZcO7TIpFe92SpZjIaztHGLxmPolevKEw73u9hdXlFz942gR5QzZYXSYX3Ia2gtnZLOHDwENbW1rTGTk9PY7+4L9XjHWfOWA8bBkBmP2b7MAO5L128bDknClTmEC0owaiIIbBM8lXMBlFS3LiiNdh7cLCnPTAMKnmv0EaWx+zDQalrQ96R1V9d/Ho6jw+n8iNV0MC45e/c3OHmAf1ozsCfxRr4nXgdSdYJjQoeuu9u7GysY3KsgKXFVdAeiP1ws91FsVjB4UMziEepgqDtVVwWylMz08jmC9ja2EG90UWx3MT6VgmVZhflRhMVPqOJuDlbtNqav3BOIBCBDHQOU5tNtFvs82Oot1soTE5g4cCCkUOD5Y0Ub6FfFmgQ5kyqF4NVlpFZree02tnDtc3O1OtV/jufa2edcx3ni3ifwLPvazj7BAHYtZqeb84azOLM1YZmV24ZDPaeBALo8MGazQEHY9lzQG8zLX5x7VCoeehP3D3VLJLMtozH44Ns7jF+TLI4C9kRTtBw8ECZRIFE5f2XH5PqCiepjijq7bM5IcKQdCmo1b+b9SX/TX1UCKMeKBE80Dm8r9Td4f25H6heVR9CRVzKFPiaiRlIJHWKMhiZS8uZkJ1/u44GWvgsjeuprLjS6euBirftBJCIRBwDfKzFsN9FsBaYRQCADiimbNB58usRFBieP8H5xSBbLZAPaXNsszhaggfAKfzdlBKcGxroMtrPCxAK5BwRUt1hJuwLXid7j2U1bbCwCgoNrwmtVR/aQKlKdsXRCMmOx8Yj4BzK77mbQMWPZm29+S4/wjNwOAz/jZWWtIU15BK4NzAZzyyA6f3PLzIIuTYwZ4HFrWUXGINEYXMj9gXcbKocMIe4T25UHJQOFBVsFFNpkwwGWZzJzrtoNlrI5/La+PgeZMgSPOGAQCwuheh0cGB+DmP5PC5dvKjvY/icWLcKMmuHsDTza5Z9Ei2iQraG1ABqkhjU1EUmZWwefrG58iEy/fHNconMLnonWgPLTY0Lqlhq9LGk/RFVKG3zB+TGwg2QGzfDtFmMF0ulAHbEVIxzE2Weg6Ry8pll2FtboWqUy/PcsCjn9dmRlF3ceBvkaRM36ZcGigzbC4U+z40af6k6TNWiAUNgARmjx2yxZqanlYPgYbhmrVFHQ6oVKyCcKU42PF9Hm7Sj45LhcYG3hpoKCh4TJecED2jbwwaZ9gD3vOFxfWYHKhyd5j0i8MgDKoOiQt6WAaiQf2fwsfQFX6of5aeYzJrnbH5uVmqOyxcuilXIjAqGm3KQzIZ4buEAZg8cRCrDRjquDYmbNQfTGnRGo6i3mmgwd0KDHg4zgpds2BjZNFMlyuHYxReeRYpZhxzWMMQyMKYkPQybMM/hxOSEshvIHLTrQiDG2Atki1A1wWtPIMEYuAQ3xmVjwPu2uL8t66LLl6+oeOLPsdAig5EbG88FbTAsAIrhasaENQ9HY43w/uDr23BhCKaMAhY+MFVhw+eZrLoRoEJOjmyGeb17PX0Gvp75erJBjZuiIkhspd7R82EgY7tZD9ZPDL5uoFap6VnO5wq4856H8cjr3oRsYVpWIyywGKgYT0dRrpSNNZnJi6lNL0sfvHV6bRW3HDjw2nMAWCmVsF/c07Bmd3cT+7s78s7e3yNQQbuvMWRSSRw9ckBKIF7/za19LF69JqamVAFURIxkRvh5+57fQXa82XdpQWSwPL33VU1YAJZnw6h+pFUCgZvKUFHh1k8MKR8dSPtg8DrQQs970EkNVBV83oP1SJC5+mDRuSH6dEHdYBJgNgssvqzglPIgFJABQR2wg1w664FlssXTMI2DVrNvcYsnG48EwENrjn0Cl+P6NjeqFPBz6pxDATHhNTxIV6BH+DeurRyE+kCVa5ADFQSJFbbKPSkwsgm8chDOQt9VdlzzOJQk9Gby50Cd0UB2IOg2VsuADQkBt95gPPTgQ/i5j/8cbr/jDBChCrGrQXKtVkKrWTVQr9s1JU8kgn/7u7+LJ598UgMl82e1hsVBUHmbBusnvw9GATI9t8HiUCAFx8PBRtGVgn6v+Dqp8+4HhJ4Ghrs72zofg/M+UMAMWWh2Oq4PwvZrNwDrAjCh60+gUioWDjvNAsc6pyFYau/HIY8xvTUoCpaSfEboKf361z+O3/iHv8UbRl7hytvhcZLEQLJBra2Miv3dEr7y5BP47Gf/EFcXX9FxEYzIjWXw8V/4ZbzzXR9Go2EhpZXqrlR/HGzmMsydSOPcSy/hf/83/xKXLjxjwcUhPJ0f8WMf+zAeuP9BpBIZAVDjk5OYm5vTms4mjrWICAm5PMYmp3D50kV8+1vfxBsefwPuuvsexBL0bW9iY21VNjQcVj75xSfxh//hD3X/yY6Awahs9EaaKmfjUj3pwy1TWpL9ZhZNCtMOzY5CBaWOtHtdgL+upYWQsvbhU0OAh/UL92UNJj0jgAN/DdLCfcTrEfYuHx7ItiHYFureCqHadr0Ttp5xvwjDx75CMc36iYQFDnC9h/Y1w5WsfLa8kfPzoPs4KDdNgm/3jFuQ8Vg4HNbnFKhpFlhsJrUHxYA77zqDe++7F6dOvkaZTwzSLpUq+NNPfRovvHhWtzGBCuZZEcjifsphOYfH3KPNysFUuzwWsflCvoLnhWn9CotqcMkJx2kWj4M1Q6WarWwDIMMbVMeRPT8ssOpYS0XMyD2wIgNQE8I94+kkMoU8JsanpaZj/ZrJJHDvPXfhwMI8vvSFL+GrX/0ymo2aai8LNLcMm3jMwBh+sa4dsvsM/PF1kM8q6wZmtElZmmC9bJk+3C95zq0e5v3WxbGjh3D0yFHLz2JuSDolAIk1MK21aNXn6wnPqdcgqjNicaSZH1CpYmtjUwAU63ACFVKUti1MlrUlWcGsveMBDNn77qLyFFjfTE/RMiIiMEJs2n4gaNCbPBrF5s6WaqsHH35QzxRrTO7PvP6sH3z95b3IZ5Sf1wcL7ifNtZu9zGCY0aWdEYOGaT+WVV2zu72Ll156FTNTs7rv+Jm3tzdx6tQJHDl0EBdefUWKBAJkJ0+dxNzMrMgUkV4Pzz39DG4/c7vqcCoBqdoaP3gEuVRGPRH7At6brE94L/JccE3RkI/KUwFb9AY3IgL7EvYBY4UJ9Ptk3LaRSGXQqJalpiDrvxuJ4NrGNm699TWm7KZNXiYr8IZqVu4xBJHEnO30sHDkEBYvX8TRo0eUo8JHoVYpa+dnzS3GcTaHTq2p8/zdl17B+YuXZR3Fml3PaTSG++5/QJZQfC6oOqctIXsjgh969LttpGN9pJmR2Gxgc30dPcSUTVisNDE+NaXnVxZqsTiWr23h1C2WAch17tTJU1hbW8H42LiUFrIaSSS0ZhO0YJ3IdeS7330Zl64sIpcrqM70jBm3AEmmEiiVS2AuNdda9mVu2ajsHLkG0CKS67QNq5RRQEWKhpD0UQ/ZLCQWyTq5if8mO46fvA6k+BEOAW6+1d/pM/DH/RJ+N1ZFvNNEJh7H1Pg4FmZnlT85Reu2pRVZwp08eVLPMAPcm/WqZQlW2shkk5ibn0S5XAOiKZSrNDFLIpLMoEYFBWvDuO2TlqFi9RXXUw3po5ZvSkUcQTzWbrmxAsYnJ4L7hNUoRlIxcEPrrfIhgo0unympkxIix9ncIdTnwRbJB7XsCX34bZaE1nNwH3Og38PQXYXhfYnX4KP1LV9D2S4he8GzK9graCjPzxzmGfy5gUIj9MEEpt2uicdDtQLrCLoh+PfzcwgErRmIz2ORyjaQX9mVWP0e6l8S24IiwT87ibje13GGYIRDU3W4+kAWUswLCSRbz5xhfcjPZQoNy+rgzEX7H3NSaOkbiDTqkXzAL8DZnFdsLzdCngM6fC8pDrhO0m1DpAZT2yt3QeHaBj6xh3Hbd1nopZJ4+QtD66c73rpt5INgqWczLwMSvMcJbcUQkOH7uDMLc3A6di1F5pXdOvt7A4pNCWszJN4zIjuLpGNKBQteD3MQV4QEorf64GD754ob2Z9ybgCzPHbgjkpoPQeas3LWabM72REG1wWTQVrJq14pWIVbbWxKdf0zz33aQD13WbkJVPydXs7//3lwR3tdNRBcUCiJZRFKaSsfDgEHkrBbUUfbp4TsKCzAmUwlDaO0qRji7Kiz+FWB2Up5lS1mNtg26VUYjuhBNna5/Kw1vOMiHAssdoaUGUtNHO4+lRwF7O3vaZPgYIrghza5gNpaADgl/ZYr4FJufV/Pciy8MZa/d/Bm5tCSiywXFMqRpapQSC4XUts8jUHjzaahoWTbGwMuDLKCjIuvy8XNlRrKDGDIrj6rLYJmY0L7IL4+7VcMjbfwcsutMKsZU0tw03Mk2jif3/ulTYIKlyChtNd3f+Lgs8zNUM1qVMfJEFS+t7Na2aSXq2XEdc3Mi71YLKtpWd/Y0L3B62iMBc/CoC+25VCQ4U5ggg0SQ2g5DPNQ2nsff50+9KiiwsEHlhU+aOTno9crCwWFvTbMY1Ksh2BD4020LKNCnACvF62f2FgtLV4Vy5Ug10ECFdmc6NEzswuYXViwIM60DTrYTIvdwLlrCNNu1hksZ5ZYYpOHEHLd950OMskeXnzhG9hZXUWsazZL9KT3UHgNQIN3P38XqDA+hiTtEGQ1xMBoZp6kzOOz0xIr0+SUPQ3iJb0dGxObcXNjHStLSzj36qu6T3JZAyko1WfzzkbIQAv39jarHS9q3MeSxZQPiEetnvhvg4Zc9gdKjgpe+BYiGw0MS97zbQ32GEpt7+myRm7oGvQH0NIHW9xQOajoyT7FLE/oX8rBhDZ6BjCeOI03vO2dKMwcBCIpxLpRJOIRpApJVGo1dJv2zHmRZ/7uZEkyXNIGfxxW0jqBVnH7+7uyuSmVtrG3vS2gYm+X/vzQWsIB6MnjRxBNmH/o9k4FVxe3LJyW1k1i/A7DXkcZ4T540nkTo9nVBPxdUgobToVBrzNalHVDX9d2Z+AdP5pRIfXKCHudx+pghQPBplK4Hqjg+jlg5DRpYWHDxYCc2UAtgBP+fl7ocYjvhbwN08JQLLBJdAzB7k8DRPcLJUNXAz8rvP1n+fuAWK+mwhj/zsDlveWSVi+2dcwuxQ3DS39NP3eDISmbgkZDDVWCAXAEMJmVE4AWD5nXvRiUAcqyCaoWZy1zPeVzaM9IGCaGStCspoYWKH5NVBhrL7E1m+vNxz/xs/ixt7wNmfQ0lk6JTQAAIABJREFUGrU+UtkEKrU9NOpls8SLx1HaL0rF8MzT38Hv/JvfQa9tQJbL1P1ZZZNGsGpQmI/Y4Rh4Y18GRnDdsUBI7gnOsvfz5gNIedobvVbPC5tI2nRwMMfP5vf1KCvN9n9rTPj/fg0cyPT70oMC9bMxZlc5WGp7ptshGstoqLjgesfdg/uQCAPh/3me77zzDH7rH/0WJg8cQD+SUFhtgmHO0T646lBR0W70sL9dxFee/CKe+Is/xuXLL6Je30e3G0VuLIef+bmP430f+PuoVyNiNVdru2i3GshkCsjnLDPi6W9+Df/qf/1tlPbIUA6DXA1zgY9+9MN4+OFHUMhNmCVgvyeLlYmJCV0z7scKsqRHcDYnxeOF8xfwyCOvxYkTFiRLZvnq8lXd9/SF//SnP41PfepPtB9KcRjynryBM4DHFDIEI7gHG0gXHSgZ1aCNrNV+7ew+tp/nvWMNvWV8+PfUazX52ZsNFJt6a/7s3mPQoykoXOXo64w+V1iHnLSgOkO/GChOJY+tL5rHa5jZ0fPZbNc1KLe1MNiihLwXH1r7s09QXJlbpt2QOsm8jnW3ac3wNbXbJJPdsjT8OARWKP+HdoHAI488oswKZVC1+yiVavjMZ/5cgb/MFEinkxqqc9BPIoNCZDMcvhsDUft+ACr0WUPjb3UaFS9D5rMDuL4G+v6gb2GdpGcpNNaysQiWbtetMX0NqnXtBFKEtVbrVgjwlh1aVF7f2UIB+cKEMjikIEtEcPddZ3D69GksX76Gv/jsZ3Dp0nn0erR7DAxGAj7y2TZikZYzWSrYGqJA88E9YfZ0Bv4EEFwscLseCWYEUMmnM97BkSMHZd3GvAQCG1J5MkOE9ghthmkbUOHnlj8ne62I1YSsaWjPtbG2qXtFatFYXwoFDjJIRKGigqQfKTw4ME4lUT13zdSWuYJeR4G79CEvcVBECypj6GvAjz72iiXcc9+9GlSLIdswoEpe0QHs472mIYxn2YU+h/WsADEpvRl2zstLnSnPAWtje57WVtdx9fJV2bKxfi3kMyju7+LYscMKHs/nM1hZXdW90arX9X2yGQNrHuuXWu0Gun0ScaI4ePw4CpPT6LeNTFMplkVo4f3lQa6svVmT25BK0wxEYwTEQ+ZTH1i8vIKVFaoNzFKWjyuH8HML81hZW5Wv/Jkzd4rARPskApEcNHINqzeZbdPG9MwsDh46jMUrF3H81An0GaAcIQBeRUf5S2Hwo+wZs9FFgsBOHPVmG9V6zbLMsnn0QHZqFMX9spTvXKMnJ6nYj6LfaTJhCpXiDiZyWbTqJKFUWR1gc7eIOFXSIcyV+3smm8eV5VWcuuVWXFlclKUwQbticQ+JSAS3336rEefiKbxy7oKUj/fec0b373eefR5XV9YwVhhHt8NnPYJEhNeC9iddpNIJ7DDbScpFKtf4PXb/MvQ+k4yjw7Bvhhczi5EkoVhcAdLM4WGdz32X3+vEsXelcvjHmaHFyaCIuvmHm2fgr+kM/HZ3E/+xU0KtWEWfTPdeRGvRsZOH0W710Aszg/nZaQGbk+MFzWFILKP6lC3D5sYWKtUmdvdqaHViKFYbiCRTaFDlls/qHm9rLkD7RZv5cI1P83u4dtORgX2urN8yWDh4UGuWbMODnaNmRiEDgms4f441Db9Hocshf0B9T1AEcCbBuovzFNaaGrbTHpwWoY2GkZjCsJn7jpNHlXUXgFJZMDEfJhDtuPfzdbi/yLI1EEJGwYFBbgWH/Do2IzPysznBlb/zM3D+MFCjy37X+gzvOfhZuA7zOPmfXF99BqQ6JOSDenaCvYcHuVvdzM/L/Zb7q9tY8fN7nppmJyIFm2LA+3z1Q04lCtZErD2dhOo2VfqsUshzz6dllgVp88tmhap6bF4Y5iUiwhCcDW/gvQj3cFkYqteza0bXEYLXqkuCcublL8wOnoC73rmnfpnX0m3VRVYJAIQcHWTPHtSgUsTZvEtqUYVS2+8+ZyMZzO85Bz0MNLG5pBMLvZ4TaTeo33nMhXw+BLMbmYXniOeGcxt+ya1mJI9Ut21QnPtn4LVkDSI1vO6Dtohe1qcNMzUczNOMlft7aAK9X9Azx9ePLzzs/eFf0/Jx82VunoG/2TNwKvjX2cJuXnMc7PCBY6Adf2cjqMyEJgt6hneahyt7TgEYYajGob8AAMlezfvcHvTAmFSoDX/Whmu+6PPvbrNhzG/2uOzO2DwxV4LFu8nq+EBz46NSwp5UA1FYPPtGYahwWkwVfgax/UKADxcKShS1oQTfeWfbTk5MhqDikhZO5VyIoU8mmLG1xU4Xum7yQB8o8Lxx4G8LDQfzXcnH9b5Ub4Qm0M+XA0BcdAi4qIGF5XrY4IgDGdssuTiL3Sc7EQvA5GdyRfKNd5AzHV2WJnYrm2TaGlHezqaKA8xeB/kMm72MrF143tMZs85iE0jkly0dLXyI9HPj5DVnwcJGUqzOwITlkJN7jlD1MKBlU8xgPTH5lG1B0KaL+97wen3kGxUVYmlxww0qjTivt9gHfzVQ4a9jTKoI+z3dVxwc8jwuX13CpfPnxWQjUJHKZGWNMzt/ADPz8wrZI5OeLSYD9Xg9NECVoqIl9ik9vtU0BoDJB/zM4UjFO3ju6a+gvLWNaMfUC4gySJwbkg1PHUzhvcICjWxNAhVs3lm4sdEnE58NMgEr2gXJuiBsl3w26OnLe39x8QqWrixiaWlJDIdCLq9iikAFvYb5/PDvPvzhZx1lk7jywSWx2ljDZxwNQeZ51YbMzT5YO4gpYbtnAC46Aiq4FvC4fGPVoFwsaFtHfHDOjZjgkXImpBqhzVUbtVJFxaCAj1YbkxOzePt7P4gDJ9hQJpFEQtJ/ARVSY7TFpOUXCwIydskkpFdjZwSoIEuuwnyKPQMqatU97G5vY3VlVTY8PB4FkafTOHbkEKKJjo55a7uMpavbChuNxroalNnk5nrLEy9efC2zYbEDGmZ1ZFkWVjZ4ManCIgwWeM2pWFOhLLWTAZKB1z8AK0aHecPzOcxU8DWAAxwLxeUaZQCvfU6+p62XBlTYQFHWFQFYpV3MgHE0Aqz40NOufSjigt+pBvZRK3r9eebruWInCBnsOGCMWa4jKn5t5DhYvhwE8EG8gMcR+ysHFobn20JcCTqRva31n0HR4TiG2S2matI5ERgzBGC8YLdnwPesIRA9Ckz40JHv7wCRsawpaY/gHe98Kz72sb+HAwdeg1a9j1SeeUhF1KplMW0lG261cPnSJVy5ckmqilqppuP3obDYv2Jok38+BCr8+juQ4dZ7di/QS9XXi+8FKpy1rGEj2Uu8C+QJ28bW1obsR1z55cNef24NuLFi2de90f1m9DzYuYyrfuCaZoW1OKb6kVFQza5hGKJJbh6uTyAw8LWOHjmMT37yk7jrkYfR7kWRiqaQZP4Kw1Vp8VHroFXvYGt9C09+/gk8+cU/x8ryOTSbzN7oIj9ewM9+4hN4z/t+xoCKGlVce7KfpK1cIW/K0C898Rn823/9L9FplYMNVghGjAA/9VM/gdc++himpub1jNIui9eIXucEj3lMHGJSrcGBFNc93t8LCwe1F6yuXsPm5gZiEVqRFUCLO9o+ffnLX9J+z+ErT4+fW7/frK5gsRLV3u/ruJ97vxdHB/S+Fwp4HDD37dzbUN0aIa43vVYHtXotNFmWZeHWlbQ+4lCRx+lfg881AphaneFABesVXmur20TmCMP9YqmIZqumAa4hgSYpYMaR39fOiDOvaxss+H3DwkQN7cB+z8FEoBeyon1N5Of0PydTcQXUzs3N4gMfeB+OHj2uYPdKpYHPfe7zeP7557RnUgWwtb0tECmfL5g1DYEODwj1bB7mbgUVm+V2mPWWB+3qHneXmBEFkl9LWQiaYUJgAPJnrwcqdN4I/GqNMqBCwwGyVUPTOvDX5jVN0SqJodLjSMSpkKCCIY7Tp0/hzjN3oVZq48WzZ/G1r30Ju7tbGlYzb4ePHtUNes61SFs9bzVdyJwI9l+jwKWDN7ZPWB0voCJuhAwCfUePHcaxY0exvr6u4QNrVf1KpsTa5/7v131g/aRa0+zP8tkc6rUG1lc3VAPlGaoa5QC8FrLUEtcBFXzuCFRUXr0G9iACMNLZQX0vb+yIqU9pocrPwDqTz+xDDz0s8EI1d5KKaWMmigzkwxyFuBPUMasGWfoE8gEV3wqpbzRR3i9jfWNdCp0zd96hwf7e7j7WVtalDo8rLyaGer2Eo0cO4eDBWfA2oyuerM/6BuTv79dQKjJ7qaEeQvcxSUPpJOaPHtM9CtajrTbKxbIUqqYepyI1I9Up7xnlLnWtn4rFyKQlQ9ee2ZXla9ja3A2WfDawIwg0f2Ae19av6bzfcdvtmJ2bw9XLi9je3hExjb1gJawbp2+9DaduvRXnX3kJr7nlFLrthoCKTquuzDDLLGGv1bGhvXK7omg2u7Jq4vXO5nKWqxVNoV5rY3l5TXvZ9vaG7LFqtTJarSrmpidxbeUqJrJZgQGlUhmlSg3Fah3xZBY9KsmTKdnV9hHDfrmG8alpLC2tiEAxPTWJ3Z1NJKNR3Hb6Fq3VY5PTeOX8Jdk10pufvdHTz7+AvWLV6j3xTGJo0raLWXbs56J97BKoiMaRTGXQpBKHpDiCWa064Rb023XoblZtxOcpppqfuUqyMY5ELDy33kAul8HvpeewEHrU0b315p9vnoG/rjOw3m/ho+2rmCyMIcq9pNlBKhFDYayAUqkqcs/W1j567S6mJkgETGByIo5cLoljJ46jMD4mdViz2Ue91Uet0cO1zT1Ekkk0OAtJxFV3c32Vcr5lzhJO/OTMiLMf7oDcx1g/zS0smMUbrbBJLgpgBQEJc7/gHCIn4JKDfqqntS4rz8IG46xhmUPHWob7MEENWTSGtduGwO3BEH+UaOhEWtkpMfw5qNH4M3wfVxI4CMG9j3uJ7C3F6g99XZhlce/lWuxflg0ZUy+keY3yWc3ayTJbhwpLAyWCdVVYywVGBAUAZ0rssWXpN8hKDbVdyHjg8Zgi0KymXNnhPZRnd3if79/Hz8HPqNyJUH/r87KXCoHN6nESRp61Y7eaVTMBzRiYS2ozNRGOQ53ovaX6JIJSBJ8GmYLBiSXYIptFlF07/3r5C3ODP9/59h3N1lgLyi0iOGtYrxuCrF2BEMgtds1sbqF+RKCMASMCDGgpOEI+Vs2tYzMCsWUShqJOQx1arhvhxs+Dk7LV0+geTJhNZOj8eQ1TGSPBDsjUIQdD/ZYC1O18ymYwEPiUGxKIMaqtwtxF971fB/678mCtd1UNehOo+OtaNm++zt+WM3BLgp5xNRV5lLYJzZbVjzXcfKi1ULPo1cPJhZ+2RtYMe/q8mhktwIHtxgdHoX8WMMzClwuss98qtap5H8t/nkFzwYoj2BWwuOTDV63UhAILGOhHJCPna/K1W52mAnjrzaYk2ByeS9o8Nq5j8YdZ0r8Y/fAobw/Dn1hUA11H3NmgcEPk93Fw7ws9F0UCJWxoebzyjA5h19qIBixQetaykepYEJDsq7jQWzNon8Fsd7ipck1xgISLPBtqNZGyv7AFXbZA2ogzdm5BVmglDO/MK/rGLwVQk0ElBYqWLUOYbRU1JJp+zgwsbzaRTiYxMTGO+bk5NZD8f3kAa1jKc0xWhQUZkj3IRZcNFItuDwmy4oNItwErxiI3cEKWTzArKFrL8LPcqKjwooI/y4KJQIWKBbLVfgBQ4UNVsY+pBqGPthEtMD83o+Ohly2BCsrQDxw6ouD2fiSG+QOHJHstMDOC2AIVFQQqOCDgLIUFBoGKSlUghQMVrhjg6WQDFkcLTz/1RTSLJcR6ZoERiXLztuEwr7cDATynVHDwc5IlS8sCY/5xOGlZJwRy6DeogYsGBhxY2DCZ4MTq6jK217dkLcasEKkpMlnZPTlQoYImDEpGgQpu7hyuqWgIzGUNGjSQItOEz1yQVno4Gf8/ZXZG3SDppLRdoV70gu/bcN+AMwvdHAyNZJ1kQIkBfCzazHIkQil8yHGplcoaNlP9YMyMON7/4Y/i9vsfRSSSRqLP4E+GhiZQrpMN7LJWU21R/cSCivcarQL4iwNA5lNUK+UBUFGt7GJna0uhqbRlILOY58oUFUcRjbcEYm5tV7C8RKCC15JKHQ75h4oKH7iOFpo28DFFhQNMpt009ox/74BxI2DS2LpsWHVfBaBCz14ouG4c7qrwC0W4Dyn1aAcZMIEKC3wjK8dY2TYbNJm0JdSHQTwZIP6zLN5G8mFGP68zbsRO8SI0hJqpYEwOswxoC2gDXfqQkklv97IDFa6q4D2n8zoCVJjdVLj/ApgzOoj1Y/fn3lkvRdrvNMhoSogta5wss92TlUtQFPF3P0a/V73gdLbwQFExsrD6+3ohOBgih4JR17TfxelbT+GXf+VXcffdj6HdjCBTYNNQRb1WRoNrfrA5ohpq8cpl/N7v/R52N7b1Tj5EdsBCRABVr8NcktH3FSN0wHg2SfhfpagYBSpsHyH7xwAWZre0GvURRroF030/oGL0PvNz4tfW34M1g7IWBNiZuog3nl9nXgOtcyq6uV5yWDt6FxgLinsO1U6/8AufwNvf/360ehGkoukhUAGgXOmAirfFS1fwxSc+i6e+9VVsbiyizXPeaCM/UcDHf/GX8K4f/yiqZXrcN6So4PFmCVTIAqWLT//R7+P/+T//NaJ97lX2XLo9zoc+9H489tjrMTtzUM8VgWs20LxO09Mz2ivVfDFYMaxxU5PTGk5trG9gfX1T35NOUjqfwrVrm/j93/8DPPfcswq0brfpwW7Xzs+lP3s6x7GIgApnBWo9GGWJBbKFrxN+HzlLzFQU9uw7GCVglHZ7ASC10sAaJjVfHKimkgNWoqqIAaAZ9iZ+rz53uFeiCa1Zgh69CR/NqODwcgBUhEZ2BKjwoYHud9qQMtMpsA6thjHA1Y9hANx2zeLQ781RwI0DXn5E7gGPvvYRPP74m5DPj6PZ6ODzT3wBL5x9AakUgQvuH6x7SNooCChBwupbyx8zlp+v3X49fADgS4VaW2EK3tzaWm3PLasgszlT7pGDAsxlGHgVB8UJjZVGFBVWRw/BVYE6QcVMRUUml7Ng+ERG5y2ZjOHI0cN45OGH0G72sbezhyuXL+Pq1cu4dOkiquV9hSsTVpJDoWy8PN/E7A/1RI4AFX5++bszQ+2+IjmD78l8JwMqjp84iqNHjyqDhzU262cyKL1m4P7vwNR1QEUYZNAerVFvYm3lGmKRqICHfrQvey4SlEiW4sDdFRUMq+f9WnplVaQSqSeoEg/7idiNfWaQcRjdNnVEJIL9UhHHT5yUgnx2bkZ149bWJhbm51Wj6JhZ37Pup3Ura+coaxmuYS3ZIVFdRRvJdrODzY1NvHruVYyP5/Hggw+gWC5je2NLKoFkPCV7IRLv+evkyaOYmMghmYgiU8ihQ6CEGRexBC6+fFHr09raurIVSPZpturIjeVFrmE9xv4sSYVIrYHCzCwalarZF4pQFhQrXdpgZVRz5QppbG9eM1V8IoXizj52dopoNNrKnZiansLe/j5m52dklcnMjjtuv0N2dZvrVFD39P+saVm/cj249Y47cOLECd1bx44eRqfVQDqVQKNaQmlvR5lXKdoqJujpzl7P1jkq7kh+Yd/JYyFx6MLFJZRKDTRbHOSx92HYNYvoDu6++wxajRrq5X3kCKBGo1pv90sVlGtNVJtt8B7guaAqvlJvYGNnH0ePn8D+flFEq8nxMdnZdFt1nDh+TPfkgUNH0Y3Gscvas1SUNdO3vv0MKlJuG9mNPSfJXAxJZ4/G3qrC3Cla8sUTAipIfmLIO4GaTCKKXquGx1/3qMCrYrmk46s1Glg4dAjjhTHdV6ydqfx9YL+On1wtDsgs1/dzQ5LL9f9+8283z8B/+hn4Z/WreCoL5DM5LMzMIJtKq//dWN/Czt4eZmdm1BvVKwQsaAPEe72NfI7PL21MO1IbkiASjWcRSWTQpzsG5xaxKOrtjp4Hkhqnp6b0AdmXsU7grMFzA7j+MjeUIKgU98FGU0x9zj3Cft5qNNQvc0bD12Emaqdn1q6cCXHfNJA2EDPUKw9rlQHpSgrIMAwO9pp8TSkIff8Lltlum83X5c8TIOH3WuaRDYi9v+XxqY8OM6BhDWzZC9z3RaKldfrYmP6Nf2a/zpmaW3n693F2xTpEyudgeTvcHy3YWXZJbg0lOyLrv0frP85nOFxnzhu/17PQeM6cvOtgzKB2Gah4h7ZHbo+lDB6pzoOqjha/st81+1PfJzXQDzkKApKcgKOezlQMJHaw7+Z8jyATr7mfc+9hdT15D0QiePnzQ0XFHW/bHtQNdn5MBWrguynx9W+yyQx5IuylWYcKICIrwNTdPDbP8pO1sI7C6ky1yK4yCSYp3vtxC1OHoFmgzWyU6yVQyZXnBmgZMGGuNOZMYk4vprKwGZ3Nd0yJofcIAe48ryIahAw3ZbvU7F73ay01ELNCZAFpNaGO4iZQ8Z++ON78ib/dZ+BoQHXJeOFgWF7Z2mDa5jsf5WZQU7FH+woDHGn9ZA8ehxryspM1kQVq8+ddxkTWvlRK/Z4WZ4V0crPgRDmwxKz3VmKCHjxmAziayGbAUHUOH42lw4Wcw3UG4pIFxeEUAQL+mT+njYUsFvrqBz899z32IR8/IxdTIfSdrgaXLHLNq9dQ28FATKxzyynQwDY0QDYMNOSUmzqHxiy+xWbUYIANTcdkXeF9hsBBUJUMLB3McoLMA7L8jX3dxTSDtr1Rardx5coVFdlkAHCoeuOXSNNhsMANxq24BCYofJLBgTFTUHA4zXDvLBtcszYiEERwhZ+djRmLAsnxdWy2uTPwjsfL4TPPm2azhDU46AzqGQ5gbEnnpkGmOxUwNgSiosIHYZLthYAj5aMQqBBCbEAFfTR5fbhxacBCpkZoQv368NoqXEmsUQPICFTwvr22soorly5KonfgyFGklFERwcKBQ5icmRVTRDmwwfrJhgwRAypoT1T+/kCFsQlaiHRr+ObXn0C01dFA3RUVUuuEEG4P0maBw4ZXG2r4f206/YgaI9lZ0SIrZmxasi05CGBjyWMmUHH+3Cto1lu6PlmGMKYY8mpARSpFxYvlRRhjYMgu9SEnBwd+z/qgxQe5KpBGbKK0idLagTZLyoNhKLBJKblJ87ln4CTvD99U+ZpmMUN/Xhuq2fDIiik20by+PV7XroWk0/pp/dq6wkx5b9eqTfzYu96Lx97yLkQjHE7SezuBZD6JarOBWrVu4E4ITCuXaH9gAEWrWbOMinpNXsks0rhOlMv7qNeKss4qMYCx0xnYu7HxPX7sMJKZiFhzG5slWT/RzoRAhW4Qk8gMmBQ+qB0t9Lh+CdywUxSKKhZM9l0DxgMLMT2PxjBmQ8t7n6W0W7p4JoY/y6M/r8JQw6WhTZIXLyIeh+E2h4geuqYwY7eiUlFj6gjal9nazcG4DRlV9Iz4uWot4jMaGCN+D/jwjEAFv+QNPj2NSqWiX1Zk2fFr+B3Y18ZGtoyh0YwNK/qCBQ2Hd2FQacPWIevcz4WvdVTHMJBc1iIhKFWgYIaAs1nhOFjIQc3okMyHj8Y4HzLIB2voCDN6dK31BsIuLH91kM2n8Iu/+Ct4y1veh143gfwYnzVK3mtary3bpy/rtuefexafe+IJLF64NABnCKqM7i8WIGRKAx/UqogPRfQQhOSw0Cz6NCMeXP/hJ+a1EJMqyMidqU0bEoJ6o0NXvwZ+T40CNDfeh6Pfw9pBg/KQl2HycS1vgy8vtO380Vud68PQwszXdP5Om8kP/cRP4CM//3FZhuSSBSQ4CI70wDFiqdRGo9bAc08/jS8/+XlcufgytrdWUa3sy4IgP57HL/7qr+GNb3oPalWCDGb91KUqM1PA+NikBmL/1//xO3jiz/89HXLDxeRJtEbnve97Nx5//I2Ynztoth3tlhoGAnG0RKCvejZnADeHbqaSS4v0wAyvvb2iQinJ1eB6uHhlCX/0R3+M8+fPodWiz3zLcjdGAtJ9uC0QTSGVpm5wezBvanxNF7AZ2FZ+PXT/DqzhDKjwa8xgy3qlpqaVzxxfhzWZZ1IQqHDrJ3+9we/h+RThJGqsc3+ubXenIYtd8G7LbNGoeDPrJ2emmSpPigoRA6zB069wr8iuLWlqRLP+NAaCrXumVhMI2zUAY1ALBGBca0akJzsb3t+8Rm972ztx+vTtaNTb+NKTX8F3v3sWmWwam5trxuTPjSHD7COqjKNmpUDSyWgzrkDIkN3hz+R1a7v6xeuF996MctjuQIUA22DXJuaemt+gRiHUGvyeBxYaYXjjaxfPmwLOE3FTVGTHNJTm66bTCQ3e3/iG14PlBI+33bDcq2efeRrPP/9tVKslVq3hfrdawwBKs/GS8ipci++3DlhjbHsiB7qpZMYUUpEeTp46gUOHDgqoUGZWhmBFatDYe0jqsJFXwYpIlIqKpAY5rWZbSgSebxF14kClUlbNoDo/WD/xddOZrJ4RKips3UhoqKU9mmrUbAadpllGsK8p12qqQUrlCk7fequuJ59rginsPzJah0ngYH5AA6Vq1SymCFTWGvqsVIr4Z+P9XS1VZRW0srKMerOGbDaF+fl5kXs6rS4qpQomJ8a1TywtXsSx44cxPp6TzUoqTeVmVEBqfmIKK1dWUau1ZbXKYROtn3i87V4HC4cPYXpuHq9892UN9POFMSwtLgfrTeDa+rqAGgPCqF5gL9TH4SMHZDfFmph7/NUrK7h6dVXAHXsUMqt5XQpjealQ+d6vffRRPVvLV5f1LLBGJfLHvoBkq7vvuQ8HjhzGhVdexS2nTqDDQX0ygXq1iN2tDeWKMYuskM8qnJvrLtcDrjmqEcn6bVOpksJLr1zC+saulG68Lspsk1VcBw88eB9qlRI6jRoKVJjEo9i4toFILIHNnX1MzMzL9555JBPjY9gS9rmxAAAgAElEQVTc3sVeuYbp2Tlsb+/qtcZoTVMuyZ7qgfvvxYEDB8nA0f60tbNndlO9Lv7y699El0pu+r92+ew0FAjP9Vv7YjKOaq1ioy31xiTxsYfpIM3eo11HpNvCJ37uY6hWywJByDKfmplFNp+zgFn20k1mtTXwrhev4O6y9ZA3v26egR/mGfhiaxf/pLqIRq2NTCyKNFVF4+PIZvOoN1o4euQIpqfGkUnFUCuXEE+w94sjnbVMnLWVVezt17G7yzD5FLrRJGoEfjlHyKZlv1auN9WXcA1nr65807GCwFDZKtGHv9tFfmwMhw8fNstet2qllTcH7wGIHK37RTIKlt022GeeajfkODBjzizsmLPp+7Lvw0OCRmPQGzkB1AEF7hXc55245O/t2QuuqpDynTOvrj2zruLm+sFjcTcD36e5d9H6kp/J7ahsdmC2cKqTQu6YWcXZDI37gfcY2idHLFP5Wdj3k0g6ajXJ12WdSFs8t7Hi5+D658NwJwopvzQM2v17eB18r3e1xShUapZJppowlYLViW6F7jkYoz2Kk1bclskVH+YOUjfHEmb4yGnFajpd65AHcfazQ0u8M2/fMWtFkjRCHqyrOEylMgzGNsJMsFyWe4oRJmVdHL5sTmeh2f5lNaWBB2ZrSgAhWECFuR7Pu+WWWF/KGpHXWVZgroQmODEgMRvxip9pYOkkFYllNDlo4Uodvq9yPUjWCbWk2V119PpuT6b6JjjY3AQqfpgr583X/hs/A3NkoobB74CxGRYLeQJyCs2hu5iY7OEiIfE+yL7EtO6azNptS+gHFwaetHih7YENJRj4lpJdiwcScS0ROhq8BbVocpOj9zczMALiShZjtM/AGXuIFWIXCR5/Ys/mFHImmTcZ9u3uALgQGOEBzcFCwDdIR31Z0JslidmJaKgjSVxTjEhrTq3xcdmh96McyrFpkwdr+BoE2/DvA4TYZPa+uHPhcaSeTZI4d2Sai92XUkAnwQ9n8O3t7ePS5csDNoEWru/zFcadgcFLaT4ZTMYm9uMjAMDznkxYwCo9t7kB8qCF0vbY5Cc1TDUbrJQaI57fra1tbVguV9Q9wRAuBd9x86IUj7ZblPuxMbEgbQ6FuDHcCFQ4S8GAio6FHJE9SekbixjKLd0iR+eGoYEhxFesNzYWQYKoz94dAhWra1i8dFFy+YNHqKjIotePYP7AQUzNzl2nqCDjVRZkHByQ/c/g50ptEKbN6+6fVZsxAZUAVMS7jBcLob0RC1Eic8wG6iZNdFYshwupTEasAjaVHFjQ75HHREBHOQutNtotOxcCwfJ5beCvvPySmjSCEmQNMqySm6QDFbxHfdN0GxlnbPLaeL7H6GDs+wEVvK00/CFjkkHiHPCSgS9WvSt+2rqnnH3rRZ8PRDm0t6yKYE8TvBhVRPA6tyxzpFGpCaRg0DDPF605HnjtG/CGt78XqXQBqQi9txNI5BJodDvymneggJ+RgwIOYchKbI8AFdVSEaVyGaUigYqiLBf2d3Y0NKasd3trWwAkrZ8W5maQG2Pjn8fatV1cvrSOSIRWLgT3KLmxYeIo2DD6Zz2GwXN8oGKQRDSws0eeUxWDylQ0pizZRvwie1SzHg54b1BU6OVdahwYy6ODMr+eDlTY/zlQYdoDARHyPB9aPzlQwQduYLVyQz7FYNAWvDs5iFTB6CBw3AAxAmSUdHOIy2tiA/Vh1oazdsW6l7WL4T8+pLSl0sAXFYiBh2+gtYHiDr55YcbzR5Z7pVQ28Eyh4MYA4r1u4IMxm6RWELPHwrRdWaRzH6xxTJVgpPWhbdb1g0d/NgbDW52LFvqRLj7wgZ/EBz/4M5ifPYpelF6rzJlhaDFtOopiMV9bXcVTT30L3/jGN/DyC2d1lHx/Njn8MlWa5eT4ufAh82BoOMinsPBj2q/oGrOoDowfP69ce3gurKkahoVT4bG3uyNmp0I+BwBYsI+ym25gI+TNl05RyPIY3ndcJ4ZAhcc18ZnQ2RsZejoYw39OcYjPLKcg+VYTF+y0+N4/9tYfw8/+g3+AwsQ0cokskpG4lJSNPpnywNrqCr719a/ilVfOolUrYfnqJexsbYp5ly3k8Bu/9Vu4804qXMhsa6JS3UGnTQXmGCbGp8Q2/t/+l/8JT3/rSURBcF0I3gCoePePvwNvePyNWFg4onPI+4LrB+1VeF6z2ZxIE1KAxuIiGXCv5HVg000f+FKpiESM+0UfFy9ewac+9adSxikk9wcBFWxCqEZL0IrJVBXeSPta4PeFGqvQOI0+R3bq7Z7gefcmuV5mtobVYU7ecFWR1roRpYbXhfx5s/WyDAi39pKEPmKZEmqcgjqEJBM2Y1wLWp0G+rQ08qWHzTmzswLz0Ne3wTNPtlgAKvqdAH7oFg2gy0DhZmCGD71tiBGedXryk+FMFmanhePHT+FNb/wx5PMT+MqXv4pXX31FwccMNyZZgyx2qiq49jIuVOdHtp0hmynUtH7O/ffr1q8RLOb6NZuAtzW8nkuhXI+ABui4Pb+Da2bIoyBQIUbgiCWa1R6WZRaJx5AmUJEbQzqV1V4di/YxPjGGxx9/DOkESS1ddFsRscNfevlFfOVLn8d+iexE3u92Tnn9uFYKRA7X1xy6hmvfKIBmfzZ2XzZDZYA9GzyftOyZnZvFysqKrgXrEQ5WzFqJA29TVPi+Mlhwo6ZYJrDBHoHWTwa8MOA8IvtGXkeCT1yveM2k1shkdD9Wz22gkC8YgA/a6zADzOwq+CzyMxCoZqh1kwSJegMHDx+Upe3e3q56ikwmpRyhAwcWtBbk8jnkxsdF6JGNSTKJ/Y1NbaEcxhnhoieLp2QqqxBo1nDprPUPrO9TCdp6MlyZtVkC7WZV3IdCgWsy101aszJTjjZBCawur6NcqkvtYMcexf7+DiampzA9O4P8xAQWL15GtxfB/Nw8nvrmdzA5NS21SLnMIVVCQIIYu50O8oUMxseyuOfeOxWqzr3i2tomLlwg6clAVp4X1nHZXFp7AoHvBx58CGQ1L11d0lCJw0xnrdI+66GHHsHE1BTOv3oOt5+5Q9kMiRjQrFWwv7slK6RklNZdfLZSei32f+wXxKalpzyV9r0YXjl3GaVKC+0uhzr2EJG0w587c+dtSCcSWL5yEQuz01KnXbl4GfFUBvtlKk3GUaqaOpb1JFndzK44dOSYsme4HlNRUS3uA90mHnrwAalrGEKeyuSxvVfUe1L18JWvf10scRZoXQIz7OuiMWVO8F7aK+5pQEhyHJ819xsnaamQTaJa3MZrThzGW9/6JmxvXMPa6iquLi3jjW9+M2rNFhavLApE589RwfE/b8cwbd6iN79unoEf6hlY7zXx9yJXkSOwTAVkm4rqmLICalSp0wax31b5c+TwDGamx6WInj94UHXN7tYOisU6dglW7NfQ6kZQo4KCGT/pJJqdLio1y5HgAklb3QZZ4AJM2es1pWTjmjQ2MY7Dh4+ILGE5B1ZUct7i5EX2ZnyemT9BW24NgjWDsdkDZ0RGlrI9X1yyYKuo4b/PoEJ+g9j3wb6P6yqH464wECBBADXFPA2zEeea7XZQTgbhZ3dlgtTk7CmkEnOyiOVqOKGC9RLBYa5N6u8JEHiQM0mACct2Vc2ufAsDKPz92NNoNhZmN3w/9lcEPbj3+lyB+4ycCkKN5zZUqhGkfqDVo4VBD+qSUNu77RDPtds4O5mRpBzLgh26e/C8sDaimwn7LKu9Ql5tAFQ4kDd1g5MvbL93hQl/9+us93U2n5wkoroGnAOe/ezE4Jm4/S1bun58f//i8ckBhqTWbseyToLFqdWFFthttUkcPa29QX0hgow85a0W6YZ5IltkByoi1kMLHNF80zKo+G8GjhjQpllVsIPU3kWCL3M61LdanavZGr8v5J7x+9jzOUGP95pbfXkNL4eakNXI2onXir0AZ1zKHonFRa5krc3zrU7/pqLih7qO3nzxv4EzcDiES7PgN8SaBSKlSIZqsugdDjVtiN2S9VOQwcn3zZpgWyRj9vPBv5eDMLJR+ED7YI1NiLO+tSgH5rc31SzaiZizoLUFwYaEfM1clswty6rgsIA/OzM7q/aYi/f+3r4QbK4ZLK65IHrQNzcFPsqNloUNcUhMcEODRcnrTYLFBVQIetgkuHlxEzClRkB8hW6aFM8CiroWABkaMAEVQp7N4oLvJYZem4oASvBaej8uOvTn52bNooCLLFmaPN6d3V29J2WDPK9srPhz5hvoVh/fe9NomCHrpyGTUpvJAO01pJlWM7LeisY0bOFQ3BZ9hiibZFBSe/kdtrXw8nd+LxsiYwBy82HRzZBa20C0mPcZFkeZJhdQC4km3s2hwf1vfPw6RcV1QAWZW8xA4YJMuy6qDEKjKR/JMHQbBSrElFNuim1y3LAW5mdNUSGg4tLA+olyeQ7f5+YPYHbhgFhOCv3rQ7YBNwIVjWpD11VWNQHN9oEQgYpkrI2nvv4FgJtG30JPATtWSk1UKEhJQH9gY60yVK8wMS7rEA66VHS17NwJ2OlZ4C/vLx7n7s6+fJR5f5PtdvY5WlYkDaigJ3UyNQAqeK+JWR6Y8ub9PrRycUaDP4vKkwnPlysqfDCljY8sjWC9Zm4QBlQI4WcwMRVOwd7K2eleKPQjJhfVM8XQcJ4/XicOgpQfYyHMrXpTIAULMF7raqWFU3fcjTe9433I56eQZMhpMi6gotnroFaz7BmXeNL6idea9wal/WTQ8u/l0j6ottDvZXo576NJxZMGC7vY2tzScUyOFXDwwDySGQKeKRXi58+taq1Q3r0UYEFeG4ZEKqxCYO2gyBLzwuwwjFVCoGJYVPn5caCC59ZZuzwPKoRcDTVi+TM68BodivmTb8NLAyM4KFKRHICKULrYEJtX6waggteS3yvfVxVV/tlNeeDvx/WN55dBYSzKXK2lQVbUAuoKhYJ+8V7f29uzgqxn4WYqGnsGaJBlKgAhZKz5wMqfK3tNY+t64e3DVP87X1sFvnJNWijt7RsTh2tQ2Cv4fKiQDsCFsTjjA4BiwE4OfqN8Tka/fE8bPf+j53xYTPY0/Ea0i7vvvg//5a/+Ixw7+hoFyxLoIkjBPbJU3NeauHz1Kr71rW/i7NkX8Nx3nlaDxvtQLNIgF9b9EwJt/XrqvpHSKoTChevs7GwDVoL8eeCrakW3NzYspu3eNTn07s6WVHw+BB9lsX3vYHK4z9v9bQMlPd88124dxOFTh/cP95lgVRSAtyEQYU0jgQpFVRBMCoGJXPP0q93Gvffdi1/69U/i+C23gQnaCa6p8QhakSjW1yp48cUXsHj5VVRLuxqMvfryWSxfXVSgYCqbxC//V5/Egw+9Gd02VQ4tVKsWpk1FxeTElKwUf/uf/ve4cuF5RPoNgODiCFDxnve+C69//Rtw6OAxA5U5ZCNo3mhINSQVYiqFwtg4JqenZVXA427UWePkpYrk+nRtdUkD0YsXLuFP//Qz2NnZkuc+90c99zfc6zr3BBdCqPWNQIUP5/m7mrUQ4ji4f0ck4qNAha3bbdRLleuACldU6Boq0HHUss3UDHwvfg6zBTX2vZkmWi2idlsYrD23PVpBNJtgRgWtHxH9XqDixntMrxFsjQjo6/6i9aFNIQZfQ7DAVK5+P1rDbCo+Kr1IZrGMFdqOZnDPPffj1tN34Omnn8XS0lVUa2UFmnPdymbyiEVTYla3+pZJ5l7DJrO3PWB0XfC13wf6nlGhNSOw+rxhZjC6h2nbM/3/AVRo/TU1qStj/XnzurlPZmw2q4yKTNpqCWaf0Ory0UcexAwH2I0+uq0Y2o0uvvjk53H2hW+j3WEmlBFT9JoRs3pl3Z1MpW1Q4uBJACwEXIzsCWbtRqAir9qJaxOVK2fO3KoB/9WrV4OiwnIqZP3UbuueGN1brGbkumW+0wQ+SNJYX1uX2og/G01EBPixjjTikBEyqGxQ5lcqheJLK2r0Z2dmVW+Y1YSFsBPsEhhPBWO7q31wY2MLR48fE5Bcq5lVIWtBEq9mZiaRSsRVe1+8dAnHbz2tz8V6ZvHyFZEcjh87adlYzTaKJdbKHAa1cPnKJSkmaE3FwdvBhUNSV43lc2g1OGRijdrA/Py0fidj2cI+aWnUQ6PZx9b6NqrVJmZnTRlcq1dENjp522tETjFLlYRsW77x9W/ixIlbUCpXFWjLdY4qWPY7rP8IhszNTSrknOttpVzF5UtX0WwaCUYEpD7PfVyfcWV1CVOTM7jt9tt0vbY2t0F7xRAbKJCHQMVjj71ONrsXL1zE6dOvkbVSJhVHs17B9vo19LtNsLTOppOYnBxHp2l2KlKrZDNiW6cyOdn6nX3xPOrNCOoN5p5B9TwBKWY/3XnHrSjk0li8eB5HDy6gtLsjm19EE9jY2RW7O5cvKGfmxKkTuLK4hO39smy9CBRzX52bnkK1tI9us46DCwt6lje2tnHk2AmsrG2gXGsgx2t9ZRExErQIlvRCT6Cw9L7AaAIVlvPUFzBkzwzzJqo4vDCD/e1reOyRe3Hm7jPYXbsqkGdpeQVvfutbVUO++up5XNvYwjgdAcpV/LvKhFbPm183z8AP+wyw/39w6+uI9mKYGRvHwtw8piamZLdWLlVw++23SfFVr1bQ71rezOrasu5vOjsUlSXYFqBYrnaQKUyiQtJpv4dMPovd/RJizFrs9rQuyw0hODLQhUF9Rsh5nJyewtzcnOyVWfd5HTBah2qwzp6ZzP9gMeTqSy4i7EdsbmWWQkY6tVpI+28glXKPclKSz3a0l7NOSNCyu27s9ZBHwD2D/8YZFT8P6zz+zu9xEMPcQUzt50oIt6Hieyv3IvT8A8cIDa+t//CsC9aUTgaymsAyzzyMmn/nHkKAl79zTefr8X25BrIOc1DBhv/MGKVy246ZGUBi/GezOg7t6yMh3LJBFNBjjH2eO1MeMng7pb5QpNVw7CI6sg9UFohdX+8Z+Ge+r/1byLkK1tI+rxHtQXmoZgfGetJyI+xL/V3IOGT9/Pyfjw8eCwIVpl4zJwKba0RkYSqXFv68ZnBGbuWxKpw82CdJCUOwK5BbB/kTA/ukrrmmBIKsGrCQxciWVESOuOW8cm7moBbPEz+D/axlXHjYtytvpIjkfLVnynaRXtsW1u7ZK+pfA/nYlBZDG1U7x5Zx4aQjfU+3N8gRGcwjbgIVP+yl9Obr/6jPwDyROIIBAeHkYku2CIf0fJhoY+APjxrIBDeI4EsXwqS9MVVxJ490y1Pg5kG2Zpo0m8DApAxwanpadidqfENwokASFuvBmsJeg0wyQyS5QfHBnpyeHIQTra2uyVuViwgtFnyhJ4vaZWmS2gZJHDc0MTfDgmiLSUwNKcEGl21pUEtGf0CfuaBKnhX8tZ156IuhBVfaxuBDXrGxQqixIbKBBUCAQu8/DOQ2BQiZCBaEzEVJYAuHlzoPRF4t7I0INxd3vXfYpLjh8lppGMU/00eRKhIW0qHZd+kgAQUurESWtfnSMBcQY4HAjxD9vg2KBARpcKml3eTkQW2jxlx5mV0NKjkQYJOmoG4qKjr0pAyZC1RTdFsawnuYtg/fHFX3YQuboIGiQgi4seG4wYiZTGZcUFR4AWCyuLZCCc0rsIMDC3Oy/6FcdfHyZclPDxw8jEQqo4Zhem4BCwcPIpPLyH+TDBB5BGsjMMuVZqeDZq2hc8LPyS8HAPhnKgJy6QiefurLqO/vId4TJ47JHEFSaKGgPFbJHIOlhuy3UimMjU2oEaZNAa15bNAHBVRLUcFcluBfTjSd/7+9tYHvPPVtbczOVOSz6ooKFi4OqvAzmprBrjF/92GBD1scSJDnYrB+siLABp60ryJzTGyNwBBkRoXOOdeOqAEVfG0VKgIlmO3A4+HQxAY7NoTlpspCwVjLsgpjDotscRh0WxXQSJew46dvx5vf/UEUCrOI93n+40hkqXJhCKytHRrqdjryUaZEn/cbFRUCKmoVZV7oV4Wh2mV511PhxXtoeWlZKg4e8+TYGGZnJjA1W9AzXql2cO7Vqwqj5qCZwBbRNw3/w4B2dFDoIIEBS3bu7P+Hqh+efy+gde4HyiNeawMtg1O9/ewPACocZPK9wodk/ByyAxmwoc13PJSAoRkw8EHFG4cGYtPa+sEmwupIG0gPC34DVKm6onKBwKrGcME3nWAOWbAsLCV97vWwS99uDg2Vd2SfgdYYXCeN8ZxUkJmfTx+0DoCYIH92YIKFr92TVtLqXtOHtUC9/d1dHRPXuUh45hyo4D3Cn+WgwRQVxm5xtooD7Q6wXTcRDfevjneEXTx6LXUuqR5DFxOTU/jHv/k/4L67H0Eb9M4OKhnmC1WqKO7t4cK5V/HUU9/EhQvn8PwzTwewd8j+1bOqcFmzcfIBqV9vMXn0PbQjJDg6tPjSPkTP0vAM8/zxewa2ZYGBxGtEgGJvd1vKMF4TX099bXAAafS4B6BJkGA7gMT7w+8zPiuuuJGqJ1iAmf2XMb/4c3z2CLhyxeTebENc85hV89btyEbmV37j1/HAI4+h34kgFUtovVnd3MbVqztYW11GubiNWmUXe9sbOPv8s1rvtf/0unjru9+Nn/rIxxGNFGTbUquXLJspm8fExDRqpSL+6X/3m1hbuYAIuMYNFRU8iHe9+x14/esfx9EjJ7SGGZvJwDGqPLmeid2eSMjeg88I93uGveazBYxPTGgvv3DunJQFVFT8+Wc+reE9vee5ZjEzyu9zA5FCzgFXT+4VrqiQndEQvLPObCgxH71OUh4IvNQ3DayffN2u0Y6JuT43WD/x3qIPtdUoQ7DC1xwp5HgdlS1iWQsCKTgH5vtx7QnvR4YaGZUaMJOwQEVF+EQ6Z+FsD8AKDgoixpDUOsbahDWHvaI9s3rDAJiFbIXhemv7szfM3Ntl4RW+n/83OTmL06fvwMbGJnZ3d6SmoPUY64NUKqc6p0mv6B7ZlgQquNfRo5tKBctucHDCTr8dkdZM+2iDLz8urVusbeNWW9n1MALBUFFh974dXgfcY82Gr2MWfQFQ9vtEdUrIdkllswqGZ6io2RH0kUoncM/dd+LUyRNoNfrotWKolJv4zKf/FIuLDJzfN1tDVzrBwtaTyYysGLT+3whUDPI2uLcFOz8Oa6jkCMq16ZkpnLnzdt0bBCqooqBS4UagYlRJIxiKACBtJONJY7u3O7i2uq5zRTUDz12pbEAFX4/KalNAZPXscRBDoIJ1xKGDB3W+OGgiQMDn1v2gCQ5xmM96cf3apsKj+QzQZk7rJPpSBUbQ1dCegAsDsvlss55J5gtYX15WZpuykgmcRnh/pFCu1jVI4X7IrIv8WF53LvMrtAeB6r8ier0WDh2cRypNOwpTbWgwJZVfBDvbJdl1MeRWJBZZx/ITdfCaW18jUJS9Tzo/jvXVdbz43At46OHXKv+Gw28CCgQr9AxFqMZNI5tJ4PiJI1LaEIhZXl6VqiKVympvrDVq+hzMlNja3tSQ/uGHHhZAsbm9o/PaCFZuBE9Zo99//4OYmpnG1SuLOHXihOph5sJQubCzuYZUnGBlU+HXM1Pj2m8EiifNXthS7KJAPIMXvnsOxVKLUBUqlbrszPhfBFnuOnMrYr0WttfXMFnIIx4Brq1dQzyVRrXeRj+WVJ1J8IQDt1qjia1d5o+cEshEi7+ZyTFUSvto16sYy+cFNFVrDSTTWdBXrIOY6n2qHsyW1Zi7DGHnhSZopbWzS9urhtYB1hq8rzXUS8YR6TYwnk3g9Y/ch8MnDmF/dQVr11axtraG177+cbDsWLy6hPT4uILMt/f38Ae1GV+hw9LxverN4Ypy8083z8B/3hl4uPgUOvUushw012lhl9QMhvs3SW+HDy3gyKF5pBIctlM5GcEkc3h297C5uYNqpYmV1R3sFGuoN/voc31iH0elqdwsLLPLc0VZJ3HvVOaD2Os29xibmJA1Hv9Ne40yC6nq4Dpo2X0czqs/CcHVInbRxSDY3nJoy7+7DbkpK3yQbeeJr+/ghIK7g/Wx+ngO8wPBlLW09zzcl7nm+iCYe6T+zLrPB92sq5MMnLZBvoBm1kRaN6gatIwB71W8fhLAHMKoxfK3ED9T6jbN0tn6ELPt42cia557MUGS0cwLuQhQMZfPi8TKPos/y9exLFkjmapGCXWiwpqtYLnO3lcExAAqqIYKuVgCRkL+Ac+7A0+u8PR6i3Wj51T6OfKZgH8O1W4BYCKAwj2eyj9+fn6PqRAMtOJ1Ien0pZGMirvesTdwMxlVELN34L3LepxENC6kPvSX/VIAZvzJscwKA1XMOt7ILTxX6kOZwxSCwnlduQdbRplZN7HP815J5y30qgZqWLC1erSgNDHKUbA2DfejW4ixRzFFcrCRD2p1zcNCPy61iEiPBs6wP1LNRKVSw4i0ozOBm4qK/7w18uZP/y08A4fYiIXNwRc4Dic1MNAmYrZM3ABM0kY5fUz2BxpKq9kKKOEgnCiElqqZEbStZkuqgWgcDz3yEPa2d1QE82fJpCYaqWEJw5wzaXkiij2VYWBcTcNvDgH5f7ZIJfRzLstSIHWtrmGHcgDkF0+GTkNvb0Grpt7gUs2FRptV8AD3QBrJxYN3oDXjBrzIqiWwFvlzfC82ND6E5sDCFy9eZg0NwwLDxdfQavOXk+qk05V3LofNfD0qRcg65DUwf764GDveBNOzlwW+kGktvFGxh42hbMoD7XbB1oU/L+uswCwQs0yDBLPaYrPCnxkr5PV6bFK40PMzigmgDc6Grv4aHOTz/IrN5Cw7MlDVodtAwAZRDVku8Jr0KCWNGLO6zjC6Xgd3ve61VpyHAbZvOl4IjAIVfp3ExKs19Jndc1EDx+ATyffkDWkqlo7YIpTDMdNjZWUJ44WcgAo2N/1oDDPzC1JU0JOXoDuvAZteFj+m4rEw82KJrAVjUzjb2QuNHgP/4rTzeAXXLr6KAi1YqJ7g0FLWT7Z58xqxQBHARUYFhxAwFi0605oAACAASURBVDL/n2AFCyiBVLyW7oUYJKs8ThZ6vGd2Njdx9uxZ/RyZdQyCpqIinWL4aF8sPj+3PsDxYYpby/ggmv/vHptkwko+O2Ipw/cl44PrgeSZvMI+UA+AUDfaHxRkzsYYsrKtuON7uB2V1DMcQEVt0E11lbIuqBRiQOLenryOxyfn8M73fARTU0fRj9IGhOcrglKlKgYQiwfu6QyiLu8Xgw0Rw9yqeh2CVM16TWxE/p1gZLNZRb1axfb2Ni6ev4Di3r4+2/TkBAqFpAJIeV0IhJw7f0nWCxyQ887mmuHn0Qe5Prw2FojZBdhwl3kpvtgP+XJaP0YGiDz/sioI1k9+3bxgHr7PDRuHrC2GX/59Dp7wdX3o7ix3vxf8ueXvzmrln51xZEW352qYfQbXi3yhENaBHorMhKjVgj9qF4lYFxNj47K4SCazYvFs7m6h1qxr4EFfUL6/s2r4OZ25zVBNZ8N4YWvfZwxY/97r2cxRG4yqqKPXZwu7W5uD9ZfPtysUnB3E6yIgN2FD/sFwdGT4Fg9WS6ZEM2BWw0nZF5mF14A5PZLhYQyhiLITuHf8w1/7r/HYI48jns8jmk3bPkqWaKOtfIpzr7yEF88+h8XFi3j2O98csIMskNbDjw2sujHfwa8j9xBneQ/XYi+GjeXuIKk/17rmZLSF8Diet/39XbRle2jPqn+N3ns33oc3DmplixhCZ/0e5u82jPRhtwW7iyzQ5vCXA8ysMeHCl8INyYIT4M9moo2pyTH8wi//It7z/veLrdeLkMGaweLiGra2iho2d1o1FHc3cen8K/jG17+Ga2srsuvg4OrkLSfx8U/8Eo4cPYVqneoGrgsdZMfHkclnUN3bwT//J7+JvZ0VIMbQXWf929T57e98Ox588H7ccccdYu8lKLsKzwufW+5LPkQms53MfO6T3CN5nASNOOTrd9s4d+68Bmdf+PwTg4BI1Vah3hgdeg/OCay28v3HG0/tQQJOTdEyCjLx8wiwuwHU8HWB+2K9UlFtxPWHX5694M+l1IkjChlT5pm9l9tV8h6z6+uKip5CjwfWcAT6aZMlZabnIdiRjT5/+vuIZZIA1EFQPMe7N/gpXbcc0k7TBosG8oTMC7EjLTdHwD33Gg58Y3EcOHAArU4X+0UC2BXtTRxq275lA896qxHyfdjAMkPA90bLYfAagPerq+D4/my+/cul+IO/B5WYr2W2loTMGdXaAYhhDRKYjgaC2trjIIWv3b5+cziey48JKJaCjIPzRAKnbjmO++45I0IBegk0q1F87i8+j5dffhatDn2zRzIqonGz9OK+GpQyAp0C6O61lh2L1cR+HPw53SuxKE6eOC5wsdXqKo9F1k/ZtIZeXoNzzx8wLAMoLmA2YmSeTCqj67V0dUVqI/4c61kHKhRgnzSiBp/JeDyFbCGP0ivLUmdSYZ0i6YTkIPcBD6xbLnEEKnjPXllcxKFDh/QZ+R5k+NOuhLVIFF1MTRQwMzujoNlsroAccy/iCXzpC19U0PWRI0dlKUprCe5HrEsYtLy+sYbx8QII2iRo/5lIod1siUCxtb4moOK+++5CLhfH7OyE7l3e8wScev046rU2djf3sat8G9adXQU55wpZHDl2BJl8AWtLS1LhEiR68ktfxaOPvg6ra+solWtod60a533RadYwMZ5DPp/CgYNzynDgc3/1yhJ2t/cRjZkShudqapp+4H0sLy1JbXb77bfrPqQigGsdLZVUC3ZMUfHggw9jfHIKy1euGCDWbCARjypPYntjHTSDixIC6PcwOz2JVNKAPrMfjKCrXiyCiICKC9jZqyNbmESVilmRJ2g5G8OZ204ijja21lZx9NACGtUK1qiUyBewV6yi048qUJ6fjee40++jVKmjMD6hjAo+89OT4/q5TqOOwwcPaJi1vrVrAEenh2g8jUgijqsrKxq8EqwjiYZrWb9jeUnKMqEqPqi3OVjlueP/RdkHdeq469YTeOT+O4F2XQqOYmkfV64s4r9469uwvrmtz3P7gw/h3EsvY79cwb9atkrOAWoDY69b4L7nLzbL+tsOaISJ2w8+lJv/+yM+A4+Wvo3x3BjyqSwKmTwSsSSKe2Xd1wR7SRpr1EvIZ6OYmMgro+Iw15xCAXsbu6jWSCSMYXu3inK9jXq7izbX8DjrLTooiJpmOTm9nmZGvJ9ZZxDk43PNO3dickLr9GjPot5pxD6He4/IeuEcCQTQwDbsk+xZBZAPvfo5h7GBrvVirGt9mO5qDZtnJdR7OpnDa19XnHr/5EN2r/G8/vdBs2dJaA0fUUP7Z7BiRx9xUDeqLgsAjAMKTsSiSoHKCYLwmhMFa8xRK07v1VS3BRKiEyidOCT1YCA4jJLAwmKjmsLBe68rDHxgb8V9c5gLqLlZAIucKKNj7XQG5FjOrgTcsw9SH2GOAiKIpZntRgIJ7fK4v9X1Mfhnnxm4SkKzSNldG0F5FKi48+07eo2BQn9EmeEEGtYssnUP9lB+HJydCFPw8x72XL2vymi7X/x7TG1hl832ZyOLhOpV/0eQw8/DqNJdqvUBkYu1rP2U2VPZOfFbQvcRwSnuXUGlw2vNv+vaq+4zO3q3gPLreV0+8Mg6chOo+BEvqjff7od/BhbYNHDx58IRs4Es0Vlj/BpgYRZQtAMg6sfvb6m5lhcscyMkWYupaFdIXaUsBrI91saic5akB5aSJcWHPJPOqjmgL6yhuB2xevjwsnnmQCxXyNmmwvfjYF4PNUOnGQBnjGTaK3BzkdUTpVy0ftKCaAF97unLIZodnyHOZDnSl57DNC4M9J01JN8GeRyKU6GhhoGMqHrdwIGwsPhiwpwBQ9VpO8Dhm0nsiIpL3qZF0BYcLnwEHvjaBF64QPGYDSighZSxhxv8d3optjm4sc/D79VQjA1yaCTdCsSteTSM4kIdACYuvvx7IpVQaJ4Ym92ugKJ8NmdMBjY1wcaCTEL55QnVNsBFvqqyVOCxmNyMX7k8wZaU7MBaLQOFGIrI5qrb46CXQ5SW/l8WUN0WTj9w/6A49xDmUcbCQP4W41DfQqZ5rRQ6PKKocEY0X6PZqmtQP1BUzC+oObxy+bIBFWP5oKhIK39idv4ApubmURjPIxE3NJvFlW3uzFOhRQbvZRvifT+gotsxBtna2iIuvvAM8kTlGcpF/gPvgxgtv9hIxwdsCClIpEQha9TuVykj0jyPxtiVX3EY4PngeGdnR+GU15ZXUSzui3VI9kk6afZPYgNG+/Jt9saH99AoWMH38dfzIZTAQV00YxR48ePDLw4COLgQwBbYvpTB895SxkrCABc96UE2OmSAm28nX5fXaMBGiVlws/JH6H3Z5IDQALLSPkOvK8jmx/COH/8IZmdPoheJIZlNIpGMaEjeaJq6hA95q97Qc245N/SobGoNITjRJfDXoFKjJouXSrmI3Z1trCwvyyuY2Qa8HjOTk8hmohoC0K6LXsznL1zWGiM2RZ9jCx8CW4M4HPyHoX7fgAoDGWhD5sxfsy/hlw97vDDUYCuwb7yAdGaLFyNeyI/uBKPM6dE/+/fws/n1HfzOYfKIHYxfL/95L4h9gDRamI6Pjw8YQjyX/plNQdZDJhnBeD6PscDqPXPXXVjb3MDL587p+vA6O/jiA0oN2cg8Cc+Wq9T4uQzssWGr38ujgAvLR2Hi6oVNmbO3vRXeh0H1dvy8tt54qGnhkJU+vIE9NGyKjH0uHDew0CPke4vpEsLUAlDhz483Qvq8ki4T1VDNi5/+yY/iQx/4MNKTk+gHJRH3l167jyuXLuHll87iu2efx8rqIp596hvao4yRRFtDXie7j7qBMe3XdXTw7EDF97s/KC3j64zeA/4aPOZuAJVtD9hFrVqxYL9Q+Ov+DveKqw+HFrJD6xu/j1XIh8Lcr5ffR/asWPOiY2Ij24+qyCebl+CyroM3Avw9ANDcQ8gE/sjHPoKPfOyn5UVO5mskksK1NfolV0VioIpqZfkynvr61/DcM9+RSiRDL/lKCdPTU3jv+z+It73jx1GtdbBfrIMuXSmypcdy2Lm2jH/23/4mmvVd9CPc04b2RPzzu979LjHE77zzTtUbHljM43OgQvsk1/qshQZzLS8WSwwZUW3VbHDw2cfTTz+NZ555Bs8++6w17oGdx2Gsnze//wfPO9l8Qe3qz7Xfv1Rb+ED/RqBCzeyIqmb4HEXNdqDZRrVWHQZF61m04bMsIhVybixifzb1/gpLD1ZQDlTwd3V4Q6CC76fhbN0ssowdNhyu+bozACxCCDXvfbeQdJbjINginBQ7/jCuCypcB2yGew/B11CzyHKRxIO22SHwOqWz8uam/zVVMNwbXSFaazY0iCVZgT+n445aU8p+napQnh+dh+DBbOt2yNzwzzkyo9BuEKwdzDLLGmG73qZy42toHQmZFIMwyHDuRsFmrY8hp4v7K4HkTDanz0uggteM4ckPPXiPmf614+i103jl5XP48pc/h0qNwK7Vx6bwsJrWgQpZDIzYXF0PTtrrD9ZkKQ4tWJT5FEePHlHw8uVLSwIAWB9S4cE/83V57/t+4/cB62bWBPz8BCr4sVaWVg1sYj5AKnGd9RPJUpZRkUI8mdGxbz57AZPjEwZOxSynRLVXk4MfeoT3jLgke1vg/PnzslmllSmZiQx8lgIwShVHDIW81eeVKsPY80hTsZJK4y8+/VmUimUsHFiQ4px7Bc8FMw54/RaXLmN6alI/y/6GYALBIg7y11aW0G7X8YY3PobJiSyScqPtaz1kbU08r1xpYmdrXxlTRlKpqq7hcO/Q0cNI5fMobmwKAKHF3De/8S2FUHNt5YCegC4zF3jc6UQUY3lmRCRw++23IJ1OimS1dGUFe7RqiSdRrdVw/MQxnLnzjHqAP/uTT2FmekZrHt9/eWVFNZF6QQ4fW03VQw8++BDGJydx9dIl3HL6VjQqZQVdF/f3lFGBThuZZEy5FdMhSFwkrFQimOsB3X4UkVgaz3/3PGrNPpptbsIJPZvJdBzZbBKnTx7BWC6J5f+XvfcAtjy/ygO/m967+eXceaZ7picqzCgLhDJCEgIDJViMBZhkzO7aW14v5S0V7LrKYO8uwl67WFOuWvAuBuMlCyVQmFGY0eTuCZ3j65ffve/mfO/W953fue92ayRkm7JH0G9qqrvfu++Gf/j9zjlfungeCzPTGItFcfXqNakhNnYKmJiekzqiVKlgcmICjVYTe+Uqjh67Ay+8cEbrNq1gN1ZXkUokzIKL+UFrG1JYM9B7LJlRz1ikFTDfcLCwo1omGqx02ctQTcFQc3nSC0ynzc040O8InLjn+GG88bX34/rFs1hZmleuCnu4TG5Cr0cY9+BdJ3Hp/AXs1ev4lQvWR90MVNjCYJZ9X/v1rQlUOHAxSrF5pYMtL3Pwv8W/dd/aZxEbxJAeS2MinUM+m0OvY1SAk3edUG4OiR9cN0qVIra2N9XDE6wvlWuo1ZhLGEezHUUkkUa51kCbxNExu6e5BvHK5R7LGRHJAZpbkIhG9aZd2KD1E4EKt2ocDsuldja0jj0daxhZrQWVMJ9DfSpnGiKeGknCsxqUtxPqR9aRAl9CSDW/z/+9jvbewGpU61X55Y/hZzb73puvU/6+KyPEwg9gOxUOmkHJfjEEMgdbzqErSbC05gbH+kS/z31cfYy9DusUKlIcuFFNE+ZVZh1u5Ee+D68hvWcyZR7zQttIjNNq0YgTVEaYatn6WCOtGLiiWRJLmZA5yO+57bl/Nh27QK71/k/OCZ7bGNQSmrfdRHoKCvbQ17GW1WsGVwaeTxFvZd21r+Q3xSYVFaY449e977ZsVF6P7FeM/GkZHPzi+eNnZG2gPzW/NPKTW8gLcBCAZY8RAMXXDjZhvJ5c1aH6SuHhNhtVD8vfDeQHm8VFNecRATMonu0Ym8LYRiYEdSwzV3ZknkESjoMT8kTUCmCKyMcOVIS6UvMcAWJGIPdsXwfIQjF5O6PiW3yNvv32X+YInGRafUikJ+NTBVoIJ+auouF6n8GCHbvR5L1vDFFmHFDaz+H+7OysbnzaOrCba5KtWS6LbcKbzpo4Q2D5OxzKcvDMpo32D/Q05PNk0kkNjsulklQUJu0zJgsBBxb8ZDxziHj33SextbWtzZCNDgtuPpb+1AQCOGBjM8PmhxJwNuK5bFaPc/WAhyvRr95Z31OTk8jnclhfX1cTy+2DNkhkvJpKwIaq3EwcpXe/eTLquFGQlUWfYL4fLqi2iSWMmS4lgQW/kQFgAzWy4CzLgoxvoupk+7Op0NCNEmPK47pkuSdVyPN3ZNkS5Ise+CP5vxbU/eAeDYtZMGfSaso4XCMAw0JFCLpCB20zqtaqspzQMK5vx58LLzc9bt4EO7ioErQS0zLGjZsyRA/0oXKEskW5LKFULqq55+Cn2+8oTNuLczH6wzBbjVAAJfhzfm6XhPK5O03zjPYMBr+cidjznJMr7EDF8uKSBiUXL17AjevXxHAz6ycDKuaXVjAxPYP8ZE7XGwsSWidwIxRqH6ElGIc5xsJ0OyVnVshypkuPxShKpR08//gXkekTtAO6HFJruGH+yl4QOSjB0FWzRrN7w4EQ2TAJpAi2F2Hz5WsSpHjm6WdQK1d0v6RTKamQCFSwYBgFKkbZIXbv2detQAWvQ/08MMmHMtFQuPG6IlAh9ltQI8kmJxRuAi/G7P51IE0gXrDe4bBU12YAZLyY9CaP55TNGEEFbrb8k4HDjXoFibE03vW+78fS0l3oR2NI59JIjAH0OmXTrDaO56DV1rVIdQkzAXr9pu49Dl/3igUNYnk/MeSSgdq1SlnZFLR9ssyFBKanJpEaBw4dOaQA7Qa95C9clpc1hwcMXdSYLXxu/9MKXmPX0i+av2vHnoMsZ8Lu5x74efFC2Qa3puzyL//Z6GP5s5cDJPz7/lgDQ/cDvx2o8nPi58XvPYEF4TMNi/ugqPD7j+vcgZUDWmd4fVDFxu8RsLBhUx9jUSA1nsD87Lzk3N//4Q9jY3sXv/v//T62tzbQCUyR0c+h4ip4hzo71yyh7H7gzzk08c+2rySw8Og+pQYBpGA7v1fYtcBZrllh0M+CU/lE4TPxOGj4OcLi92NhLBcrFA2Qs9fh9WkEISvmh4NVV2JwgRPQTwCAoWpRvOPNb8PP/tTPITMzh0GKlkg2nGc4J5U8zz37FM68+DyuXb+EU08/EYZjca3x8diYgWBUchCoGO3rw0DDmgxbK/g1CoDp84BS4JFBYijkdfz5PvXezTqrUtpDubx3s/VQeJ3hQPyWgeUoYOLFOfces0C0Lx9EWgMaZM1az7gvmUKAQz4Ne3iAQ86VCAPhfuDek0hE8I73vBM/+dM/jYXlAwIqBgN6s+8JsKQCs1bZwwvPP4PPfeZTuHHtKna3NzXcJLuZKsQ3vvkt+LEf/2m0O8x9qqLTpqdyFrnJHK6cO4tf/oX/Gb1uBf0o1yMCFf45BvjAB96PO+68A/fff6+GmgzM5WfW9Rn2KmuE48jmc/pcvJ4LhaIsCQhI8xq6ce0ann/hBTz22GO4dPGC9hb+vo5leDk/3qP3upqdoHzze8OOsKkjeQ34+xm9r12+b8c/+PQP80mAgfa2uu7l/cbVrhmGvFpTZIo7vy+NNW/eztZcKVlQ96L+HrO8Gn4eNdGtNhq1uoAKTZ5HrmW/j2xNMBs2+1R2H/KepVLQSDQvr/Sx68yA4qHKI6i1dEz6+0MH90y25g/I5pjJZbUT60S3PlOt1mnrvuMQ1wYCNJ+iPQZfS4akeq96zZAa78Ae34/dZ2EdCfeDgDw+ZyD4DO+VsI6ooQ4DGt4DXHQs48U/u+0zfo3w/DqzkvVZRkAFAZgUOj2SA8awvLyIhx96QBak3XYE3daY1ESf+tQf4OyFZ4BBa3/f0bB9H6igEsjvAh8i7e9R+3WLgxU8c6zp7777hF6XakTmIJiiguAd73cOS1g3GgnGhyRqvGPW1HNdM99u4Mb1NZ1fETHGExr60tKNRCJmSXAYJiKI7KpSeOFTX1K2xf333YdcJmf2GSG4m7VtjrZsgwF2tncFpPD61joajaJSLqsOaNIaKJdXrTE1kdXzF/eKUuCyFhibmMSn//hPUa81BFouLR0IVm0GDFTqVVy7dkUZF5NTVBEkuT2odiVDf2tzTUDFW9/6Bhw5tIhWs4pUxjLumgREshNiLRe397C2vomJCdqC0paR5AfWKMzKSWL16nXMTs/qGhkbT8n2qdFi2OwYnnj6WakzspkMBu02Ttx5FM1WBSeOH6WjqY4/rYd2d/dQ4+dIpnDfA/cJhOO6deq505iansaJEyewtbUlmyX2X2RMcxBJEg7XJYZtzy0t4vzzp3Hi+AlZdxJM2d7cQHF7k7G2GHTbSI8nsDA7Q1PCoac69zbONBkPOoiM4elTZ9Bss49g4c8sPFrFdpHLZ3D/vScQHbSxdeM6Fqanpdp44fQLSGayaHb6SGcnZdtEmz3yDC5evqy8jjuO3yWrpUwmh8l8HrVyCdW9Eu666zg21jfx0rlLWFhaUT3JXJYSswJT4+gwJ449MesP2orEWV+PiRlcqzdk30ZVCa3pBFJzPyZI26ai4gjuPX4Ez3z1S3j9Q68WUeq+Bx/EztYuNrd2cec99yqD4/mz51DvtvFvNo3k83JAxU0L5vBOHUK0I9+5/ddv5gjc1ngAb64/hUQkjm6jjWgvhmScGYcpbO9QWRhV7TM/m8bBg4tYWllELBHF3MqyZgOFjR2UKk2srxexuV1FswvsVetSInG3YN0QD7lLssCL2ADXfkbHCQs75rpPy7i5ubkARNhchLUza/N9gN7IcBoch55UPUEgYnL+oblIy2ySuS9ofQoEU5Ebw7yF+xDfC/cSgiYiZISAaK7/TtJj3cGah7/Hv7s1phQYIU9DaqvwOUQIDYRRznickOf7tAMKGkKHLwEvITibjyOZlWRQt8hygEafiYp2DtVDL+Q9HN8PSba+/7rGnjM61nTq3UmC5YIqO26zpNKwPdRaqt3DjMHqUKvhZR0eyEcOhozOXPhzzotSyuHg3Gc/f9Z6EascRHqIhBDvsM8aOBByBEkC42NHVO2mZLdaiP+d+gRVfvbFjArODESiC7bxIlQE6QO/z3khldqetSo1aSBVcg3n3zWTEGDCXsMIVFLLUUlbr4tQIaCGoEvMciRdZSK7054Ry2RpKwd0e07N33TczMaTx9x7SM6nOGvgvumqW3vdcI/Qbp8kVYJgJMmMZK2w/hfZLxC+HGyxjE8LDGe9Z8fxdpj2N7MX3H7Mt9gROClPcVs4eFNzsVW7GIJJuQi4TI6P4ThmfmEWJWZCMOguHkO72Q4++3206TUYApG1uJou3gb8PXo7d9Q40ZqFrPV0Kilbm8mJKS0SUdrXpMYwNzcjb2eXi0tZ0O0G31YqJCIaonLN5RA8Go9Y+A9fQ+GlxlRztJ03MDdKLmZknwn4kA2P+QkSyODmwS8uykuLi1Jp8HhwsXfFAX/OjcQ3O6kNQpaADwYNfe5a8E8YnnHhswAi8wPn362JS4sRfuPGdQFBHPQRtOEx4TCDTHo9n3sghmBkHsf4mG14/Llvrlz3PaBnn0FtIdNkpbHY1pCgT7/cmqGyZD8KYCFazQGZqgJ772T7yfuR/n02qONrmVWCBSDyePOAE2ghwKLGqkfWHBd4hmM3taFxf2l3mrjvTW8YWkrxWPswm8ePx3LU45B/96acQ2kh06Ho8IGZKyoUBhy85xcXFpXRcf7cOfmYE6hYXjmIBIsMhmkvLiM3NY2pmckAVPSRy+VDNgSvEwJMHOYYmGaf3wYoww2+Zx70lWoBp7/yKJIdetoO0Bc70I65Kyr8vBMsoN0Nh6leIHnx4cwJHijPR9HQYzDQtfjEV59AYXtHYBOLBG58sn/iMIkD3gQLN2d+Gqucz+3HyYO0Rwfl+jlBFfqgu5/liDUH7zFee0MwjIOhwHiX3HTMVCM+LNUQVQwQDlUMKPMgXxV6AmOisnngQEsARdMGJgIq6J3eqMnr9O3v/h6sHLgnABUpxBM8DhV5JasQ4Gv0AjuD56vTRLm6i8LODgqFHexsb6NcKurYsYlmeG29WrF/V2u6dzjkmchlkUnHpKiIxcZQazRx8RIzKnpqYFmLUnUyOki0QRuHRzZ8IuOWQIXOF6g0cCbOzVGJtwIRPCYOMHjDeuu//RrwrWUUkBgdnPvPRwEI/pzXgQ8bR9UWNw8LjQHkvzv6s5mpaUxOT+k5eOyYCSLrpzCsjPSMMU5LBYYf/+iP/wSK5Rp+7V//Gw3kqWrx5/XX16BXqol9z3ffaxzckyVFsD/zgbd7u5OZqBJReQZ9lAqFYO3C9csGes761RoZPN6HFnhhajo6dKeHvlusuKJChTPXPRWfbqdjA/fheXK7mehA4P3dR47jf/noP8bU8gr6NPuVhI3Dqi4uXbiAL3/xEZw/fwZra1fx4nNPh+NIm62k9kRlOZC1oznwfoC1g6QsqsXqCaDUzcBZAFYGX8f6Sd7adm2SOcz8lvJe8aYhKK8jNQMjX7JA1JDagm/9WvXH8cg5++prr8l92TTXhLGEgbf8jLrm3N+fR4oAeFAaMNg6Gu3jvlfdh//hf/yHuOvkvQIqut0YdrfLqJNYMeihuLuFLz/6eTz+lS+iXinjxuo1Wbdw4Mzi/t4HHsDf/omfRTKZR6FYRafZwVgmg9xEHmeeexYf+6V/DPQb6EeZX9XTnudfH/zg+3H4yEHce+89WFhYugmocFa7ANtYDPmJiWBLyHWqPMw8ou8+LaloQ/jII48KJGUzYnWDARWj5/Cm+z00wQ5mjyoGzJLSrnOeEwK0TryQ5+9I2Lkaq1Frr25f/sDW1NqwX0AeHxc8k0cBziGDfhSoCIoKWqOpsWJYdsiJ4mfw7CGCm9bO3cxMHF1jWHTofgrZZnyv2UxWe8VeqTi81/x687VYfW6wnPSgiAEXzgAAIABJREFUTa/DzEbNvkwEaOeVn4Xh0wrGHB9XDeYNuQbbVuTp+rTn4C/7cxkkKUl+AMv55F5rseb1r1FggeuIDB+1L3qotrFPTVFhqiwNabSnMdPAkZ1gSeAqp9BsO1DB905FAT8H/1RUXCyGpeUFvOr+uxVaajkV49jc2MGnPvVHWNtkJovlRdmxtPwY7mW8R6WmGFkDHAyzNc8eNwSwgs92LpdRIOvMzBQaDapZr6vuT6YIVOwrKpzZehPoy3cSYTYeSUtpAVYEKlifa1iTiGjPISGGSgXmipCEZPUUgYwU6ufWsbSwqNNFsg2JRByMsFYeY/honaGpDOJOKEOp2WhpIL+zs40MldRUHNMClX1ItIfpqazsXTe3t7G4fECvkUil8Sd/+Cdo1FtIptI4cOCQ+h+eSQKjVA5vbm0oPHpicsryXGhcxCybThebG2ugEvetb309VpZmlZtFxbgpmLlPRHDtKpUkcRSLe1KbN5p1EWLS2TRWDqzItu7Ms6eUK8d94PSp5zGeykqFWm+2cfEK1QYZrS/JaAQn7zqOYnELR48exPz8jLKSzp29gEKhJNXQnSeO4+Chg7JsXb1xA4XdIirlGl7z0EPoddo4c/as6mHeF+ztCGJRVXDvvfdhcXEBa9ev4NCxO9Bp1HXN8ng2qhXEogxxb2Eim5L1Uq/NgRwfYdkofQ5t+kB3EMdTz76IeoOe8wRK+xijEpEJFrEBXvOq+5GMR3D9ykXMUAEdi+HG9VXEx9LYLuwhmckjPj6GYqmMqYk8tgu7CgqfX1jC5avXkMtNgDVMqbiLeCQiAJS13eUr1xFnvsp4ErlMFnsEwvo9WVZqGMmBVjQiZjgBC+67lUpVqkzty2T2ysa3i/F4FK1qEa+9/y7cc/wQ1q5cUID31saGVEarNzaxvbOH4yfvwSAexxOnTqPR7eLf16eHe2kQN42QUmz8+PK6g9tqhJsKlNv/+KaOwIPbj2AyPYGpXA7zU/PIJLPY3NhWLTk/N4tqZU/2uNEIbZp6KFdbOHxkFtkMM75IzCPRs49CqYloPI29WkP7WqMblEEk+Mh5wfKlxJgf9OVioZxRkoswUE7pzOzMMHOSSjfuJ5pHeJ0SZLyyQ3ZShzLmLJtivwbdJ+xw3/BeQ/Mdn/P48J39Juc5zLJQPoAphPn8xq63wbFCowOg7v2rg+t8XWUOBVWDHh8svPkZSMzgfIRfQzKKbE8NONFAOqhArIfcz3fwPZGzE35OJ1BwIXClAp/D7a9ZT7i7hc8obHBv7H+ROGRf65a+ZnHkrH5ThtoX7cBZb3lf4wx/6xVM3aL6JcwHzMbcbYathrUZjs3ZlKUQ8j0JAsiOlGaAva6AAD6fKxEc8HXylWVC9G+yfnrwu0pDtYvNsAxIIrHBLbz43LKhJeGJ1lNSiwbL6kDglUrC3QUIDMgCLCplnEjZ7ZbqCxFrBZRZ7qORkIF4lCoYI/fqPAncIpG4HeysrNa1Y8AZAxWCzJII8wER9KzW42PUj4WQbQEZvFZZTwcLKX8ev54MqLFzZiRuI3yyDpU65naY9je1Ft5+0LfQEXh4fk6DAQ2SGfBM5kyrpZuQiKjCteU9SOsgst+7mJyawIGVFbGZyc5PMr+iUcduYRe1BiW7xiQkY42FLXuvoYyfi7dCk4IdU1goufBz+Erf7Gx6HAcOrqixZ4M0vziv97K7W5SSYtDnYsob3OxzGNQoxqsk3ftDBrGxkuN6/z5g5/tlWKT88hypDs0lG31uBgyu5uM5cGXDI4JlsOHgAjMeHwsBoRwCkoXI/6Ma0rskUHYeRHi79LA2lJqNDX9f0sAAnPB16OPMZoyFOYtoSdNpLaEgqoRYYgooDRZOsuHSYMg2Ai5sBEXYDDlrn5+Tx9M81o3NKG8/WZxE5cfL4sHQcw55af80bqQ+/U9GZEvDrP2hgDXZXCf5WbiA2/DBUHJuRgIKxJLloISWTS10GKTd7+g88f/73/SG4UZxK1DhlhjO4nOQQoBFi4qS/eBXH8KS0c8my4AKCweem5lVc3HmzBlsrN/AJK2fDhyUooJAxdziMvJT02qq2QxxQ8lPTIqdoQE8FRXyHLYw7VuBChU3vbaACrLiTj32KOIMtGIDJqDCBulUCfEa5vt3r3EqKrRlB6asF0LO+CYLWJttsEvh43gfXrx4ES+dft7yKWRvEFdGhSl7YgZUKG/GVAw+sHHWBYsb3dvh+hGiH0AFNoZ8Dh+u+GvbBmzsTRUrVJsI2CJY0Eds3GyddMyC1ZQDOW6FNBqyZZ+RjR4tFsxbnZ7pYpY0m6hXq2i36pL/f8c7P4SVAycBsn7SvOdaCqklcMB7gGqSaB9SR9UqVewWtlEobMoaq1GnLQz/r8ojnV6plfIeKuWSGnVXFfH+oBVALpvA8oFlsSbL1TouXb6q8EOyDRGh7/fNqoZ9MCB4ZsLyd8RYGbCIph2MrVP+5QWgs3n4HAYM73uNqnAJ8mT/PRVaNwWZ3jzcHx1A3jok9vfpA05Xt+wzYe1V+Hv+WB/A8vu8lzjY4cCE9wCPJQePXoBrsMkBaaSPQweX8O53vws/8pEfQ6sbwcf++b/C4499Cc16bchMUnHl65dCeIMlXpAre+ErcCWwuXWNBEWPfQ7CIgZUyNak10N5r6Bzah7tBtL5/6OF+U0DePfwD0M5ARWhABxaP4XAWwFPI6CBF5paW4dABYvYCObzM/iVf/arWDhyFJ24ZSVxytNudHDmxRfxuc9+Bms3rmFj/TpeOv2sWVjRU5xDNF1DNiSllZSYRaFhGwWd9MlfRpKu60+uf/tAjbPFdJ5VfgeQLQLUCFSU6Fdv4M7oIHg4PA/gxOhjRq9H+wARgXl8zK3XoCtvbPBNUNVUB+6Hq5EL90OxWM2fX2uJpAZdLB9cxj/4n34er3vDm9CPktkGFAt1DbT6vQ6uX72Mz/7ZJ3H5/Fn0Oi1cvHhWQzECFbxMjt15An/rIz+BlQNHUSxWlXUUJdiezeLUk0/g1z72vyOKNnoRAhXi+IZbb4APfvADOHBwGcePH8fhI0eQSjHTKMjXA0nAmz6y2q2x7KNarYlIwaEvsyoe+dxncfXaNfz5n/+5BqGjQIV80MP97c33cM0IGRRGbjD2t58ns1syNi6JD6zhnJUlL/UQlO3rvN/ntOukxwwZ4Fx/fL3xNSEq4COw/4ONmgMVznQzUcV+RoUC3akui4fhGlls8rtuasD8zQAV2nM45EiYsmMiP4F0Jo0rVy/bEGFEUeCNZihtQj1k1/V+vWLXs//v6xvrHLKsaY/D1+Ix49do4CeBCgLPwyaRdmqyOCKwRvM0sysz4wn7zLb2f61NhB9/euf7/bV/jziAsr/+RqRWtbBPs4EzsYXvAxoqBCWenzsOVlmTEazg3snjNzc/gxPHj+DEnXei1eyjXY/jK1/6Kh5//Avo9ssYDLj32PqrHB41zqwBYmCNMpqBo/tatglG/mHN6PkfZnUBDefvkn1IBvV6G1evrN4CVJiiwoEKvx51LAJQwedK02IpEsP1a6tG+AlABWsX2iBRucEagpZStHJlRsU466yNGoq7Bd1/K0vLUh3bsETpaapxGdzJ7Df++9Kly1heWlb9MJHL67kJfrRbDeSyadBhRDYSvT4Wl1aUgxBLJPGJj39CQAyZm9PTMxpccFhQbTRUw19fvaoeieQrgrK8/3nPcV2jurffa+Hbv/3NWFqYQjzKAThrdJKtxtBr91AoVlAusUZhfZmQrWm7zcyFnPoi1pQ7W9uq9bqdPk6ffl42SMxcu3Z9DatrW1IbcJCTjsdxYHkBkUgPs7MMsJ0VQWl7cwfnzl3Aq1/7MPITeQGr6UwKa+vr8pkn+DI3T9JUEnvcH3Q98HN2wfWBaoL5+UVw9sO9l+QZrYu9vixlqaQkaWc8FsVkPo3JXFbZYwMyYmNWG7ORIBzX6Ufx5DPPK5x3b6+OVMZU7wwjz+bSOHb0sMhrV86fw+GVJexubVruSjSGapOq3qTUGVSIk2DGTA2qYecXFqSMXVpeVo3crNWUx2SEsQGura4hPk41TlrMWgXWUk0l/DesySSBcT0cmLVZpVoVKEJVYr3ZEKmM5zWdjKO8s4m3PPwgThxZxvq1i5ibmhDZbnl5Sbkhl6/ewB0n7gbHSl956mk0uh38fmdea4/WrLB02B8GYobqLNhA3fy9b6Exw+23+go5AvetfxYRkjwjcWTHc5ifnVPWDWvGAwcXMTGRQSYVxxj38ZjZhCazWVm4Xr+2hmqV+U0RbG6VER/PodpqidjQ6trsgWCrLI/Hk6HvJSGjawpSuj+wRozHMD07Gyz3WkZGDbZCGnIHprnb5PDe0IwjWGhzrXWgnHUU713WJ6wzlHGUTGkwzPfjNZDXL9zjSVTlGuj7qQ3faScbFNyBDT8kDoSBMH+unsizM0K9zJkTgQn2lcoWDVaDRmYyG25lhgbrKeWSKtssEADlOpLQ+yfh0O08OTA3UgD3ICPW8rkdvPCZBP9kHcdawd8jv0crQssWC8qvYBvEY8zP7iRGBZSz7lK/arbgnpvkRArrMc15gr/H80nVshwWVJexpLT+SdbrQUGi+okAVbAi5XxLhEWBNdA6z7kE9ypZUwUbXM94eHEkTJtABZ/HLaI8x4L1HGdoAlncuov5fn3mEnLOaHWljo0rd0PtzLpHamARXM0hwLJWxZoyhgvJuK6m4T7S6Ab1DvsUI5XxOiTxTlbRPFas12TXZaCD5XxYELYcBAIJRH10cN+Qw0TYd5SNOUI08nmMAzteayr/1hUYAby5DVS8Qhbb22/jL+8IPDQzFaxp2grj29nZFSuIKCCbHhZa2iho+zM2hma7qQLt4MpB9LtdLC3MY2KC3to91Gol7OzuyDs6FkupOaKs1nwLoQKPDRCLXVMANMW4GZcUros4FwtK8SencODgQZw9f06SwTuPnxB76PrV69jdKcjbmvJ2Lp0smjkYJMDBQQ8LPMkFna3J7zib1hligabCxcXQdDIBacdEFo1Z/2igy0CbsDCzCbdxElQk8xMpp0MWCWbvpEWdMkf6sMapUAno+dCOJQyXZKNkIIQVqIGR1yMAYJZQZB5osyFLieGwQarIpoZKFg1/hArs25HwufgZJPMLXn4EI9jQcFjGhjCdHNfzcZGvVetD+xB+Np5f5ZHEYqjVq/ZcMQskNxaSDT94DNgg8nH8rBooUUnAYSMD1+OmvGHz1WgxdJcsXh4zs3564E1vHC7Izsb3TXNUrqkNOlgcSGnRtOBl/s5oATKqqFCwZiQqBhWbpjMvvYSNdYYbZrG0cgDxMYZpRyX5zk/PYHZ2GogYw5jXHdF1Kim+GaCC4Avi3Nk7eOGpL6NbKCEuRYVopQqCZKPnhZaGTRyKaPO2IYpySsJjnDWbYEZKQOP5u7xXeB9yQPzkY48HWwyGHMcwRlUFrcPI7kqQOW8FkbNhfbjDf/uxdnbt/sAYCnb3QZX/XECKsiWCt6fuJRvOGBuYRFPLtvAN1IfDNoSwz+hy2OFjFKZNNoCBMQotjJDdXVUB2WnVZGHw7e/4IFZWTiKaGFdGRaNZFqNNntSplIq60m5R9gTVUhmNZk1gBq8RFnkEJWj3xMaZGRV7xV3UqpWbgApeK7lMGlOTKQGiiUQSpUoNFy9eVsNOH2heMxwYeLEwOlQkcLvPuDVQkEGfRt7gWnLzWu1DMx4Ls35r6xgNh4SBUXTrwMufxQuZ0eH16MB6FLTg7+j4hoGqDThZFNsQ34v3W5+Lj3dgbZS16wMyZxY5g2bQ7mEsMcDy4gy+64Pvx0c+8uNIZqbwL//Vr+PTn/5TlIqFYegwn8M/KxscjfmCcmLUb9XVXRaYGlRgDqZoBbLi2ArKPspkyDbNJo9h2n4d+qCRn8nBmtFj6QNPDRBp1+WAVLB+8jBts67ZVzdo33BrqsCQ6VNRASCXSONX/7d/gcMnT6ItSxOuEVE060088+RTeOTznxVz7erVi7hw9gXbNTQIoY0bwWKTNrNJdIaRDzP8vJnjzD5g5UM/Gyhyrbf70tfV4VUYArpZlPPQ0SKNAJ6fk9Fr4dbjNLqW+HXlx0+S8aD6+1qwzG4CW9+Y/xSGobLwMhBdSgo2M2Et0Plg0xDtaWD1d37u7+I73/dBxMgU7kawV6gbG7fTwpkXTuOLj3wOu1sb6HeaOH36WbSbNbQIkA/6mF9axt/84R/DA6962BQVjRZ6UYKQSTz1pS/hN3/9XyMWgArax40CFd/zPd+NlQPLOHDgAO64406FFktmPRJGr/uA62vK1lAOY6mEJFuZ4drPPv2cVH3Xrl3D5z73ea1PbKQd4DCgYp/xf9M5EIhmgPLo+dR5DsGr/DkHvHzOUQUfiQ5+r4rcMAqGkEQigkrrJtBR5zh4Imt94P+BNWdNZ1AS6MYzVoPk7ZJSDBAlE80Vd1To1i0jyGZu31hR4UAFSRccKCu8PBHHtetXvy5Qsc8HDFCI2/PpBJnyydUiDqLxPNHmkSA0zxuHDFSKqdYIjDwZROlzBSXK1wEqqC6UCsTBxFtKcweVtG7z+UId5veI30eeU6FBSADtbgUq/B534JXrpe9JCWZVCaxIaX/k9ULg4PChRbz6VQ+i04qgXOjgTz/+aVy+/CI6BCr6Zs9pw4h9oIKfmXW1kZUMfPfXtvdLz2vL1hJYoUBTYGFxHnfccUzDgUajhSuXV1XjUk3higqvJRxgGa4V4YOz5qaigoDt6vUbZs/IummcQclN1aUEKKje1eunkho0Mz8iVephe2tLv8+MCtUqsq4doCs1p6nQ1JMMIijulQRYsQ+gsrvTbmnfZh1LyyFeyuyB6s06Dh8+qtqNqopPf/ozAiIJqFC5y3vAVAZAcW8Pxb0dnReFijfbAmalEqOF5/VrIra8+93fgXwuLVskKjnYNwiIabaxem1DivG19S2tO3t7BWQnskinxrByYFG2n1evXcfkxCRWb6xjt7CHXG4S6WwOW9sFXL2+KpYpB0bxwQCHDq6g12vh2LFDmJzI4caNVdxYXVUd+vo3vRWbN9axtbEJXkONTks9GusE1iY5BlYX9zSYIXFHWRq0CKP6VkQDDl4G6h0PLK/YOapUsb2xoePX77UxkUsJIOk0a1pbI7LSHKBNFmk2p0yVRoc9Vw8R5sJEE1jb2FA2Bmvae+85iWivi9L2NmbyeREf1jfWEU8lUSiXMZ7N6T2PJ1ICFHYLJWxu7+Luu+7G86dP49jRY8hm0vrMvGaoXNze3UW5Vtc5433DqpbrNoegvKYZuC7LGSqCaQNCy0IOExt13cN0DmCNQrCK9oMp2se2KrjnzsN47QN34cbl84gHAhQD2ZudAbb3ajh85Ch2SyW8eO6cAoh/s5C1vjLcY/tgxTcCKr5WTTG6DtpK+0pWXPx1NmH6r/vZ39p8GumxcUxmcoj3o+i0OijslNFqAtn8OMYTEUzmCRT3MLcwI/eMlWPH0OsOUC7sod4cYLdYw8ZWCXuVJuqtrjJdmp2WBrXcM5UPEGpYrr9cRwgQEKTgGJj3/sz8nPZ4hdQTGAdEnODsQlvBiC2QW99wa5d9se491pR21ZMQ6+ABX5/9sjHhbYBsta3lSvC2sOxVq7mNnGskQu5JDm7w3hahNuTcGahghFc6d7AXV82jXtgG76xtWVd7bqoTS5w84iRBfp/9KV9P1spB4WB9t80iWGOyn+FnVJ8+YrdsbH5bg6UWHKMlrw38+aXXEfhj5EHNjqQUsHnUsGYIubNS3ypA2wAbvjfuWVSHc8BOoEXKQKpZ2EcF+3P7vuWkOUnYM1Z5TJ0sSXIbMzVZr8qad0ThbiHVRibQeQ/B1TxvPE6nP2GKM37d950Wpu39ooMwdszMaonzG9aPbidttsKsSfeJhqO1WofAGjOdaFkvC/KoyKakUlIh+IaHX4tcMomrly4pe6nT66KwV5HTgsC5cao5iLxzrtlDjJZcIdOWdZGBNLQVT4XciijqtTrGRKB2YKKva5Wvr7lWoOApIJzWUwSWRNwyhwE5UgQQzAozq6zZQ+lc3FZU3FKF3/7nt/wReM1U3oraeBRbm9sKiONNUK1UhjYGXOy42PCmrzYbKBQLGE8kBSoQeT90aAHHjq0gkxlDs9VAuVTH2TNX0Gow2yIEFLHB4dEi6ilPQA5ao+h321okovKujgj8yDPgbmoa61sbYq4osCyVliS+3TKfUwIVLE7pjygktG8oMW9q3sj8O9l8XCw92IiLJT8LG2cPK9ZAK2IBknvFot4XPWrluS0fQkgFEBuzTUT+chwqcbNhSKbQbttwJI2L2cZM73oOqCT5F0u0r0aA75WLvWR8YePjBsClnkMqKh34Xjgg5uaeyqTNHofyNCH7xs5XuE8I16GPLV/f7Vi4YSr0Owy7bZBp2QLKBmmHoGw2hanMcEPjBsJza/jHQBL7eoMWOSYl5KYo9n8ANfiaVmXbJs4Nm+ew02WoIIt+CydtdehjaJ6zRI0ffMubho2vKyp8iMjNddT6yZmDAjCaLflec7Dgljn8PX4mbuqdficEu0cxMz2DQbeLMy+dkdye1k+U78cFFMSxsMyMilnMzs0IZOPnJVDBa4aqnW8GqGAweDTBQVIPq2dfwM6Vq9DVFjx8eZ0QqLCAbmMiKNBXti0WjCTrgsBC5s85aOAm5rYLLBC4AW9vb+szn3n+RdkY8frjNUCgwv5Ouyizf3K5qw8ZeL48tNiHm7y2bfO0LIB01u4NH4TbEDp4gJK95p7bupT2fSxj48Z+9aKIv89/a/8MQIXbkjmAosKRIdxup8WJIwayfWqSbdw0RcW3vf0DWF65G5HYGNL5NKp1Ag51pNJZHcfyXklNNgszFmtkPrQ7DflME5Dg89H6qVgsyuKGQdq0ISIgwpBXAZiRKDKpJObm8piemRIIKqDi0hUBNDa0SQRPSzI0TPHkrI6hf7qUE1a4DgNXxYbezwixX7Phshr6WlXXBotcP1dar25h5Y7+e5TN45uPH2/+2y24vPDzf4+qJew9GtPYbZb88f44l/WacsIGfu5DwPczBD/MNESKipnpDN71znfgJ3/qZ3DwyF34f377P+B3//1vYWNtLXiZUiocGhENWlW5mt1MAFT8fYyuA8aAzgwfY+/FMmCkEosAlT1aeTSMAT2iqFBmTfCTvRWo0NIVWFEauEutHkLT+8ZE0vlgUajBpT3e/78VqOhF+rLpT0YS+D/+6a/ixKtehQHzW9BHu9FGYbuAJx5/HE898RharTrOn3sRa9cu69rnZ+J6Sk9zK8QHGMRNOuznahRUMf3g/vtxQEmfUYHT+2HiN11PmtpaTCePTa1WUU6FX3+jIMNNxyZ8bjWV7pUaQkb5VlqBIeYSbGdi+TXK5+I6QMCbAyFXVLghEItsgZ/B0o2/ZxlIA60VP/KRj+CH/pu/iXR+Bp1uFOUS98mIgM3nnn4Sp559EtVSEc1aBadOPYNSaVvvk6HIHOB9+Ad/GG9723tRrjTRoxKUeUbRGL7yhUfwu7/5G0OgggC7JtyhA2BGxZEjhzA9M43jx08gPzEdcij28wL8vJgqLY5msy3/YBI0uBf/2Wc+o/Tei5cu4tFHH1X9QBa3Wx4S0Pbjfuu15RkVDlCxefPzYiidXY/8OdWftH30ZtRzMPwaGgVYWW/xmvFAcJVmauiN6Wz+/R6kbYpR/szk+yMZFUOgIkbhmbIGFEzIBrfTHQIVhkl+c0AFn552RRzEVmpV2WLqM4R73kIK7bPr/Q7Plt27vs4aiGIEDV/X+HgyyKdn5hBPjOt6ZKi4Dwu4NyjDRgMTA0QF/n4DoILn062fRgFmP0++v0fC0F9Wcp5rw3VPgOc+oi0rMH1eV1Twc+6r3nzt9XvewHEDKvhnkvtjPC42+sL8FB5++CGMxdJYv17EH/3BJ7CxeQX9QRn9Pi0XrUZlBWrXkl0DBFW4L/H4+L6yv4fYdc01mTWEjjGgEO07jh3VmkzFwZXL1wQOjCfHNIzn/xzoD8HvQOzRdclXj1GFHEdyPCWi1OrqDdV78oxOGmuU6xXtS1nnkMXPNZO5Mbz3UiWycaPY3NyWbRhVDFJOx+JIJuKoKmcuJUUFA5S3d3Zx4OBhVKpl2X42GhUNnTvtptQoPP5873ulMu46eY9lZWQy+KPf+331AVOT01L8KJy+S1skoNFqoVDcUb2ZyWbELOaHo2qU5/zG6lU0G1W8591vV65Tp9VQn5DO55BKjqG4W0KpVEevG8Ha2gYWl5bR63W0XszNT+HggUXte+cvXFLGGtewr371SczNLerc12pNXLpyBRMTk6ox0skEVpYXletAsCCdGdeyceniRczPzWN6ehabG5tiSzPjoUWlDvcjX9uHQbO242hgFwLkdc/0u+odaZ118p77lH2zsbbOQgS9blvBvLn0GBbmZ6SqHlD9To/vsXFUmg1EeB1NTiI2ngbG06hs7SCdnyBrSqovBmSTzZ0ZG8eVs2exMj+v57hy5Qr68QgqBFoVazEuxeLywjLOnLuo4dPs9AyuXL6M6ckJTE9Pq6clg5f7QY1K1pBnyADyKO08+tA1pixGKuqDrS9rJNV7Ue6XNV1PfbKqQ5YSV4pkIoJop4EHTh7D3ccOoFLcRH4ih9VrV7C0sozc9DwSuSmFcSv/JR7DlSuX8UunK7aPhzU1bDujfwzXt5v/8hcBEf91B+Jf502Hb7+S39s3fuff6j99XenLAioWpqaRT+UxNz2N69fXlFNx8OAhzWO4PjFbplwpyQ1hfnEOnU4f61scFMfR6cdQrNCBISNaB5VksbG4ht3srVWXh3w3Zo0SxOR9Y+l91iZRUcF7UoHOgUTEmonAqNvkiGFuG5/dI+F5LYCb6mXLzPKsALNyMlWAgQK2lxnxyghhIsoEhYbyorRX0ZbanCn4vtl/W/3JfE66RpjaNxQWxtAPuQZmf22vx9chX1BCAAAgAElEQVThUDqfp00WVaTGqh/a+oRahPuFuWEYyUOKa70eZwQx5fNwj3OShbkOMBci2MLSerzV1Ofk/qq1Kqh8zbaItqrWk/sqoXmVSHEkse47jHAtV/5BzMivzBtV9iPBi7ZZWjGTQTWV1n+zwJPyQYTXYBkeSBj6zGGgztfje+G+KQVavSY3E6kbaP8UMhm0joZzrD6E54JztmgEpz4+Obzl7n3vrik36Oqgus/qPdurjITntrb8JQNX6HTS1LWiKsOtK3nMgzK/3jL3EcunY93aRioRRafRwLu/49sxO5lHebeAbquFNuu2WAKFUgmraxvad/aqVREl+HfWFrwPeG3RItnVug58JRnuTuVIsBnT5+BsSDMTm6uIhOaWVYForXp3BMwevX7UmoZjLiLAbaDiW32Zvv3+bz0CD+Rt6EvWBxdIFmFsUoXocphHfzoySYLdx+5ewWisDJ8gI0aIXx1Hjy5jYX5ShetEfhJXrtzA7k5FxZx7B+sGDQgsJctkbY3z5uYQPkijeaNpkUbfpLXZrAYYlHZR1GCBOJYBwLdAFF8DVoa6BmkgB/zaBIJ/MxtwMbgCOq3BmHwT7XFcFLkgcxDPRZJIKDcT/j4bIW6ctAXxBV6ovHzvbDHkQIDMqyalemHoTLWIQobDkJ/PSQm4mLIMlRJTjIuysfH4e9xs+N7IhCSDiSx6Pq/JkKnkMLBCrx+CpllUk2HlYZE8b3x+s0exgGKeQw4wnNGoUOyh/ZR5Njqrv1yhtzZBFGZPWM6Eb4QCSILULE3GY8JClPmmyCzXxtinJyUH/z2BVlRk0JaJFlAMoaSy4oE3PRyGDPRmZL4BF/aENXQErph5ERi4o4oKDpfZ8LmVkDfObJZ5fuXRTTZ7PIaZ6Sn02m2ce/ElbG5uYmJyAsvLK2atFYlhdnFeGRVk0ceo/ohCnpksqKq1FiJgUz1AtcZrxIKhfOAxHAxTxpeMoz1oo7m3i5e++lXEqNKJmSUNf4+FEQsOfj6+thiqHDbxOuO5Y0ZMGKQouFQ2B2aNokCoMPRnEcfi59knn9DnZxPKZpxABdF4/p9kKCMZ/rxng8O1Z5AQ8CJIqKFLr2+2SUNgwoK3aMvCeyoRHx9mMnAwxqJI7PVQ9PHc8PXFIpbqxgbNPgjeV2rsM4HJrFW+SGCH8GPRN5pjL+ZCsADaK+ygUS2rUIjEkviOd30QswtH9XdmaPCearXrGsiwMCQL1n3e+Z7Y9DOHgsMMZlHQ0oZs/lKBnsslVKsFMSGpyuCaY7JPUyHlcnFMTU1iempWORgcsnQ6IZwqrFkaGAdZsjH2LUdAA/cAQpgUNhIGlQZOqajV5zTmENcbSZapyAlBsMb8oI83w9OYYWIsbQ3wR6yghBOFwnY4+xsBNlgA8TF+TkYHz/53v2/UM4QgOT93o4DFqHLCB35c880CzELA+dJtquESEUyks3jNXffg7//dn8Nr3/g6nL58Af/0Y/8nzr10BpW9gsI1bSAXVe4IATt/PT9+w2tSRWhPa5MAI5i6h6A62ccEj82ixo4r7XyqxT0VfLRY0boagIx9C4V95qIPhA2Q2wfovNA2OfPNYIANhu3LGxs/lhpKah0kyyiBn/9HH8U73v0+gWyNegf1SgXra9fw5JOP4cXTz0hx99iXv4RajQNtY1FpkK9CPvjsKq/CBrHahz37xUQk+p6Gx0FB5e+d7NAo1xup5/Y/BxssFetsniRFpj9rQ6HzGlJzLwxyYwOBAvDmwKP72fv1Hh7rjd8wTC5cj8M1QUG9ZhHnVoW3gqK3Ammy06HChakU0QG+/dvegv/2v/v7WFo+gkEsjbWNHT1naa+E555+BpcvnkOzUUG5vIMnnvgydnd3ZNlBxQivs+/+7u/F+7/7+9CjFROVngIwUvi93/ltfPoPfl+ZFr0Ir82bgYr3v/+7cOwOWj6lcOeJuzA3v2TMtWD5RYCFayQHpZHANuY+xGNd2Sup5vjyV76CYqmCl156CU8//Yxdr62mMdvEoA/g2Mifw3MZwDFveOTjHLyReTZdccNz4NeBW3353unXl1+7SllgflQAE/h+tWeEpjzKQPe42R366zmA6oqKMFpWLcbzwL2DSkqpXIP/MoEKHn+Cy4p6IHkjvAn73PYPkVF4QbOW6/M5+kjnsjh+192oNmu4cPY8BqzH2KAKL7QQQu4JrDS85uJ+eRNwMaI4EvEk3CdUg87MzA/Dsvk7rLWc5d9XiL0pZW1vpp9wyOHggIG9ZQBWSazhcIONsPbFjlkQiBEazqcDjQ4g6Tl5z3OtVtg6RLKgdaUGFyK3cB9O6HOqJR9Rxnm9YOuvXa8KXKcCZSyJ8VRK9WwqnUR+MoOHHnoNJnNzuHT2Bj75J59GoXADiNa0iPC5dK9FQmg4refCvS8GZAAo/fPaMSLAnUQ+T9UL1W5mf3jHncdwYOWw1i+SPS5dvmh1CcO0x5nJRqarqTNHASX7O8+jDT843Cfr/cYaSQjGrKTqmvV6s1VXXc2BjnK6xphpkVX2WK7J2n1Mg4DC1o5qLwIdAtxIIGq1iIZoUMz1kaHLM7PzIrrwNUqlIjLpFMrVEmanp5BOJ2Ujcu7CBTzwqlchPzmpDJCP//EfK3R6YX5B9mS2QLMfiGG3WFA+1tT0pKzlrFcw0KvX6WBt9SparSre8553ys5obX0VR48elu0Ua5pMJo/V1U202lQnd3WcWYcT7F5YmMHS4qzu071iSfVTtdrAs88+h6XlA1IFUAH6wosviVih2jAGHFhZUu20uDiHhcU57OxsyQbp0IGDUvau3lhDrdqQFVpsLIGtwq4AElrU8b7hte3kKvaEYg7T2i2wXglOsjanomJleQWF3V3sbGxoTaXaOJcZx9zctMhb3TaBgHHldQwScZQaDeRnZpSxwSVge2sHOR5T9UQx3gSmouXxrTeQGACVUglbO1tSxRUqFUzOzqJab6Dd6mF+dgFXr16X1dL83BzW19YwNTmpMO2d7R3dY812FwQN682W7FGU6yL+GfdDy6STxVnIodLaG1RzrMHF2A5rVr/TQ3I8gUSkj3ZlD6979UkcO7CA7Y2ryGZTIr8trxxAenIasWwep589he1iEUfuOIaJ2Vn8vU+eDcNEHynu1xg32z/d2rm74uIvAixu/b3b//7rfAQeKn4RaeZjIop0IoeVhVkUi2XUa23Mzc3i4MqCyCEc646nWNeMITMzo0y/zbUtVKod5VOsrhfRYIj1gOqiroAKkkJox9bvDZAaT2Iin0exUBQITCWSSJ8h22VialJh2iSUMQeIYIF8/YNKgefIlG6psNfu5xn4HaK5iCywR4bjHRuAu4pAdYaUAD0NrNmz8efcV/h97kmuajegIcw7pKIyRbPvvV5rm/209azaO2NmzTxJoFfrB/e/1rBX8b2On0nWRSNEMSOEWa/C96EajKqNpM00hvuvnD4CQBM3RYarP1ifKBMkzEykIOQMKDgiaN8bCc22oXhQsLCPjcbQIpFUtkSmUtF8iADFsLe0zE23Vt//M6ilw9yQj+dn8hqVsyauYyIrBuCHazvnXyIrBdKT3h/rM+3VRsbluX3+kzPD25WKCu6j/GxunbR/LxshhfWSE105byBIYkST/XXS+zrLQuG+TftzKj3o7DCQswtoU95s4L3vfDsmshlsrK4qG0nKCYbR94Er3Gd4jbCuYa4Y69LEGBoKGO/qmnain9ncGsGD70Rz0XB+RWINqhTNSlWPmWUW60O3eledFb7v5COVHlKOhhnEbaDir/Py/lf3sxOoYCPJ4n9mZk4LrLEfrRjl38kCqVXJ/mXQWB1s5KKDuKRGQip7LUQjVAn0QQXV4uIkDh08gHqDGRYNDfmFFtK3LvjF7u2VsblVQCTCxnsM48mMNj4CAONjDOQh53EAop0c5ip/gc0UF6puT42YQh+ZB8CBfAhj4uJNVpz5041rRsVmw70DtSmFXAd+Plre0FtQCDQH+PT8Tya1iDLkWgtnwqyQhDZzs2lxIE+vYg58LeRbQ+V4QrYJsk2RN15XTRMHytw85F2YTMmbkQ3c5tamjunUxASilPFJGUKlCF+vJokYWU4aKDVb2CvuyW5KOQQ9y/TwzAYx98MgScF9BG4SFnqtnA0y2fo9gUA8D/q/yxBu2ii1la8ha4nAPOPCR7ZYo8FmhUHTZAmwGSDDjR618SEyzpVXiyqvASLe/Z4NYsR14jmnHVZLigoOZx988+tMBheh9RELEWPS8WR1uq3hRsMG04ctYn/eAlR4ASCgglYWlO7zvcWimJ6elHf++RdfwsbmJvKTE2qieExoDTO/uCCgYo75JwGomJ6d1iBbQEXE/DarNcsQ8IGzs2C1QbBwGIuiPeiiU93DuaeewoDS8AgLDAcqTNrJ4T+zT5TVItZqRECFKypcBUEQgwx+L1j8dQlUsBh68rGvGErPTS8xhiRZfglr3JPpJDo9kxPG6R8+Ah6Mp1N6TW5wlOUmogzDDIOYAbNcOCAfE5jBQSuH7z5gabUoQbW1wAeKYinEqcgJjMoR/21eR2KhDEwBxH83anX1XQrGFDg30HCBUn9aO9G6rbizhQqDU3ldJrN4+3u+G5PTBxCNJaWc6nSaGnwpRD7IZXlMlF8iK6WmwAoHKmqVsmyfaAvEwGAGbVfKVfkxCxxVURzRYCQ/MYbJyXwAKsqyraCPsQFx+yx6Lxx1bHiseD7JwA2Fgg8L+f54jAQUBhayijfeK8ELta/rRLxgkyFHA4OZCo4xs12xQsQGSvoKGLHeVhA5jBKV/XEOzt46EPIhlx8/Z/0a8GIMFAekfDjl+4CeKxRFtOjRwIl3OAeU/Q7yyQyOzi3gb334h/ChH/gb6KcT+OWP/Ut8/nOfR4mDha4xeDlQ6ZO5ewtQ4cfOhtiWwWPvwdRcLI7HGWia4O8K9ghZMDH54df2yiaPFYJj52x0UK/Ddwv48PWACv6eHzsDve2e9S/egzy/GkaGb4pbJRBlgH/wD/8RvvMDH0K3F0Wr0UOpsCsFxdmXTuPK5QtiuH7p0UfQaFZG5N4+zA8scOwDOXw/DgBqKE1P7QDS+5/+PnkdcS+SzdxIgyKwKVxDslVSgL0BFTeBNcrXCex6l2OzFghBez6AHRb8I4x1X7d07HhN65piKPF+FoBfg36MR69JNRXeyFFhSc5ev4u7ThzDRz/6izh6x91ANINCifsSsyqKeOHUaazfWEW9VsD29hoee/yL2N7eQorKwnpVdlLveOd78P0f/mEkUlm06l0BFQR2f+ff/t945JOfFIj2ckAFFRWHDh9QTXDsjjuxtHIQmXRW16cG/CEEj0BwlFlBJEVwr2q2UC1X1PAxW+jU8y/ghRdewunTp3UP8Nrx8xYbUQH4sfV7zq85V1KMAhWk2UvBIoER/XCtQdT6G9ZHZ9/7cbVL1RR+YsPRzjEAFcPrK5pAJG4WCm594Gv/rUAFlYeW0UVbT7N1UFwuQZB2R3UjrSMZJsT6wNeqW4EKNda8XkItwfX+0NGj4J58/vwllHf3EBHITg5nGKDL7pDv1QBgy0+4+Wv0GvW1m3XhxOS0mPj84nHgANLVZzzmfE4Os00ZZNZtGlQEYMCtuiS3D+CM7jUeAWeA2oIzBANYE4bDbyCRiB0qJNAhk2/AvdvWYRrl+7kmgDMKVPg9rfMnIollmGlon86KtUiCCxn9Y8koHrjvHhw+eCeunF/DJz/+Z9jZvo5+pGrWakPVhgEV/r+gAwEVFvzt+76GAcqnSCKbdfWOeTbfeecxLC4cuAmoYCilWUQRhPfa04CKUcDcwA4D2KWSSIwrL0FABTOqxhKWq9aqSWFByxBXD42PZ5TPMYOMkSfSWdSLJSSTaZw/d9aGUc0GpqenNIwn65F/MiQ7ncnq3rYBtNkikslLeynW77xWaLP00OseVgAsCSu/9f/+O73HpaWlYQac7J1azJcooFTmcC6rx7OuJdAej8bRbjWxsbaKdruOd73r7YjFyPRtYIzWT7JQ4hqfxMWLV4BIAt12yFsR+XOA+blpHDy4rPrp4sVLuoZpX3bm7DlMTc6gVKkKqJJVBC1X6JstZjF7qhjuvPOohEJcEydyOQ0V2z3g4plz6HIx7UeRSLOvsrwWJ01NM4i6RNCV72PfXzudzgrcIagp5U2vj6NHj6G4sy2V/JjYxG0kYgNM5LOIRnn/s+8gESmKCEkwgz5SE8yiyaFWqeHatVXMTM8aaajR0P1D0KtZbSBDdUqHa0oFlUoZ1WYTu+USphcW0Wp3MTExhfJeGcViRTU+B6DrN25gemoKkxMTIfMwIdULPb74WVijEuRgxayhUrDhlFUX69eQ9Wa2MHH1ygo6ZS4QVe+1GhKxKFLsA8pFvP419+LYwXk0qkUpP7Z3dkAS0N0PvhrtQQSPP/44VtfWMTk9gzvuOoFfeGI75E+MrlujoMVtIOJrFvX/xG/8l9NxeAj6K+/cvan2OCbTWSzNziFP5R1iKO1VUK7UFKadSY1jb3cHW+sFUkSwciiHex+8X2tYoVBCqxNDudqWBVS7G0GpVkeLeVftpvYgkg4IzMoSSDbZNlNhX825AIEKzg7yk3lMTk0FBrnt2yTJ8rF8nMAEzXQIPFtos+rCW5TE2hedaW5CdwNE5Mxgg38jo3GeZb0X91jLerAcAA6U+eXuDuqfSVYN9qhSSWpgHDOXC+YWjgRqc40olUuysvK6jeuF9wi27xnIwNezTEfLqLC6zEBHfkYnJvI5uSdZ5paRjbju8PucybC+pPKD85h8Pj+sXZQPEYAKzrr4ntyVwp+fsx5lpQaVBWsR5s/ye8xoIhjN73HPUlhzyDozyywjwnntan2D1QhSmGvWEbfsiXGzGW+RwKua3hQP3mPaEJ/ZGKaK8X/zGDhg9NJnLMOHX/d9ZyEcX3t9HjORU4K6lsfYCHp0JDEAylxb6GbCeQ4dUZitaYCYgJdWA7PTE3I34Jyt1ahhaXEeE7mM1IF0d5ikRRlncI0GJuYW0I8lsbq+iQ5zZDs9kZC497LnYh0yNTtjVqIdyxXh+ZKThgBwqwmllhFAZUHuBCpULtK6XgCGAVY+x2Pvq88XMmfVRfPvstEy4MZ08rcVFf+J28PtX3slH4H7smnJitlQZ3N5G0ZykaICoNtVQ81NxnzSOMEYoMFcidi4VBBs1DinoxdpLEo7mTgOHzqgxZPSvq2tDRXKbIq4QHERY3FNJhCzLK5eX0epykU3h2h8XE1Ns072eBX06q8HXz3uMoNOTyiv7FqyGbSJetJXLniJUvnAzYEbCVUO+h2CGJSgxRiSTdlVB5VyRQN5IZEazMbE0ibAwYWFzQUXcbIiDQUls9UG8JQPkxnFDYCqEA7k5TNo+ivZ6AjJTlrgMd8rFxT62XKh5PHkYkkQYjyZUJifbLe2t7FdLNjiGjaQ4bDaLVq4IVDG2Kb1E5sDCzvP53Iaghf3irbx9wdIZ9OolMpq3LhI07OXeRFsKOkfzHNLmxGBAwz8oWVFo6HjKsZaLCZvXm5c6+vbSCZ5XGL6jNyAeHw1BBAD36SGfE/1GlU0psSgVz9VFbRIEoNTQEUXD7z5YbOS4ZBYDGkOxhyoIIOallHWJNxk/cT3zRCncaoUrHnme3CgQmyGBD22I5idmcKg08X5l85gY2NDQAUby7E4ByoJzC99A6CiyqKLypR9oEL+xsFaxwc6BCr6caDD8ovMz2eeQadcMhZwzDYh86C0ITQtDQSeyUfQGKu8Jp2RrKZIvuBkUtrrOVBhgdBNPPPEV1U4EJgy6yeqKQxgInPR5K8RgXpiDIhdHkUykxZQpUKJj6etU7Be4rXLZpmvywaOQ0Veg86W5EZrBZNJ/7mB8ljbUIFFmL3maJHF64KsAwcq6FvM9yPFlq6ZGMaYi0H7jVRGlm/lvV3UyiUBhMlUHu98z4eQzs0hGk9iECcLo6n7j8eIwwoeBypgeM8YG4ZWA2YPQUVFlc1suYRSsWjKitKO2HkM5HaggudGg6uJcQEVkxMsMsq4du2G7BycjW/1xc2MerH5Q7CkW3V5seWyVgfaCL7oPRJEFBhpg/hRoMJtNzQMGDPJrDOmR4EKso+/HlDhe83LKSo0qB4ZEI0qJvRJQ8CaF/dfO0yygl2EE34erXURncdmp4FxAoDpHN7y8Ovxkz/zUzh2/0n81u//MX7zN/4titvrOjcs0L8eUDEKspiFkAfjmn+0hgdhcJggkDMWV5aP7w31clWsbG1I7nk6oijwz+h/+vF4OUWFgzVqjrj4S1K0f/55X8rzdqhTo7Ueg+bp8drFz/zcf4/v+4EfRKPVR7Pew87WJp4/9SyuXr2E7c01ARWPfuGzaLX3gQrJpMfHhyAlh1U8z94MmPo3ZHr07D70AbIX/1qH6S9L0HxEAXUT05zPE1jMDlT48/o1bkDciE2XFrF95ZAfQ10jAbDi9/y68+vQ2MyU0hvQMhx4h7Xbr7FRZYpLuSWbp0XToIvJySx+8Rf/Vzz46ocQjedRJ+O43cfGxiYuX7io5rpU3MK1a+fxxS9/AcXCrnxx69WyZPNve8e78OEf+hGMpXNoN3oKMqWdzG/8+q/hiS984esCFQzTPnL0kOqhpQMrOHT4mKwhue4KqKI6jdkAXMcFwlorzXWKmSR8D1evXsVXHv8qnnvuNM6ePaO6gjWXX1sEKvYBRWum/d+yqAz3JR8vxVVovtXwqGGxJkfWBSOAFr83yoQfriECKqiANHsmARVi0ZmHP+9PqhUcqBCg5ICp7sDQEHE4HuN1ZmAUrw/J3oOagGx2AhUcmFosJ0OF7cp4OaBCrGX1n5bPMjUzg3sffICzSWUzcQ3VokzFpoAzElWorLCQce5Rt375sfFagf/m4IBSfWYb8Hrkfex1hu5n3h9UbCj03cBsCsEss4x1zL5NE8+/mJdh0CD3/bDG7oMkpn5is6qhRJimKA+Nm+SAAxw7PrSgUaDmEAAiEcjWWgedBFQqmNOACjXtXJ5oJZnOimlPgko2l0U0NsCRwwfx6gcewub1Iv74Dz+O66vnEY+zxnEwl4Mlq7/MvtBCwaW/0rW5f1wFbLCWSSZlvWTZZz2pEY/dcQzTU3NfA1RYDpcpKowkY59l/5q31xBQodwugtH7QIUCUpl7UW8oh4p7P+sdqh9kd5VImh1ksaOBPdUOrFFZY5PYQPUvB8r8vWbLhuSlcgWNZkuEJ9ZM2WzGLH36PeQnstjcWNfzc5jGWpfBzAR/8jOzePHU83jqyafU4zC8mfVzejylQf/29ia2tjewvLJswyfWUyABIYFGvYatjQ30ek284x1vQyTSRSrNGp5EsQTKZYIrGWxu7mIskZayk5cKr7lyeQ/3nDyB9Hhc7+n69RvI5XMCWj7/hUexuLiMbG4Cm1vbuqY4MJESvV6T5VO/38bRIwcVdM7alOs/h4qFnSIKxbIURDdubAu8ufu+u9ComwWSKYOC1S3r8oFZ+PG629jYUn4PVS7ZTE5EormZGeRzWVw4cxbx6ECkMypHlpYW0GP2YZzDuDiqDdoDn8XhO+9EMpdFJpuTMqtWrqm24B7OtbNcr6LTYnbRQH3XVD6Pa1euChDiPdqgypsKDa7gPZLTUijslWVHQxIWCWxUVMxOT2P1xg2dK0KLHKS1FKANKZGoeWWf657rIiSR8RvAfbJteV3KXjIWQ5Pe8ONJyz6JRQRUtEq7eONDD2BlfgLr1y8jk0lKVcP3N7O8gkFyHLubO9hjdlqtiu4A+JVzbs/yyhtqv5LnFq/s93arKuaV825ftf05pONUVESQT+dx/NgdqFXqKptP3n2XZjURAmwbayjXK8qfyOcnUCiWcOXqDmqNrgCKTG4SkUQKlXpDqicOo7k+tkn2DJbE1sfTnrOhNYwZZnTUYJj2wtKi7IY1aA0KO5Eow75gjg4GcojhT7eMMNgX81/KQxIbaRG0X/9wnbXB+f79JAeLbkd7oika9u1m/XGuSrBagKTb4MIxYj3lJNhsmjlp+/ZJJFm4st/qi7Eh2ZL7nLtcsP7lcSIIT1KlgZ+0nLN6husLv8+6zBW03F81eCdTnwNv2XFavSMLc+7HgRzL/VhZIL0+Mrms1Fzeh3r/KrJFUHVQoS7CBJUMdCwQsGPHknVhr9PTfELngvO/8DPvNfha7MVVA4RQbc2CohFUCegGlTb7EKrzOLPQWTGWqvXtQUUhNTdlpAKHTcHH53n+k7PDm4eKCtluhRqXcwvWrpofBesk9uMEcUS8k2KDTguWp2mkDCOdqa7hGt/vIJtMgBZl6bRZr5+8+zgOrCxjwLwiqv6KBRR3d6W4KFbqiCXzaPfYe8VQqTdx4dJlI8yEbKcjR4/qNVTnKE/F1BWskwXwhMBtfUaRzsIsTQCKut7QAxr5RqTDQAz0Hspck+1ccXYi2yr2Azy0t62fXjkL7u138pdzBE7IO9YGv1zgNPgTa96+Z150ccmt+DWeGkMqk0I6mRFowMeyMY0OesqxyKSiWFlZRC6XRmG3iNm5vG6iKG84AhrdrgbLkt7FxsSM3CpUsLFdRIMMIjF22PASsWc2BKVb1jAR/SfyKPsVMWqtmfKAWCLBzgyWXVPwFjfwxRQQ2uAkzbdiwps+NQRB1u5NFJsYNeUaDHJzhCHzvb4UCGADEiP7yCSFOlYJghxjCjNiE8Xmh+E6PVpdRUwSyAVSqK40/SZ7p284ZWSyHAmBi8ri4AZBvg+HTkRow6BXm/agJ+CBw2C+PjcqAijcyAg4kE3Op280GbSU0gZANQwbGQ6z1Mgpk6E19KonA5yADRlhBBx4nLnZsdm04M2OFfTcMGV3QLsQA7TIQGMjogByevx12mh3mvK5ZDNrxYopKhyo8EG+N8oENUYzKngunDFP1jQBM7dQ8AG5rt+ehUVFWGjFIpifm8Gg3ZHtzNbmFvJTE1haXLIhQCyBOSoqpmcwtzAn2Uh+kXIAACAASURBVDaPy1BRIaCCCDxQq5tsUl6aIS+Ff1cDw0FBzICKSKeBK6dOobazbUBF3KSSbJy08dOvPEHrmiSiCQIBNgjivWA/N5sgt34SUz8M//knzwk/34unnsPOzo7AOLLYGPTHzyQf59SYjr1YtQGoMHkjBFRQosvjOcYwxKgFbxvrOSoGPwcQbP7og8WN13IBgjomFFM+fPEMA1e9jL5XG+zeDFRQOmwDGhuSMssklhxXOGUqk5f8slopoV4uoV6tI5Obxtvf/UGkMjNAbAyU6rRaVBnV1JzzvbFQ4nrl/qBUYZERUa9XQDUFMyrov7+3W8BeYRdlWj9Vql9j/cRicWoqpQZ7YoKqmiquXFnFoB/YIrcstaNDXRZv+j8MxEcHriqMQrFG2SjvY7KEOMSU5DXYiLhHuCs8VF0x7DcMrUcVHXZcbTDlQz+3UBl9m6OD9tGiXYVNaAZGgQgfgo2GbVtNuc981fOIXcTZmg2bBBRm6VVLT9MOppNpHFs6gB/98R/FO97/nXj23CX8k3/yS9hYvYJGLQzlNRaOacjoIIG/lg/fJUGWXb5lfyjsNQTgcV3RYCvcR1qf2z3USgyINUtBDht9fb8VYPLv+/Gy4dstCorA0rE//MncPM9+cwgUuMVLYPdwzf7+H/xh/MiP/gQqtRYqpQbWrl/HS8+fki0Ir/N4NCKgotkuDf3pHfhzwK83sHXG97TR92t2NDakHmU3qZFJjIccnBC+Nurjz/caMBcDvZsa6o9e096IeCHsx49DaH/c6Pny64DfG1VUGIOLe+TY0Puev6+mLigBnMXuMmcHj/zY8hogASI5HsXP/uzP4b3fZWtCrUVboQ7WbqzJE71W2sNuYQNnX3oOj37pc2o86HdMoIIN13u/6wP4Gz/wg0A8KeunVp8ssjj+r3/+MTz32Fe+IVBBaxZeUzNzszh67DimJqeQov1eq6WGjms6rZ/YsOtcRSzTi0gtGbinT5/C1nYRjz3+GC5cuKCmgw2r9hWqipxVF2yGBC6EuoBNvV+f/NMDGnW9mphiCA75fe7NzOi97gw1fwz3YfPWN1UFv0/gWtcTg+TjHBhb5sbol9ELTJkj4gnPLc9zNGGj9gDWaa+U9ROBZLN9VP7HLUCFHieve/5sgFiwfiKrO5XL4XVvfAPuvusB/M6/+21UikVEHKjgIkTyiOT+PO7cL29eqEevVbOAtwdwjctm82Le+9Dc1z8NStQtG+A3ZAz2Pe+C52YUqKAK1lQkdi/6z4LSKnxeJ7KEhUPHQco62qFSsRDkJK6qi0bsXOg8jwAVxiS0NdyBCtZWZjbJYOAU0rm8BgysBXn/TE3m8ZY3MjS5iD/9o09gfeMiEGENZ0Md1ZTc+4NiWeR6ZcqZ/7Pdi6au4J9SQFO1keJ9zfcI2YbQ+imTzmuYTbD24qULqgdHgYpR66f9IZGpbg2oMOsn2gOtyfrJwrSTVGU2zdpRFpkM006ngvXkmBj5mQaJG2Yvxefw9XRjYz0oexrKvuALkaxDpQ+z79rtDnL5rAY19z9wP7IT9KQmWBBHfnpadS0fI2V5rabQV9bA6n103CK656nuKhYKqNYqmJyaEPFLwHrPwu5Ze+zubqHf6+Dtb38rxhL0Ry8LxKGVIa+HdCaP8+cuIRYdR6GwhzlmMgx6KBZ3cZRZORM5DQRXr68im8tJHXLp8lVMTc1oj+R7o8rJzlkUpb0C5udnpDa95+47paxIjAdgLxZDZbeMPVpdXlvF4tIB9VwKve1baCyf7+qVVZy85y4RpNj3rK2t4cjRI7p3SGS6vnpdn29+dlbHiqp4et2PJ2L6k/ZTBw+uKEOItSrX41KthsLeHg4eO4q9ag0zM7O2TyhIvofVG6s4dOSwyo1mqy3bXPZALz7/gpQxVBhzbdzd20MynUEqk0W5XMXS4jJeOnMOyUxWdq9Xr1zB7MyM+lmuybx9KjWyu6mmz6JcqxmIHiWIZcxf9WZKVd8nA/D7CtlmRgXV7wRT5MM/wDjVV/02urU9vPHhB3F4aQa7mzeQyaQU2H7sxAnEUynlYjz59NO4cm0d9z1wEoeP34m/9+lLtiQMdZnDXX5Igbil/PwL/vlfTjfwH/e+bj/6lXAE3lj+CpIkqvUjUihNT0zJ9k2ctj5w4o6DGIvxWo9hnHOeXB6T8/OoVetYW13H5lYZhVIDrU4U9VYPtVZbCizaPmmQTTtdRJCh1TTzbLq2T3Hew72aZLlmp40jx47KopD7vjIMRokrsmi0gbfv18ob8/szOAXwZyILBftaU2QTbDZrS6kxRG4ykiz3NK5fnIX43EfEPZHtbDBuZA8LYDZLausLfN81tZqT8uz73uexH3U7JssQtefz2QnfgxQZwc6Kz8senI9xQMNmDMact5lbICYFYqYpLwws9nrbLczNLsrzR2NywOBMaJilE4bnNtC2Xs7JSHwts8608yeVQzdYQyrTgzOdoPAfrldGVLW+zM1AbV7GzyRAm2BTAJnc6tJrJNaWUpUMzD7VhvokM5oqgs996k+nhrfNPe+m+sxej196/pH8QRGmwvvRSC0oOPhYvg+dt1EFCJUMzGCZzOKee06iUNhFsVjA1ERepNtLF85jbm5GNwZtBHlOr61tYn2nhEq1rj2gJ5vLtmytOLvMUt2iur+mY7+8vCwCZZVEiWTKzoUAk30SGI+9jQKttjPrJ/vY2ouCjfuwzwpkcv5cvZn2+mBhLBLs4utuw96vhNX29nv4SzsCdzNcOXjHcYHK5fPY3dlRg03EVSxoWdHEFRAXSxBp7piMmyzXtsnXedulUxyaE7xgOGEHly+v4XUP340Di4saGGQz4+hps+GG0TRkMUJWDFCsNrBXqWNjexf1WkuFJiW5cXq0cjjNYXSH7MpgeRILstwgR5OnXlBPCDV3O6KAwhtDlMPzTmDNWFChGm7rwsxKKQQHufxwOOQa0HvcNmBaRZFV+fBDD4ul84UvfllSsUq1qsWJ7CQWs8ysUEZFsMhTo+yLuqypTDFAdjmZwVx0O27pFNjwsgSiJDJGVUYaSwsLGjKvrq6i2WlicmpSw4RRmwYfbGlwH4moQGdTx82gUq9aaHezje2tbTU6bEj4OJ5nNuFc1CmdE5ovxNukkraQBuaiwsp5Lk3CpowLZoIo3yQmcKTVbiiMm97UBCnYLNHa6YFg/cSdiMN2HiJr+KJq2GwQSd9Fk2aajLODLj0xg8KGP3f2ujy5CWwRXedwMx6VjJXSvbMvvChv2onpSSwuLFpTHk9gdn4e2elpzBOoiNGZvK8wZTagBk6Q6UDbMzIfWMyQRWYAkzNamaVA25sOOoh2W9i9cgUbl9l4kGluG66HrNPjmvYAAiLI1iSwEIAKHxybJ/iY/HN5/dg5MZ96t6a4ePaMGLoEKuTRzGsjMLHjDHyHbfoywxhptCjtlKKC71/kaAOgeO2LnS4GKS2fOFyk/RSBLzJQOjZoCmqMW4fexgjZL2iGA0/ZZJjVE98/FRUCKXS/8X+GjnPYkEEmN6UGt1rZ08CxUWthZnYJ3/aO9yGdnUE0kUR0LIK9vV2tG5OT07reeL4dwOG5oTUUgQr6PdN2haoKNuo7m1vY3dlCvV6SmoKqChasvNfFQI6RpUgri4wCMgk8Xr58/WuACv9sPkQVgMDifIRp78XFrcNx+kXzfPGcEGgixMp7jXZyfu17GLeGTvTKDOdehU0AQgRwqEIxGbTei7DO/aZ6dHMYPV/+dy8shy1xUFp4weyDUR/eaygW7Ec0t5fDkTHpfXiayFCpVUMuNoblyWl88EMfxA/92EdQG0Tx0Y/+As69dArlIqW7/Nz8DAZU+O/78M0bgoBoBRY+d5eQmcCAVLLBaXlCezUpuWLaGxh4pqJNzPCbt0g/H86wHj2Xt4Il/rkFGIzmj3ydQahJnsnpNBCO5+/+Vz2Ev/1Tfwd75Roa9RbWr18XS5esWtqT8X0+8vk/R7P1tUCFDyh7BAw56A92cTze/qVCPnjz+mcTQCm28TgioyHuN0njbb0WGYDrarupkHkHR7hH+XB8/xq2wtl0PPsFtF9HOpayBbk562PI/qER3UjeBo+XH2OF34V1yq8BewXLmNJ7paVgrI/v/d7vxY//5E8hlZlCm4GOxTo21zdR3C2gWa1ga/sGHn/sETz2+KNqCHOZLJrB+ul9H/gQvuf7Pox+JC5FRY+qrmQC/+Kf/TKef/KJbwBUvB9HCFREY5iYmsLho3cohDZL9mC7LRYxmescrNLKxJhcBlTsbG7j3NmzZqOSSOFTn/qkgApXVFjjFBOJQ+tGCKHeb/psL3PAiI/xNUHnKwDC1qyY/ROVR7JGk0TcyCdcu/3+tTWAHsYdvQ8pMEO439BqKKgj2MD7ORwOlUPjZLJ1EkfYkJsKtUurNiu8bE/o9vTZ+T9rgAHlElJS2hfNI6UMGFWIqX8eoBcZCFx/8LUP4W3f8T784X/4PVw486JCPul07T5RgghusXjze9tBM62Vwfvar9lUKovcBIMaDTjzYYTuZcnnb1ZUqLCws3QTUGHJhwYaqvEfWSNuWnvDmu0DAllW8Nxw4ClgxAgDbodH4McXMa0pgXnq66PXP6zFjUhj6w6b5dzk1DDoWgocDPDWN74VVy9t4POf/Rwq1U0MwNBwsyOwa9ZACw/VVvCpAJDhu7C7kvdNYjzUmzbwJgt3YWFBQEUizvwW1tkvD1SMKirs+WyYw2MgC2iqmxWQncSNG2sCPHgNDoGKkYwKDsl1jVJRkcpg+8UbGmizN2G9xFqdxziby2ggpGHawHy2eRtcu3ZdA3LW0Pfdf7/ATdpnst5hXUSggkopEo7UJ9AGI4DDUkbSL5rMU9XZUd3bFy6cF1CRSSexuLyMer2FWMRCUGU7WdxVbfiG178W0QEZm7SqGpfVLWtsghsMtsaA1h+Wc0fVdjJFz/cMpiZy6tFOn35exJut7V0U9/YwTaACrPXNgsJYvD3tN5k0FW193H/vCSQSUbSaZl/EQeHq6jpqdQ4ReS9CQ0SRaYI3O8lavAIIynhNSiDBBnAp3Ye0fSEwRAVKu1FHh4SmVpOsNFkCM2Po4MoyOu2G1ol6pYFqo4kLly+DY0QGa8/MzWNmcgpLC8tSnd5YZ7j3hMAjrru8FthbFXYLyp9jr8VzzzyO+fkFMbm577Muvnp9TV7h9Iy/dOkSlpYWZQPGHBpel7R+kno1Pobdwt4wF0rBsrzPFGprNifKw5EVm9VXdq1yXU6YZTL98Glt3GliPNLFg/fcgfvuPoYr58/o/TIMfHp+HksHD6IzGAioIIltZeUAqC39+S9v3lyo/Gf/6zZQ8Z99CP8KP8EbSl/CzMQUpjI55JIZZLhubu/KXYGr/9wMyR17qlFpv1hrdfCah18ra7XtrQJKlRZqjQGqDdrecKmPyc6p1qyJEc/7m6AtHR6cnMa9t1Qpa9bA2pK2m3ccv1NqNnfBMOcJG4g7UdPvNfZnvBdlMcmgZdb+mkvZ3IPrX35iQjUX171A2NefbuWn2UYA91k7W6j0fv9ihBnLD+UmZyx2u9f5ugr2dpV2CME2sMMePzo81xwiWCE7iYj/Zp1hYAKtio1QqNeRksB2cFMkc53hjC1YRQYShCs/TVVhsxH2saw/STDlv7l2ez9OJaBIncHlw9QItt9KPRvIJuypjQDHUGfLyLIcQlN8mq25WWqr7wuwqu/dUpczk4PgFNfIkL817GOCzSX3HL6uXSdRDe1d4eHH1lUGXhucHs2oeO+uZRB2LQ/V7FAti1WgT7AKHx3Syx2GdXkAW3hOSe4VQMLjgy4mM0kcPnxIe/f01KTZBxNAGx8TYbfIvLtxqqVj2NwuYK/SkKJOQHWMKplgvUm3DCqI6g1MTORtVkW7z4Hl7XKeQvd77VUixnnNbtcz54BOAuIx53mUzaD6A5KU4gJFCJ4px0x5iCQz0zHGAA7NJG4DFX+FV/C/ph9tgTZOYVDNxZsL3ezMLHZ2d+VVx7WZm44zzlJp85M3yyTaKWXkSUi2Tatex0Q+h36P3oJAuVxApVjGa199P7JpAg1tdJpV3VTZTEoACb3w6+0Oqs02Gm3zfLt8dRfVegutblc5Agw9k7yLkj0u2mEwYgy+nmRxXOhYTBtCb4N33rf8PHxvXMxYxMqqRGHG1lHKRy4MurlwcjPIZLJ6LH3m+EW2OjcXFuKUsPExC3ML2N0hAkuPVhsmk/FlwWyUFxsbTUh+CIumTQI3q2a9rpwKKh7SqaSekwNs47DZl4UKmQUVF3WGSs3NzqLbNPBhhgFX7QZ2CjvaqNmUcSHke+P55Pf4O/zcBFaYMdFoNXDw0EEUiyVsbmxZgR+837nwuQolmTLLKioqGJhIRpLYRgQnWk1J6xXyw42WhUethlK5jIWFeczMTAmk2NzcQKm8pwEF5frMOSDIRfune1//mrDpmw2Dh00rf4RARZeh4Tak902Jx41WEvxf9kkjwVQaptAPk8xQ+mDHo5ibnQa6PZx74SUNhqmoWFxc1GBf1k+Li0hPTGBheVGNBhmNMyGjosIAbfCcE6gwWwhuWl4A+GCTkr1edIBupIuxQRft3V1ceuF5dJTZYgFXo9ZPLAZl6cThm5Q3Zv3krE4BFWQfRGJiL3ghw9f7/9l7DzDL06u889TNoW7l6qrq3D2hJ2qSZjQaJUTwA7uAkcEBYxtwkHhYG9lrWHa9tjEOi2yCFvZZr+21hVmDWdtgCyFZBqRFI2kkzYw0mpw7VXdXznVz3Of3nu+79e/WjEazyPtYeEpPqWuq7v3ff/jCOe97zvuSxPJsVy5fkikriSEEUyQqMISUX8uIV8YyV9wbIYylXFYdFQqgCOCC3iV/x4MFwF2G4QLuc6oQBrjnM+UXEyroBdUkTEKTEkNDMD3MPa6Dc+S+EbTK/IwWUYFlPQF75cqYlSvj0jSGWGjs71m92rL5hRP2zm/+DssVx8kKDRfFtbUlHWtmZl73hrHB/PNOH8gsOm6aSsQbaKM3apI/29pYV7BRq++qi2hnZ1cJvUyaQ1A6NuZBCWbaBAMXL14+kH5KeFTEbSIGVtLtT6JTIU9MVujzM0SFgjPkUGo1JyqMYJX77QGXqi8d59NzVOtsJChCy6qCeP0MpBS6wrinIYg+APq/ckNLEhRDsiVWZVwjExM/NwJ4qqwN40k+G4BsMdBnrSrnRUoWR9I2i/zTAw/Y+97/l23iyHH7+V/4Bfv9T/yO1fcxP2+rtbU/SPt1yA/J12++D6pzXLvVr8uBVwW+qhZ1MFF3MCQwqf7A9ja3JQ8FeRERwyRBkSSPXo2oUHAYJI/iaxyedEmY5Ff8O4mTqq9YbWXAl7XxqVl7z/f+CesEoLi6t2fNek1eQ4z/ZqNun/rkJ6zbp5otGNIByEH4hntBR4UDgV61exXwGdRYfJ9zokAdWcx95O2YM+F8Y9eCzj3MTQJ390po2Pbm+pB8jR2HkXTgyOp2cH2+A6I9VDUl72kc8zFJi4kKUnKSBrqGPYpjK/577b0VKc7TT5FA9eyeN99tf/Nv/7QTm6mCbW5U1bUJKYlk3PLyRfvkJz5mTzz5mMC9cqFoXa0JXbv3LQ/Yn/j+P6vn0qi2rYcXVilnv/SzH7CnH311ouI97/keERWcY7FctuMnT0uucSxo/4qoGB01dMgtQ4WXey1AoF6+cMkuLS5qX8ZU/bc/8tv25NNPajCxjypRJCkMskoibRIyUHpcdCvEDr5A3nNfBcKHjoohUUXSgmxA1uMRN80+kAyK+9erERVxv8kgCUnRgToVDrxK4viLJoiSJ9K8dKDbZ6UTaIoXO133FUA6EKKCropAqvJDNoAFMVaS545rA4hIyhULdubW2+xbv+177PFHH7PPfuqTNlB3ZltxBS9OEhVxb4rjLtlZMlxXwv3NZPLae9wU05NCvnTeXIfmnQP5fs4HRAUrz/AL6adAFquQIxzHzyWuHP5qKk8jUaFnQdYqcmNERAX7t88TxvyrExXxWqL8EzJeoS9XySrXhTyQPKzyBe2Hd73pbls8u2SPP/Zl63S3rW9VyVtGUIbP8yo/HzeS30p0UCXXQu4LcRuEGL/Hz2F+Yd5Onjzh5z3wTmA6KpAZih4V10o/DdfPQFRQFQgQAZhDpyWV+56YZ6yYc+kLZIZI/omtICrU9ZMtqHP1wqMviqhjDE1PTdvO7o4dP3bETl9/vS0uXhRwTRy8tLSi/RYPtlYD8/O03XD9DVat12xvf0/ANhX7SKuub2zq/CHN6Kggnot+bswN3s8XUks8l63tDXv57Mu2urZieDvg49Bt90Sk0OG5tblue7vb9u5vepsNuvjY7Nrk5JiVykWPYei2avWsUWtLxunQoUMa53RUHF6Ys8MLC5ofn/7MZ+zOO+7SvoMEEwbU5B4A+dwzlxlpS/pqamrc+t2W3XTmOplbjxGj7+1aeXTMzp6/aEtLG/KrWLy8IgLgHe98uzpDiP2IVcgX8J5YXV21O+64w37n9x60++59k33+oUftltvO2Mbmho2NVZQfbW1s2H1vvtv26XTIkRvsSwN8Zu6QNff3JPHU76bshRdeshqFXHj1rW/a5saWHT1yzEZLo3bzTTfZzu6uvPU0N22gPGdufk7Pan2d/cqLXyCjIZCIR9a3Nu2mW26xLzzyqOUKJTt69KitrqzYpLpiBra8vCwiD/kvxifSb5D65DYAh5qTocJXsiHBq0nVwZJtc+8OyXoANAKUZhmbGcul+tbYXre3vfVuO3powjZWrohcanW6Njkza8Wxijw3PvO5h2xru2pvfeA+m5ibtb+qjgqX0vvqX18rAfG1vu41Pu7r9OfS932zZU4yZs32fu7Xvk5HNZv4e++zkWLBehs7tveBX/m6HfcP+4FuX/o9dduXcwWbn561+UMLtrqybsePH7fTp05YuZC1RnXHqrtbVm217LmXXtYaVAd3SOesWkeGrm2WKVmza1ZrtqyNp4TWZABr5lbHxqOMeLenNYUvtPchJ+rtph0/eVK+CMzbCK7zGuYaOTFYijodtCZ6lwBzEzAXYJ2/getAfNAVJxlOupvyqHU4aM/6JWUIdVU4yehV6V70xN6uwoOQP8W41dUNsu6Dp/3d93jvEPAiG/IMzos9ADKVQtlIAiRzMV4r341EcY7Ld1J82NA58TP7ihfbuc+YA/EH3RYq1g1Ff5HAiblrfL0wMEkLez4BlqB7WUfay7ElzhP5c7Ay1qdYpY9SiHLLfl+4FvukYlOIE4iU4HnEngI2wXH5mfvO/ggoHz3xWCN5pjw71mv35OjqvyGhY77i/nVOfoD7eEF0kDkSUZC3xz5SGU7JN33Htu41X2Bb7tuAoTnjxgtqYyFyVKRQfIVRedP3+Zj3UoxA8W+vWbUzp46r8BhSG0KcDkfk1Nsd5MyKNj42HnxPkbLfsHrTSQoKMSHARTyMpNWNKIys2dL5cd8pRJTXlQogOpKRxEeKfZ7nIcxF+bRL68fuTWGyujdeJMhzIjaK3iJSMglkDe/p9VyW0f3V3uio+MO+jv9Xd33HZVbW0iLDIsZkZwYR7O5X3QySRZTFXd4FGYC1lAFmg61Jt7fbs3wWQ2MYQFqdWXQAfPqSNZiojKujYny0ZKdOHLFOExkY5ILq0mpnWSX122/UrNns225txF48u2iNdsfyowDsbjJIsAnIqmpxkvSRgQBmr0pzoIauA4ADbXq0/wUmXcy22vkO2OtoJsziRRU5GxvHcOYbAqHhzHWQ9BBrrMp6r/IXmB8WXhY+3RBtyF21V6uFWsw5fhgul+IViCyc6FcXtfhQecMixX1m46UajI0AEHZ2ZlYbjyq8MrQytqktdo1DAHZ0+oJWP4sbmyLPk6orwBIWce+G8FAYNluLpBLqlI2OVnTdqjRGloNWylDNzbPkeiuVMSWG29s7+sZTw6Wf0DVsWb3RsPm5OSU1dEyUR6nCGtjlK5ekkRx1nTEE5Lxvu/+eUKnspu3ShwzGlWxYAhsDUBJln/gdmw33m2fDV7LDQRqHbIbAoOmRA6Li2ee08YqoCB0VI5mszS0sWKFSkZYwNSH9lNn07LTa8/eqbq4XiQruf5SbklQ7m4Ha77rWHcHutWsFukb2du3cs09bo0Fghpk5FR9upg0AUVRi5NrxPGc2/GjAFQOZjHwJkBHzasMItvB3QJ/1lWV75plnPUlHIoEqasl+la0fwBuvosTTwU2WBASnUyIqFNyEboshMJUF9AIwyQhMgahA15ljAvi5DvaB1M8BYUOg4VWxfEUALZKE1JhTcabKD7RMpWcfjEF7HUvlsjY2PmmVsUmvKKxXReJBVBw+etre9q5vs1S2ZB0On+nZ6uqSzn/2kJtYMjaokmN887M6dtoNgcCNWlXfe7s7tr8DQYF0FuSFE21801XEF/eoUsnZ2HjFZqZnVcW5eBE9Yz7Y50UEVZKAsX729pDhvhHBWo2PAFp5RWhO84P1QP4eAnlc6k3An/eaeGKuJqygxZkgK+IcVdcQAGGspE4YmV9LVCSB5CRYxwlH4FGgdELKiN/HZ5oEkyMgF5/jkKgA2M/TRdWwwkjKJgslu+XMTfbf/48/YTfefZ/9i1/+kP36r/6KSCgIKYgKWmaRsOK6YwAex7uCYzq7ArHm3h0Ovg475cL9ibqp6cGI7W5uOZAgo0x/ZvErgpfxv1+JqIj3x6spvUpnSNh8FaJCgCH7i8gcN0LLl0btv/3u7xEZI2+eTkeyh1SbYix/efGSPf/s0zLCjVIyUaokauwORqL820Eb/PCChGscjMshqCySBVmgCKyGqq/wRl23xquDgsyV7a0Nr9RnbQh+QyLYE51Seruu5WoN/iSpE88ted/UfSZT8EjEOSCTJCfiOIzv4++eWHF9KUuPQFT07ejRw/azH/ygTc0s2EimZGvre9JX5n5iVr64+LJ95Lf+nb344jPaC9C1N+Q04wAAIABJREFUZ+PF0HH+8FH7o3/sj9ub7rxH5uY9ijIgKn7uH9nTjzzCaNR+ehCN+Hn+8T/+fXbq9AmtCZDLR46dsBPHT9hEZUxjg2KO0XLZvYVI9sK6S1LWqNYEtpJkUrH84Q9/2B5+5GHvGIjyj1qP2ct8XYzVYcN7qQr2IMkUqgj9UThBRW4Sn4ES6K6bvsbfRaIiJukxDoBkd7LRJaCYy3H9zoY4RHrPknUKmr7B74j/9i4v961ySaDM0Nx+2FGhPatpdYgKdubgLaGuJ5LmQFRwDZJ+iEQFgD7ST+WSnbjuBnv3N3+XrVxeso/91n+wfrdpNujYINWT87bL8x3MA4/lPAF2jeIo3eCyU/H+IpNTLFWkIR+fR1y7SSF5EhkVwHjlW5KoGGru+UANXbNO0BD7RkIujuv4LClfiYSvDqoOQ+9CHdC8hXdAmLfsxUNiL5DE0acirvF6tiSp/dAREvYQTH4hKki+89m87exu2bHDx219ecsunD1n/UFVHRV9y4bn6NJdvg85ORiLZri3sesi3mfv8soqF+B3FLMA7h8/fkykshMVHTt77qyIileTfoqdLrGjgjFCvC5ZywJExbKSfj4fooJx1G7VBXDx2cQngCQjKc9R1p65okQCQKBQAjxp2dyhQ/bmt96vJ4rO9N7unggcChhmZ5FVAtzyziFJiACAtZpaB4k50yUMnHuKm+lAoCtCUmNhbHF/o54Zay6a7hhwArJvbW4K+GjVySswA2/a6tJljd93v/sdtrW+brPTU6ZOWORR2t4t+tKL5w0ibQ8gftQlWGv1fd1fQBNivytXlm18fELedlcuL9mx4yc0dogx6CqB7CGX29/bsVyWQqesXX/6hNVru1YIcr+50VG7cPaiLV5ZtUNzR6zR6Kg7gopTnjFAi3dZD9xTL5+3yuiYDKLpDlVhVrFo1XrVpqenlPvhxYRHIbreWeQr6RjJZezY0aPW6rREpDT324rpCmNj8uVDgk1+MJay9bUNdakBCJUqJVVJk8dVJsZEJCGZR9w8OT5unWbbRiGR8nlVFWvFTqfsytKKjkfeAvh09NhRAaQQLqqmTlNdbbaxue2V3/WmYjjPO5yMV5FZ9J0ZuLcaX5KaYWYi96kOyr71Oy3Lp/pWzuftLXfeYP1W1Rr7u8onIMRzxZLNHTshQAszbTp7TgDUFvL2Nx7e8P3wNYmK4c7/Nf+Qf8cdVvqj77L0sTlLz03ZoNWx3vKGNT76Wav/xv/zNR/nD/LC6V/5Kcs/cLsOsXTD9/1BDnXVe+cf/ZeWmqhY98KSrX3bX/m6HfcP+4HeXnvE8umsfCqsl7Kx0Yo6g1CxyGXTNj8zZvOzEzY1UbF8edQa3b4dPnrE9nb3bb/atAuXVm1nt2m54oRdXllXHE9eKekgdQSEAstg+qs502pr7QbYJb+luvzI8WNe2d5zU+cYn7MXxP04AvDu9UkRI/msd5drDqbcX1MESfCurNXc+wu8gs/1zk+XLORfXh+LV6OPQIynYvzp5AFFmL4HSNVCxagoSzS1Z3us5NLAwmcCCC6VB/b0KJMUfOQA9PlcsB3WTAB3Jz9dKskBbopXPB+Kks3Ro8CJVbx0RtzzK0pOQZoGEJt7H3OmmCtGwkZkUEJaCZKBz+H6XK6qLeyH96ngtQUBH+QswbsgBChODniYnw9d9A2tv/w9xiduHJ3yY4RCQOIBivXU0UDxInEaSgtIIgWJY/ZH79pwuW9+/8zvHHhU3PpH1nWuyViW+xalu1xyCpLJZZWUrypEczktL2j1nFCqIXi3Djq2MDuj3y4vLTmuGFQ8XOGDsQ2B1LZT112ndXpleV3H3Nnb98JSunK7wcdD8RuG8rEILyv5c+4Jz6lSGady1KW9glqNzkdxo3dVs/9wb1VE3KPIAULJr8EVu7yAL8aX3vAXCl4k3/0GUfGHfR3/r+76pmpumKwqnLDA0JFA0EfFCguwM7dUrfSUlKNNCwCdyvgiIbY3W5LhGYA8FVy9LpWG+Dm43h5V99OT42LsqYo7NDNpszMTAhfRlCfDoPWMLqqV9Ya9ePaSNWETR5jQkBJp43+eRYWMlnw5aF3z4Ei8+WIB1uYWqhGvlafxjY7F0FnrCCTH1jr3wHCNQZIaXxiG6af6OgDceb8z3ZAcHuS6pi9VeehQA/L2rFwcVRDui2Pejh87KsmsZqNmo+WSKn2o+mGzpdqbJNPbvTyBZ0GHFHGDwJqeg1ocUyMyvOYa1KYXFnhVxWZS6qTw9kFv4Gdz4nlKEkqVsibw3Fl8kk+XizgANJ2tluxHBJnD9QHAC7wmBQyt0kpc02b1Zk2qFNXqvks+UPnch4XuK+m69R4nKlh0kSpxtthBOe+ggJjySuJYUcHv2MhVCUArfgASYwW0s+odeVRw7bMz09Zvt+3FQFTQRn5ofiEQBVlbOHLE8sVRgV9mJB8Dm4KoqNZsv0YnEYTVQEEVzwK96ugp6UAIiQ2gq+sZ0d7eb9bt3HPP2O72uiHClJW/R34IeEKiaWOTDJm3b6IzHFtQOW6UWRNkJeCQJBbCq+tVY5tr9syzzyjIwRSbbqZcOi1QAtKO50dHkJ4NrZ5m7oPhOKHOhfEkUg7TMwwTJXHjmsZsuoAWEF1uCkY3hW+YXnXGZ0Cg+LkC7CWNxJKgERI/dPpoXslrhTnaE4HChs+zm5iakimliIZWS0RFozWw49fdbDffdbf1+ikbLZZlWHhp+ZIAv9lD827sbgPb2tpSYquqhG7L2l26KRrq4CAI2t/btlp1zxr1fWvU8K3ATHtP3VLqbAjE02iZDpKSTU5OKki9dGnJGnUCN0pdgx58CHyiHIaArSC/EjeOeP0R5I3gM/4NAKoOLrl5Gb40IhxCK6cnrAkQN5p/XdXRwfh2coUxJFA6yKk4qAZwdmDGmxRuF7gZKuHj+SariR2UOgCoFXTLTNLbeRXQB/ku/hXAhAlcvmid4D+TS6esmM3Y8YUF+4vvfa/d8sA32Ud/93ftV//lh2xQr8OaCrBsQ/BJF9dlhWKVE/eLtQ0yNJInMWBmjMQKaAXNQT9WiYWNiAyDnAXkvJakiNc2DGAT/i/JTT95DyJJEcGLZM1jnLNqIReg37OR0C2kOZYr2Lu/9Vsk88BcJAmgmwbwZ29nx1ZXVm1leZldT2A6GDlrMEAZgBdrezTzjGPqquDEcc6QQNEWHNd5yGiqx1wKxkFlvx/ax8NeolZ66f42bG19TXsI+6TvF2GzS4yVeO1KRkKgHJNLjZGwtjjY65VCkYCLVenJANvBVtaShMZtOG5MHH0yUDlPImfq1vzAP/xf7JZbb5Nvzepu3WrVjrVqXenDv/Ds4/Zb//7X7MK553QJgJd8BnsGuu63v+kOe88f+14rjE5b19xQ+R//ws/bUw9/lnQ7uCgAaLsUDZ/5A3/m++3Y0eOSASRpmZ2bsdOnTsungmSUPYn1i3ueL48p7mDfY+/VHGm3bWNjU/f0N3/zN+2hhx7SY6SqLV6nJ1O+XoOgqcpNMj7h2QXt/tjlMkysw9y86jkEcs3nxsFa4tX3Poel5RtNjZFxCd5F7lUwYumck+iAxh71uEwm1ciQpLF60LubwPiCDBXEgdqtXAqJNV+eV6EymjggUoexks8lVTw5jOA9L1K3Yblsh48etTvvequ9+PwL9vTTT0pSFPNp9T2I+PD4NDm+tT9LY959G3x9jJWTPovwzcoV8jY+NiVwXZ+vk/PiFwIYJHQYu9r3VN/iY0KdHKGLwmWZwreqUWJbv19XbHtRkQjRQphaWt34mEg2SuJLT3ZIQA7nu+TyDoAAb7nzeFdeI8h4ad13wJN7AUg7v3DYcrmirW+sq8iDfZLOLt1DzkbSA0HqQV5KgUz03dkT4UBUQNp4J40T5JFc5l5TTX/06DGveNcxKOBp2bnz50RUMA9lpq2K1Gs8j4aeSRC8TrpRgAFRsbKyqmICxjdFH4DUjXpVMWM2l1ZsQSwIKE1hz9LjlzXXAVqYlxzvplvO2HU338zN0rWuLF7WPk/RD9dHLMKXum7Hx0U4Mr6Jxff399RZDkABQUDXAeegwq1QVKDnQPyrTtiU5E4JTYhB8VR77pnnBb5LvqTbtfXVFet2Gvb2t9+v+YFnFd3VFPhQuFWpTNilS8uKO/b2avLE0zPud2320IxNTc/q2V+4cMEWFg7b7u6euj4OLxwJnaVDYQ7FiNXqtrp7xyslO35k3gZ9OlS4zykrlit2eWndLl1ZsdLohO3t13UMCjbKpVHdQ/ZTVdGmvYqWMUABFWvexvqmjU+O287ejt1w3Wnb2FgXMXL7rbfY7taGcj/IYqSnMLOm0zlHVXajI5+Kta1tW93asnQWv5+ucpHqfs0KubxNTU/bhcVLtru3q1ipAUCItJM6T5CrzVmG4dnt2ezUlH6H1O780cP21FPPWKE4qnO8uLhoR44e1RiC/GCf7FIYlcnb9taugDcIBAaLSBDF9sivuGFvWKR9XdaeyX4f1tLgu2i9jt10+oTdfua0Wbdm5dyI7W1tWIeiK0ZKNm+HT12na/vCFx62Rqtnd9x1i1Umx+2v/f7i19hR8bVCE16EMPq+77HRH/4uS02Pv+Ibm5981LZ+5B9+rQe96nV0SRS/8+363WuRHv95iYpR615YfoOoeB1P8a71T9l4adTmpmdtojym/e/C+UWtQeVi3hrVbUsPOsq36u2utQdpm1+YkWRNOksleNqaHTzm8nb+4hXa8a3DfGCPCnusYzTkvxR5OsmpgkPiXIyfez35z5D7ag8LRRuOM7kUUsRswFdYq8gh+Rv7AEVn7CX8DgLSCQ3vjofYdqlqV17wON33Z17rhtTunRCJjigjrO4IOgOykPBUujvwHQsTWUPk6aXzJb7ED8k7PthLwIrA0AD/WSNiDnJQwOcgtn+GF5MI0+A6IJZDzKYYRHu7H8OLZaMvVcBkQrU9cY5kmoi3QhcCuYbkl8I5yc9PklIeV/JFzkls5sod3sFBLMO6x/EwpGafc8+PnkB1j6KiUggFUB4juM+FF3XJiJxnGOJZdZMQmwRsTnE/ncFZ7m/svvXuNBXwaf93TJHPeurjxGf+deabl7UHQfYcyGJ5DsT4EhYUus95TurACZ1wXLV3X7jHh3I2OnwyA8ulBnZ4fsGuXLmiYlCXjwTjRFUELzsvkiCe4rPOnTsv+UsKdPGdICaCyIsdEFwDx2Z8aDyz5ypXaNnE5JQIO4Wkysfc23aYT4YA2RVNkH1P61yIR9QdEiTJIhHFvud+u47fSI7qDaLidayIb7z0G+IOHAuVv0yUMTofkDaCsaVgTbIkvtmwYLGwkdBBVIyNlyxXSFsun5WmP4n8yADJGcAzNoaOqiCp0GEiwQbnMylbXVqyLq1RhbQ2xhuvP2EL87PW61ApB2ubtcWlbXvu5YtWpYJeKHDB2si0DFz6w5NFJrtLP0l+IIBsAtp6fQ/aabnK5dXG5m1tXm3Hwo3cjbeOF90gD3mpvtnk1KQb3xGgh04ENgvMqcWCsglps+orEKYaUVU2qZTkj2CF5QeRT1m+kBXxgDkwvhAlfAXyRdvb27WbbrzRZmam1Qa+tramhZlthIpvKodUVTDoK1nn82vVqk2MjWuh5XxJDhUEyMDJzSQdX3JmnnPjC2KDNmra/LSJalONr2urbZJF0XUf2cwxScRsCiCyresBeIkSRRAyWvwD6OVt5rSkOQtO9XC+4GPAZZwcmKR6vN1t679vvefNQ0aYY8UqyEhURLNVnoMD5O5REeWPovRTrBb1rgNY8khUpOVRYd2OPfvk09JgHx8ft9n5BSVFJIHzh4+okuvIEarzPdCYnJlUO+bufgNOXJq9EEHq+FCVtQ+8a4kKBzcHNmg37dwLz9r2+rJRXwqrntxQSaBVTSAPgpSCrdgdoiAsdDUJ/FQRJ2bMKW+XpGuI591tiqggOS6iC5wvqmuJsdmS+bm3WjoZ55uX7hedR2oJDXO5TVCQ0bMGFPYkzJl+2KaJiUmvuOgS9CB/1VdSj7QC90AyMxBJfXxDvOUxVrK6xqiDLmoRbbZUMehJfVfHkRBIr2dTU1NO1nQxXHOTSgoxrr/1Tjtx882Wz5dsNFeyzMjAFpcvW1vST3NeMTwYiHAAoBbY18XUqi7vFL6Rktrb23ayouayUswjqvSY3xAWsdUWTWknKiZ03cvLK7a/z5p0ILFyUMHgFRuq/L+mGm4IwEWzWQW9GatXq5pLBGwRDKf6UhXLQas0Brb8G8kf/52DXkNALuVBobcuO1Dn1fWBqADUisBf6CrQe6/ZkSJJEUmVWFGUBJR5n0DOIOkSj0H3AGsfX5K0k/Gb61EX81mbHhuz97znPXb7O77FPvfFL9lv/Ma/sf5+1bIdAuiutdIAjQCEB5UhyQ4UkeahasTHlhOpqtAHEKICiOQn+PBgtCmTYgyOA1gXn1e8b5F40Mh8BTmv5DoU3xtB4GgqG2+ht0MfGOzq+VCtGcHhlNnb3/lOBaiMNZ49QTDnR6U9MiC7uzsitJm/IiqQVIGoCP4Dgg0Tzy/5+OL5v5JsFmbIXkvkxFMSyNY+CUkd1gLAsc2tDdecFxjpFdWxSjh+JqNHyUfoEoqdQAT9eg/7MV0lIirce4EuRd8nvOU63lMdPfHfyfGXvF4RWGKHnR2jivcnf/LH7Vu+5ZuxR7TNZs+qta61agP5VDz28Gfsw//+V23lyjl1rMV7E00OZ2dn7U/+yT9lJ2641TqDkhWKFfvn//v/Zl/6zCcsbS0oI1WSC2xWt9OI/fAP/Tk7fPiYKveJZcbGy3bq1CnjWACq7LWsX4Bfo+PTiicAH3e2ty2byqgIYXNzU2vwRz/2Mfv0pz8dKgadBPQ7HSRHAokpebywfmiMhXt87fiNHRVxPYkko7pQVO3nx+f+RglF/lvzFiPAIAsVK9RUNQh5mkkQ0ZhjSiohgP/qdPTOW/kZKOHyBEnyTty3wGrhKSWiAvJQRMAB1XdV51fQu4tjguugigySn+SwWBq3c+fOqpqRtcO7IjwRJ/+Ne48bJR6MeZ5ZJGt8HDvFzPs6/abWk0pl0jKZghch6PzckBE0F/k0v6esdYnxy3WKqDggZdwPipPxzhS/74GocKbQOsz10Akz9FrTHKfAw18znG+Jn714xJ+XCJVATBMD9PudYMR8IF/FuVFQdGhu3kbHp+TRtb62qviI9ZJjxTkY75f2IO0nDkaoizJUZqDDTGGKzLdDh432emKYbFbkPnMCaaW4D1HIc+HCeYFExJ4iKrJIeRx0E8Vr5XxZj3it4pccJGLJVlfXZHrNOUaiguIegINcDuDcpZ8An4lj1p5ZsV6nry7OmdlZSY5S9X/LbbfYoaNHrd9s2h7zEinXthd+MC/piuinUrZ44YJtbW+rY+BNd9xhK0vLKp6anplR/gKgfez4cflcQc4Tm/MsOD91jbaJfSH3uMa2pC2feewJa9Qatru9I6Ji6dJFSd9+53d9u+1s79rY+IQ6qtc3VkPRlNm5c4uWL5TVoc6YJz7r9lryVYOoYDwCeN95xx12cfGScgY8D5iXECsRQALkwC9wfm5axWFvuu1mazer8sRg4uC3ce78ol1e3rBMjs6NvkgJSAA6fZdXlkXQEJMRxxE3XX/dDcoV6GSlc1DEmDqYpyVPRU7Htzq1AJ5SAysX8hqPyMOwZlZrVJgW7fyVSzqHliTQvBNHBKd8dnJ28fIlyQOTk+JhsVevqbgD2bzJyqjtbmza9ceOWxl5305LRVBzxw7bE48/JQmY0dExW1lblVwWBQBo8dMZBwnGv50OsRjgZEcEqzxMPDgYkqaKX4PsLfdTMjKYB7eaGoPSOU+bXX/yqN11y/VWSPflVYEEKTJil1fXbHbuiB05c8bazY498/iTGktzh2et1mjaTz68FnTJk2UQ1wRqr/M/IRLGf/ov2UjO5ap6SxsC9JFgSh8+qFCu/frv2u7f/mev8+hmYz/xZ2z0vd+j91X/2Ydt72d/9VWP8Z+XqHijo+L1Prxbr/yepftpS/XyduzIjM3PzttLL0HeZu22W8/Y8YVDxhJG0dfa1patbe5oP9zY2rGNjbrtVcFCKnbi9HW2sV217f196wCE430jL0MKSsZUDAE5zpYLKMw6rBiZnGnEbOHokVC535GnBXku81zrOflSozH0jiIupcJc+IJMsr2ohtjq0Nyc5itYAXEegO7Y2Hjogkgrx4sS0sQUDoZ7kSBfrJ18JpgKewGxGyC/4vBQmCYQvdnU57PPgIkR13BO/Ix0XLIYyP0wHLcQGR4kesCJWFfBf7yLz3NDzxmRru6E+NmJZDChGLcQEUZTZX6nPEiEgxdZRMNs4nsRPXSu1Gp6O+susRrX6ASQA/HqkhgBc2pYIZdTHo20Fud54w032IULF/U6VCYg4lm38CFzaa1BiNFyw89WYakkP70bgutRTkVnCnlaUHfg81hLBfQHwomiAy+M9PhOeVy3Z2c/fXQ4xGNHRYxbI17kOeGBVHjcj3mj8pEQL/EvMZ/yjZAfpwctm5uk0Ag/p4b74LLOB0l0xqs6eTJZO3rsmK2u43XZ1DEajG/F2jnFDcQjjHcVJQT/COIAMBK6g3nIyA3yLOlabtLxEzA7xYuQfcHUXYXSyi9d3cbJHTpm8LJwxY3omyKMVoUY5FlvSD+93jXxjdd/A9yBw0oSHKSEoFC7vwLvgQJ+AZQkLZIGSCuXy+cyNjZRVPCczqBlS8ESgSatcgNpRmPSOTpasEzOTRZdox5t/BHLAECh65cyO3X8sN11+802Qjt/z7sSVjer9tLFS7bfaFqrN7BGB9MgEidZm3mlS9BnFo8/XHgAe6j09jY9Ejwt/uH1bEho13rC6kAEFUmA03zBgAJix3Y/wCl5DKB32HWAvt8FjHETaFX35wsK2tNqn3P9Paqgun2qOF06gMoCWNp2Ey1Dbz/jPiL5TQLGpsRijpl4bGEgOGCxjwuYNlaIhHww+0s5ECOJCRZ+6Vi7JJR3I6RFknh1gC9sbBpo8wOs0AJPZYE0DBuetPMlQIOAXdIpLnMko/LA2JNARKkoJZD5vK5f15ElqecZmrU6VLQxtgC3Way7qmKEyLj93vs8IQ66j9cSFer4CN0sr0VUcBxv6UMCK5ppkzjNWHrQV2JABRgVI7NzCzLBI/GeWzhs5dFxm184ZJkUo6hvk1MTTlRUacFkQ4OoQEM+GnsrixkSFb0uevueqFK11m3VZaK3tbpkWQxggz5lBIAhzET4IA8S2P4oKcVzitJdRIZ9SQq5Prk6ECArkGQbtO25559Tt1M+m5PeKCELmoiFsptLxnsWgR9//m6q6obd3sUyBDBFiKjWQNcHoBCJCjcLQ/qJ6kOAEZcd4rwZMxAAkkELgGgSACYJBGwiyIv+Bmo/pdI2VJ0AcnBPBDr1eqq+aXdSdsNtd9mpW26R4WElV7bUoGerW2vW7g+sXK549cBg4CBwkJXqdSEnkX5qW6vZttr+ru1CVOzuSPIAo0eOT0DMN1WUXnlJ58cBUcH5bGxs2dbWnnwqesHoLElUxCoZX0kOksx4L7w7BuAvVrz0bX93V4bwIjhUde8ycJHgGVbwh2BToy3h2zAEcUG5QmWI1kN1VkTZENdUjeBv3IJeiaiIhASvjRXXSYA+/l0amQLLYr2vY3pRLoY1EUAHfC6bHbFcasQqxYL9wA/8OfvT7/1R+72HHrJf+uAHrb69Zek2hGjXupRDUk3Sd9mbuB5EoudqwNoJAbVsS+ILPyN8YNy7R63HdCuE5AYjXL9vOuqQlIgA4tVj9AAcVGdX8Bty8MzniI4V1qt4P2NrtneG+fNPEhWdQc/e8a53Gd4FADwQZATCnH+zWhN4Xa/XJNd2QFTQUVFwkFQV4U5qxXuRDCciwBhJySHoLdkKztmB5eS1+k12w28nv/q2v48WOCaEvi4kyYSrPi8QFXEtc6LiABhWHe/QQNBl5DyWOADM43qUHNNJwiL52XG8YrvuCmdulvcDP/Cn7Ad/8AfJBmyvk7J6DXmhgW2ubdqnP/lx+8iH/7XtbFxR9W6UFGCu8yyZ19/+7d9h7/q277RBumL5UsV+/UMfsgf/038wEhaXoGS88JNX0r33vX/R5uaO6H6yT46k+3bs2DHpn3M8nidFASmS6WLFtnd25T3Fns8aff78eZGx7MsPPfQ5+8Qnfs/l3SLho7HlMYzmQZAS8k5G71RJkk3J+cyEi5IhvCYmvfE5JNcPErFoDikDbYDaIO2VJPy5Ztg2yTuSLMnEPnjEaFy6dwNJk2IsFcg5yE6XA0RF9M75akTFVePsFYgK7i3znSr31TX08pETdSLWn1KYc0O9aScHuJYhoQPwGYjDa9dSiApGFRXshULlK4gKgGueuc8fil+iVJ6baUeiAoLRf/bJ1R842BAloyBifXGQ0obOWmShukiYJy5LoWq8a5nk8LCvJSq4vw7oemxFQUhc8+M9YF0cm5i0mdkFSbheXlxULAZA/UpEhcZYNBwPhuHDdS0QFSKP6bqR6baPT3nazczY9ddfLxAnGpUCHF+4eEEJOwBRsQTxVLBux2PyuN7HdcvlM9yzBWAKv4X19Q2rVuu6n8QaxHd46gAQ01HBGGH9I8YgHm9eqoqoADjKF4hti5Yr0F2d1Ryl61Q60EilVus2ivee5DAGAnaeePIJm5icFgGhisZOW5X9tXrNCuWyAxBG7O/So6q6heyQTNWSzc7OCRRqNmuaP3SvPPXlJ22AZC0d0cjmpsyefvIJe/c3v8129mqq7Ielbreb6hrA3Hu0PG4XFy+L4BifnNCz3dvfscnpKZuYntW6duHCorTjX3zxJev1BjaFJ0kubyurqyJRGFSlYt6q+9s2NVmxvZ1Ne8ub79R/Vyol9+vL5OzsuYu2urFn6TyVquRKpnunLqHBQMQFABcFYjyHQ3OHJH2xt78wgkjMAAAgAElEQVSv4zNuS6MlyZeNj1es2aja3MyMrS5fluxTMZeVb12ROBCfuhTSti0rVsbt5cWL1oUooFN4fcvKpYpNT80qdiOv2Nzass3tLUmw4ruyubejGJd9s5TP2UShZNlB32Yn6cxvqWiuMFoSeUOHP7JuxHgUmTG4kBLDy4OOn431LXXrkANlc3l1HFNIlSR53IfCO5qVf3E/AiipTnzGLMR2r21H56bt1MKM3XTDcTv3wjPWbtRsambaRnI5K46OW2Fswna3a/bZhz6rWPuOO++00YmK/bUHL4dt+etFVIzY7Ed+1rI3n9RxGx/5jG3/9V8cbuWQGBM/86P67/7mrq3c/xeS2/zX9PN/OUTFa3dUIH/V+swTX9N1/UFe9P/X5/xBzpH3vr3+qI2XK5YZpK2UL0qy+6WXV7RenD4+ZYemKtau71s+M2JjU1NWnpiwmRMnrNNo2fLlZVtZ27X1jX11VTTbA+VjdEp0QgGBr/+sc7gkemxM3ASQLn8mdaGP2NzCvBfJqcjU5YkjWcAezvx36TknFCTvRNxfx29zVPkbuRtrtar45WfZEUHJ5/DzMB6VmbTvmU4oeAzDa5jjXgnP3u3xthc+eswfC2BjzBaLXVlv2Md4bVTfiDmU/86Lc5yo8QKfGKNFgJ1jcELqYpAfKdfg8Qv7auxo5yBU9scOc97vx8eYGRDbPyMqTcS9ORIWkvNGUgqCP0thcV1rmZMJbQHhRJL1vX39ns9Fcnx5ZUX7KveBbjXlsqh3KH+gG7upLpWI3/AveyR4YZSaYlz5vun5VLy/bljt8sb6zCjJHnzYYvdwsqPiTd/BXnBQCMKxhBWFHEyeGpkDk3R1NKuzBHA/q5+FhXCPlZfTWluzqQrXYOrk21hb155HXk03vAj6Wk0KE5xTvdGS1BlxieeIZoVSWXiaMAGCGIo+oyQrJF7G5aFd0hsiAS+OjLo3kT7jC6JOa3IgUFR4SdApyTPvclGM0/LCb3X9SenDVUc8xkQGzN7oqPiDLpJvvP+/vDtwPBg2x8WGRSpqvsdkwmUlHOSQbEkqbdPT4wKdCbpajbYSdCb35KSb2HGchflDtry2ogSMY3ibfN+yqrJEMqhjxVzKHrj/Tpus0I5tqjqtNbq2u1+zerutjZCAnrbkdndgjSYbEEQFxpG0EqaU3LtKglcfAywCFPgG4Vrcgmb0OjcHIqiNG4YDt96Sp4nPNYYWxNgGHLsV4uYnogKfiE7fTdNEEHi1oTQHWakCAMFrqURn885lMq7lnqO6rKONQywqgLQkIVwTDyCA8yHBimCO+2K4LqNMaQdo3o1K+w/WGzkKNl/AdteZTVur01FS4Ru1J9U8C6Qnoolv1JwWKJ3Qp1eFNGbnjbqCfirj0ckFZAO8HC2PqvJ8fv6QzrXeqIqcECnRaXmXRdcr+GCVBWQM+nbrm6/uqGBoRVac40SwNwIvsaMitkmSnCYBrkhU8AyEAKQwG5+y3IjZ048/qerl8fExERW0j6dSWXVXoBc4Nz9rqZSDuxNTdBQ1rNpgo8pYpztQFa00IEXWuN6hy5pQmdp2KYdAVPTbDVs8+6KtL1+yLNWBIeiJ58qzREsX8J2uitj9EK83dlTosxjXkvdx464Bor79gXVSXXv55Zdte2NLm28uhTRSyauWQ5dRBGT5XBlB4ukROiriuAbUjXM+mwNQlyJvqDbJSf/YX+tEBRs5lW5+/d4JwryBqBDIADgDuZXQzed4gBvS3gxVwi791FEwwKZMp4t38HglLMFfp5ux2+5+i80cPy796bF82djrd2u7VleVhuuOM265DiSVHOjDFBGiAgmpllqEq9Vdq+7vyjek06gJLOY9BMWYQ0YQszKKGX1RHRUQSnt7VVtZWbdO29eTqM0/DIoCMKjMPlZGh7nDfYsEYTRPdR1Ql3/yIGQgGZVrCR5VBQcvBpd/cYOzKLfjjSpBhkmfGyphBXjx7dWpccwNwaZX6KiIzz/ZWRHbsDmvKBXD6yAihkRF9DkJwDSGohB9CsTTZrnMiI2Xivad/8132l/8sR+3y1ub9o9+7h/axRdets5+lXIt62H8rmqg4EcQjpX8/GvvTTTJ0+fkgqFraF1GMoxgUXJUIeiLu20cW7HifAhkhnUnvk6Efehu8SD0oPvlK4gKR0A9uPTwc0hUiPixgb3z3d8koAmiYn9vX4kXY59K6LXVVVtbW72KqGCvyUBOAxBn0vK80ON+BbIi/o61MK6d/qxJsFwWTIUFCSJFYyJ4AUCOs1dubm5IruS1iIoYC7gUjJMUyXOLHRUi4SAzR1wazvdPv4/xnsbnEI+ZBK2T49U7M4k33BuDufGt3/pu+/Gf+HFJa9UHgF59azUGtr66ab/z0d+0j//2v7O97SXL5KngdnM+5jjeIMyrd7zzXfa93/9Dli5MWq4wah/+9X9t//E3fk0dFd5vRjLrMjTIW77vfe+z+bkFAYrsg5j5zs+jx3/cOzVHzCYnpywLidZPy/uGZ4vMDpWCignSaclrPfH4E/bxj39ccclB0hx8P0KsAiLuTSTBSD54rcRnHMeqKsVCsUZ8DtdKXMbfc0+TRKTmWIKoiPPfSboR66srIMhfhj3Bk3GXqQPUJT5xMF5mYTqtLmBFICrk1UH81gLorGoPvbZLZxgNMy4TZCW/Z39hb2D8rG1semIXiifiOPcE72oiL3lfVaGdICp0z8K87vabWtPKpTF1VXhHhZMgcAvILroWU5Be6LkWdbKbgz3NX+GFJ+pC7TUDURFMuEPXiQhtcnLlrAdERdwvvTzygKk4mBMOGEfppzh/9TtkuxJERVzzBfTQrVks2cyhBY21K5cvqQBFRFggWnh9XBt9fjoRzTVKhiKSvKxL2byqCuVhI+LGqzFJ5Ofm5uz06dNBZsGTaOLQixcv6PwgDCAqAJEiUXH1PGe4s3/4+dB9zLlvbm5pH45EBbEIHWAAOjz32FHB67ne2cGYzC15EADxkrdoU73P2B1oTO1sbctEm8lO7O3SFgO7dGlRBq/EXBhJA/ojgcmc530YRgN0U627u7tv8wtH7NiJE5Yjbu937cknn7S777rHpVrVodqzva1Ne/7pZ0WMvPX+t9rFl1+2TArwv2kzUxO2V2vaXp3uZ7qjkYr1QrH5I8fs4rmLKrA5c+aMKnCRoYIQ4H4Tvz/zzHN29OhxW1y8rNchvQVg50amLnFC/N3u1GxyvGLIE913zx22v7tlpSKSFBnLFsv24kvnbHl9y9L5stXqXrRx6uQJu3TpUpC3Yo6U5U3HGMZrgvwD4pDPZS2j8InirJ3tLdvf3bY333OX7e1sCcQ/cfK4uuIoEmEdZA0HjAPi//LTz1hpYlKFaKurm5bLFu3EiVP2wvPPiwxmPi2vrVq7zYaSkbyke9pLd9JKmYyNl0o2MzGhsa2GoExKvh3pTEHdIOQnFMPki0jsrqoZiWI0lpsWHV/KpTDlpXgIeTWPnxg/ybV2hOKhgXvsebGSF4UV82lrVXftzXfcbEdnxm28mLHdzVVdM7kGHhWTc3NWmZ6zZrNjjz78iADDhSML2qP+h8+thNT660NU8PwWXvx3OiadFKvv+pGvAB1mP/JzQyJj53/6x1f5VdABkXvzTcNuDMiM6i//tlX/6Yev6qS49qCv1lmR7KiANMm/+x5LVUoeNyWOnTze+N99r6Slhq9Dkuz3v3QV4eIeFVcTFYdf+g0dpvPcBUsfmhzKXvVf4f1fcVPMLL6//eUXLDVescxpZIH9q/XQk7b5Q3/3K972SveL10ZyaOqf/KQVvuVevS95r5OE0av9/g8iz/VK18fv7tl80MZKo1bKFmyiMmkzU7O2xBwZn7DjyCDjAdVtWrvZsKXVdWt02i7ph8dOu2etbspq9Z7tN3rW6kC+p4TToMqtLoC2e3dCNtNFTvcFxZHk9b67upTsiVOnVKGvzr2AKQlf6ruMnsgGfAWC5LgkElUh796QXhyZ01oun9TQ0ahikyAB5JXx4DK+1pPbO+HoUtba83gfy0aafL8joDvGS3GP8lgoSDCHOC12JkRiRuA2BAifGQgQzj8C8ih28B7WZS8mdIlISHdYUoqCyYPVzRE6myMREkmT2P1P4aJX13uex/uIcR2Mp3jB/RhE3oSiANZ7zpG9U7JHGI8XqOr3ItURCADwpUHwAIF/5XXgbIOepZAqDnkInRqKR4VPeHyvXLzZ1BhwLw+66TyfZ4+I+UK89yoKS8h8Rekm7lEkIHjNlUduGA7lU2+/OMyFYk7BHyMeFDtOIpmRHvFxIUlJ4WzB40Fy9Ai4MxCaNjNZUV4OJgdGiYysiIF80aqNupXKYDYZ29nb1XgGX2i1kZxJSekF8qa2vy8vKAi+dL9vBeIkOnfp+iee5L7o+ZiVxydkTs85yduDc/Taa4WAnHOUUY8ERqfVVednlznYaKuYwAkQLyagK5jnIZ+lN6SfXm35e+P336h3YKrRHiYk0RxPZALVlaGK1CuofINhEVWXQAYjzqaqxvly07OeVcZGtVCxWEMisJA2Wq796UAJ1UVMyp4ALeD5yijt11SQ9mxqsmwnj58SKNrsoG/cUPtvo9m27iBll5fWbL+KnjQgKhIBZREmaoEPld3eEudMI4kVx4ryCTLzjZX8SjwdCOKHmLglK2m9BNUNj5zx9kpEFmokeSL7TpYnNjSA0xAP0lUc4RyL3jYozT+MtIORkdrwfcPkHqWyaOC2xZLHSrGJ8XFtnl5p3hbgFQ2WqBZT+1d/YHrdSEoA7dvf8TZ79ItfkoQUIKtMHHXdYHgHpE2Smecpcm10kLBxUb2qTggZMLshN9eM+ZzrMnaGLLX0W8WYh2ppNmrMgVIu/8TvkeiKnRW333efrpn7FTUEYyUzoHbcaGLLZpStSBIVvJ8NkMejsYoOPHp9Ga9CnQJwLhbs4Yc+L4AwSVTgPzF3+IiVyhWbnpmyfA5A2GxqelIdNiIqRpCdCtJPwaCTLMkleFxagwp+eaQE6ad0v2trS4siK1LB+CsSXzGgqIxVLJMrqKtDsgNUgwdGPILbVCMzFggOouYlwBJzpzlo2eKlS3bl4iXXckYqIZPVs6BCn4DAux28pVQgM8eHQIqGUrTKhoDAZbw8KKRjgudP5SMm6/4cwGv6mkPeikqlMtILrr9I9eBVYHiiIoWNnvNxyTgHdmVUhV9Dy1tpR0fLSs6jTAvnnMuP2W333G+lqWnL5Is2UahI+mm/UbV9teAG/Wwljm2BgqoK7lHlUrdWs2PNOt43VZEUeFQ0m1Vr12tas0jm6cRAco11i/OnowKigs4bADKCh+Wlddvd9Tk0BG0SJtlaNwDPhlIfDtZLRicE20giAcIRsMaxQFDD65AjUEIZQB8H4g4q1b8SoPZgnfXO1w0qgXg+3k3lnRVOBvIVn0sEsCIMpvMOf0/+HEG8+K+SSUD30FHhS6HLInhnnY+zvZ09J+zQ0lcnkQlAeNsDD9jf+Kl/YJuNuv2TD/1z+9ynHrTObk3a1T2IauneH1xvrDKPeymfFav8WX/iGiFfm9jxEJIDkAfavAUUhXU6nr8XcoUAPLTaxnsbrz9+ZiQxkuC5XpO4Z+HmHTz32LLL50TPhdSI3XPfvXby9CklEXQVAdoyF9rNpr304ksiKgbIeEHSBFm5SFQAloK7JM8z+XPcd2LnTqyKd+PbrICd+Pq4nmo9QP5QY5EOgbrt7GwJ0IpdPcnr5jp1jEg+Blkovx0HAHFMpBzg9LGYSQeviyA4lhyL8blE8uLa2Cn+XoUF6Atrb6F4IGVnztxgv/RLv2gDkqFUwRqNgbWbZmsra/Zvf+1f2oO//zFr7K0JJALI5Fh0s9DBxVi688677E//0PusMnlE/jcP/u7H7d/88j916SeenUrjkRcAnB2x/+5Hf9QmJqaVCGCKV63tqdsMwh4AjFZ+9vdsvmitnmn/RuaFPYdnGn2VVtdW7eKFi/Zbv/VbLq2ZkL6C2Nd8prpOZoxeba97HGKoWKGXJO80B67pGIpgfJKsjmtMJCuU5Il09k4q/TewZCD4ZFQdJAIjeR27KphbEBXy1VE1ZADkBynrQWgnpZ/aHfmyQAq7jNCrgHEJoiI5Nqanp7V37de8qj6OUXXTxXEleung66r5fA1REWMtdTf0W5LWzKTzNj4xLVnRKP3E3Otrvjv5qyq8vscrGsdIP2k/g2UNXWbOEcr/wc/Bv90q3a98kKb72OcaBj2M7yhXJWm5r9JRAZDtWlL4noSOBPmOHJhpJ+eYr515mz40r0q85StXrNGoae5zNsSNSSLW55yTKOHUA1nlHXv4QHg2fSCLw3vYK+kuOoaRtgfTAeDuykcBUgQQG0lR4oGk9FOMs50Qp4vH4/Ao/UQshgGyE+CeZ1AMIwnAzIjmncdQBf082QFcZv+lWtbvFRfDPM0VMwKPL1+6LACb2Ml9V3yOrq+tq8qX/QgQDMPlfK5sxQJVjA3b3dmWrBLPk46AcbpVDs3a2MSY5QpZ+/JjX7K3vvVtAn645mI2a9u7O/bY579gczPTdvLYURUmZSVN68Vgg0zORienVO2/z2dyndmsvCM21zdUVIG0SZTZ2t7ZtHptX2vOgw9+1m657XZbXlqThMTM9IxVxsckhxJNoNvIrlrbxkZLlhp07b577rLq7pZ8IzBybrbbtrm5Z2vbuzaC/BVxJ/rk9bpNTU1rP6XojJwB+SfG16mTpxS3YcBLDEWRFn57dM1ksikbH62o8AeSstNqSBIKk14VVOVz1qrVrLpXtU6/b8++fN5SVECn8qE4KGWlQknzh0Is/E241meff8my+ZI6HnyO0oU4sHIuZ3PT01bCF2jfvSxmDk3bCy++NJQvBYQ9egTSI21LV5bV/U/82mi1rRVAJuZeq9nQuFfnThsvQZdLYX7JqyasN3TrOCDmoGo+M7BBp2533nK93XLqiFXKBbv44vPWQ55qdlo6/zNHDlsmX1Kx3YOffsiq9b695f7bbHx60v76g5fC+vD1ISrGf+LPWjnIMrU++ahtyofi6mNT/Z+/3w2uW194athxMPfgP7lKGiq5riITNdivDyWfrt2zvxai4tr3aK3fr9vK3X9u+KcksXHt6yEQNv7E/6xffzWi4pU+h9+9FvAfiYpXe/+13SnzX/gXr+oB0nnuvK1/90/IK2Tsx/+MDpl8f5LASJ7X5M+/34rf/Q69/loS6dXO6/X8/m21h62cL1ljr2oFyIqxSQc/Wx2bm5myk8fmbbyc05rRG6HLqG+Z8TFbuXjJLl1ets4gY9V6z7b321ZtAsKOGGI9kjBl7e97BT3KFdX9fUn3IS+NXB7ALF5HzCFIYYpFKS5EEhnSnYJLFbDRQQDIry66juHvR1xdREEgB+FQG2IrELeSgpX/pqt3gPnggyEfBBXmuDeW9lsVkgbZ2oD7qBs85F3Md+IztjpyatZDcmM6L8AbwEUgXnirGxxTpe+Frt6lTEdJ2jsKgsSSx04pkczKb7U/ga0gf+v7VDbjsqt8idShCy/Id3JMYhDyCPJyOhmiygOvjR6pnnOSq4cYki6JWl333PMo96ukowLEhmJWeVMSl2D2rRq4ge1v7woLSGdzNrOwYPvtlrXpxqSDEulqpPLUSeP3OsYdMb9lT45yq1yP4h0IxAReFn+nIiKkokIuGWWlov/g4x9DTtK/8KgQIRMKkPgd9yxiRnqRJMCRiSff82Ia7iN7HeOJOAJFlyzSlezTOYqrK9ZGmrdet4W5Q3Zp8ZJyW3I2pMInZ6Zta3tHHSgQ23gNZXMFN5KXwgr4546VchToZe3k/IJNj5atXa2J9NhsNGx7vyq/Irz1xlB1yeS1B1EQ493JjGHwVPcBw7uQb2YW47jT7FpmJGfWoWsjKwn1Hnv71Kjt4iWcyjuGyd74BlHxepbEN177jXAHFvopTcAod4R3A61ibkztxjOwphANakNSRbMnhwRv6Jlq0QmAMRuPJ2MZ26s6IMf89HbvICMUnOwbtarlMoDrDRureCvt3KEZ6eVtb28JNLz55hut1SZZrUrb9MLikrW7Kev0UtZo8zk5a1MFwMRW94QzvwScVO4QZLveuyec+grV2NIQDO19bhbtnRQsvJExVndEAPWolIrAL5sy1++seQDbwsLJ4s2bWBxJRNHWZuGG5JHWXDqtZAnQ1KWpRixbyNletaoKLrVDBlNbTjduANo0IV8ApwsF26vuKjhA+ueB+x+wZ55+Wp0kR44csaeeflpGxTwDqnO7ep5OFHEOcVOMIAULs2+yvllyTVSvSXIjS3LWUAUpyZNaqYP0DpsGPgHR/FZSTz28KAD7A1GhjgpPqNm8b7/vXp13rPyLm5kWa7xFAuEUrztJVPB3ggDeH1sjXT4Jw9qWzLQjUTFRLtvnP/uQ2kVJqGcOzatamSRU2tcQFdNTVii4kWUkKvYxURYbH6SfXoWoQIc2VkECqGHKtLOxYudfet4GaAtLz9srHzxAQdKgpAAAdp3riO2asQpf446RRZUD8w49ZaSfoOIJDtI9VYmdP3sW0R/LpTNWQLYF49O0V35EyZP4mfpvghHpe3rwxVf0YNG41i7n1ZBIKxFcCkBXZ6YHajKMD5XSnDdrA2DntYlQnENoBAscC22rAmWkkQ7x2NTzi9efPK/xiTm7+c57LT8xYdlc0Sr5UZmTN7st26ODot4adlREokLVrvJEARRuW6PWFEFRre4pua/X96wtL5qmvgHP1tfXRVRwn5AxKBbz6qig84Wukd0d76oA5CSgiCBYBNQF7gQNeV1zqKznZ9ZU1sGhCZY0Rr2qXJ42mFAHIzjpccrj4Ss9BZJ7yJBUEBnhATEVzQfkmcvd+fdBNb4vea57r1guUWWvv4Ugnp8jGJf8VxXXwSeDawgQnmSXONbO1o4TNiOcE/PArFIq2h233W4//fd/1raadXv0qcftQ//s/7Ta+rZ0QHusDZLfO/DoiB0c8RyTwHyc66ropVJHZsRU3wYvC1UX+/imUlGdNg3My4OefMI8OwmyX7tHJ4mKeL8jUZEEl8NN19vdyNb9KURUhK6+e99yn11/5sbgUdFQoM7+iSTQ8889p24GcMyriApkKAj+iWkDOaK9JtHFENfL2P0R94q4ftMxRsdhrIAaEvhMZmROVDXWl0QR4CW/1nULAjr40ueG8e0981/Z3TEkQ2LCJQLUg+kDobC47R7o/F9NSjl4GsdpBNtdLs6ln7jH/H5ubto++MH/1aYPHbLmSN7qddb9lF26cMl+/V/9C3v085+0/d0VJa2AXIwXKsCY86zFt9/+JvvBv/SXrTiGtnHWHn7w9+1X/o9f/AqigpCGqqUf+7G/YqPlMZkSk6giwULBwokTJ9RZwWcorkA6U4bbPSXdKijoUAHeUnKFH8nK8op9+MMflkFsJKddK9iBZxmVy4vo6o6KmKjGJxPHKOtLfMbas6NMWWIfj/dUyXkw1Ja/SvdA7i3OdV0HcxjAWOaIxHUOuHtHhQPVJE4kV7EjM3ZWDEZ6TryFlQZAHfknzLQhEFkfYs3+VfPuFYgKzjd2kzbwOYOAC4nnAVFBlTP37kDe7WqiwuO95Lz1v5NkI5mEZGHWxsemdS1DokKG2gcdFX4fPPaLREWY+G6G7YtA6EU4IJEjUeHrB8qotOZ7dxHBhTy7g4ySDCcTREWSMNR6zsx8BaKCeEvfgbhNkszsYZVxJ9M21tbU2aIEPeVFKarkS8xpxcJhnsdOFSeHkCmgcMnlMPg/1gX+Bglw8uRJyRD5/dHqrXgMjwonKgpWKOFPAFHhxHw8T8bskKhwT0433y6WVDQSiQpAa/mz1Q+ICohIFfRk8wK7ynWkJqmkJ+5wSSbuHBWoxLCA6uurazY+NWkj3YGVKmPWpDo0lbIrS0siWyR1K7+M+MzxdyHeQDYzJ9mndK5o7UZLYLu6yjNmjz76iH3Lt36r8ibW+Fw6bRfOvWwvPv+8LRw6ZNefOmmtRsPymjd0KbfswuUrli9XbGF+wZaWl1QIsnhhUR0KkEzxGfAcp6em5LkBSVYqlm1nb8/KZbxbztva+pbdcOONGlcrKysCo3ytRnZlX2bWpVzabrvpjO3vbNpoKa8OaXzSNrb3bWl9SwDKIJ3RupUZSRkFNQ8/8oSdufGUXbl8WXErHYvIfCFlR9fGI488Il8S8g3WaToMGrWaXXf6pGIvlpGJsYrtbG9I+nd6asIJLUvZ9u6edUbSVm31bLvasEJpTHOMjpcK5yYDWFPXxoXFKzY6NmmNVt3NzHNZyyPP0uvZeLlsk8hy0MEsAitl5y9eVBESY+jK5St27OgJdarTnYPcE3G1PA/TWe/0SpnAT6YfayDEj8tpjCh2VRcLICpxmiqBcaADXExbv9sw69Tt2Ny4TRYyduv1J21rbdVGINbzOWsPzKYX5m1q/oh1+maf+dSnbHJqyk6dPm3rO1v2U1/a9jXq1UjcawOU1/jv1yPLlDxUEjinI6H2f/1Hy77peit91ztsZLQoQmH7/T8vgiNz3ZFhlwAge/fslasIj+Rxk8QDHRSN331YhEf+HXcOuzqiV0YS1I/dFhyr/Ke/fUigRPD+tYiK1ueess7TZ22kUrLS975bHSLI5279yAdeVQoqSVS80vuTUlnJ6+J+NT72WUuNjaoTJPqARPJm4cv/SveQ161/94/r9iRJjmTnS+x2GVQbtnzXn32dT/+1X37v9kN2aGpGhtpT41OWyxRsbWVdYDseoqlBx7bXN6yQTVmulLbpuTm7+e47rbq9q86meqtv5y6uWKMzYuvb+1ZESi2dtlW6iGzEJioTwi8WFxeVH1DgRi5UqzXkSTBCZb6N2MmTp6w0WtaaxnwiI2WOxcI/KtldfjqlKnfWJEB0l5J2opfXg/OwP0l2cMSsWquLhCXvApAvFQvqpnUlCgfE2c85PzAB9n0H93uK3SBI8RhFpk7yvB+6BcQAACAASURBVCrs9CISPpP3QLjSZQYALrJ9BGIi70oV8tFwI2yNXUlTBR/TIKWnIkfley7Z5PhRQrKIjsCie+NE42hJQgVQ22UwvcOUL+FbxGgiDTyuk7SRVBJcxl1FKZKyo9DEZa/w5FG3CJhJp22jdHzsVm1qYsrarY4traxaP5PR+tVElp0OiHbH8hQ3ckxixNCBEnOPWHwQOyRi3kK+TRwipbwghRWxihjrxPdE306u/8sfRarPv+7/Xu9WZT2GRGcccH+J7b1oErn5svIsigPJH5qhay5XLOhzIYgk0YtHE+S0Id1aFo5CAd3k+LjUSSgmg4yfOTSnzomNzS0RbTwrsEg8pFB4QZJLRNzOpuUyPRvNmt116002Vsihf269Ttt66aztoebQ6lmnn7LN/Zpt7tVsbHJaBVfNUHgSi894vsJXsmaZHIUT25bN5K3fQtYipYJkZNZbvaYVx+j0huBwYkz40RtExWsvhG+84hvrDsy2PThzQP4A4Pfkz6+FAFhgFdXB5p0FJLvaYABjU169KHY3n1eQiyEdgSMLFEktgSIAIpsKlaUATN4yT1UZaiDIIDlJIj6BapV82t759vsFGMAi05r86JeesGqDVrSi9QaAySnrDTDvcbNVEiUWdTauuDCr1a7bc4MmwFZvnxgmjZG9JUkRmAgLHAgWN+JxQyDJGQUQINbLxaq0SGbErgqAu3J5VO+FmWXDrcCytlzyRsY+6bQz3PtV6TZSRSByRVU9rmVPa6OAXvT4ZHLuFaYAdWyYqsJWhbMTJwegFbXVSFChfZizWtNbrzlPAVzaGH3TH2qw+tN2MoVz6LpRNvdFWn0kMdmMWHXpGtIdwrPEK2PgmzygNruRJJ8QexITz+ZJMk0FQdduveeeqzoqhuQI1fdtrzTgepPST5wn4GMkKrTJB71CPh+SS23ZNOYYmr0TNjMxbp/91KdV3QrpNa1Nh2TGTTrzxbI6KkpU24momLCd3X2r1mgXJYkxa8SARWScgxUksW521XTN4wCo5dMj1tjftpefe9o6DQcF1DIaNMm5HpEsAiK96oKxybVyDTLYkolSWi3srgfOuOvaSACwBjlTZd+Lzz1vg25f2r8FJdA5649AKrknSZyz3Ft1T0ghzSUhvOrZiSL9PZe1/eqeQClAAggG/vW/M2LooOkqeBFoITIDk3fMyNBqDOBLALoj7MhxCB5E/Am8DDqMIdCkU4GkUxszlZEyUsvZ1Mxhu/6WOy1dGRVRUUzlLDXoW73TsH3GQGgvZq7KYL3p89Iw9pb0U9Ma1Ya09xv1qtVrEBa71sFsrdXSOUFQIP1EVSBfBfSNCzmNE8AXGcam85IkQEogAkwR5B+SBkFfPI5hHx/BRD1FBW0At6KOeVg/Iqgo0B3fgnCfkqB0EnRLgvYQfnz52PJ7GkkOL3i9mqi4irQI5xfXLd45rBRO/Bzfo7Erubisgn866AR60g1DS6ykMrYDYMq195XwjBULdurESfuZD3zQaszNjNnf+ht/05bOXZTsDL1smMtGDdMhi5LYPuO9jpXffJbM6NWu7eekQJ09I4UJq1clkbBIzzZ4VsQ9TEFz6I64CtBMfGYS7I3P0sl2J5mGAKKzQ1ordf+AX+T/4FAs1/fmt9xnN9x4g6T3AMu19vd6qriHqAA4xKMCooL1m4PQUZGi+gnQOZBLSWIl/hw7KeJcj+fm509yFYkKEhknt3X9IswAZqiI3Q8t6AdA78GtCCRFIEmk45sAhA/GnAcJcZz7+VABfUBUJO91fJZJUjwJysZER88ewFBtPHwCwDng6Ij9/M//nN10623WsJxVqySGWXv68afs//61X7bnnnrYqnurqkoSUZGmc6ThFXjptN16623253/kxyxTnLZ0pmhPPPx5+6cf/IClrGk9SL/QUQHwVR4t2Pvf/1etVEQLv6y9DKCU+RXln0hcOW6nN7Bqk73Pq/WoZINcZm0jBiIxXF5ato9+9KN2+cplzfmFBSSlMjIzV9FEkOVS+3bQd3Yk2WO0+BXHgGs++/2P9ziSPMn1KDmXY0eo5mAgLuLf4z6RL1K04Am4E33uS6RkWmbjHiZABvGcAVIZc33riKiIklcki1Rbe7ctJPerxMav0lERSexOn30nEhWg2cmOCu/4jNeb/IQRy4Yqs4N5q3HFM+q7t4NZRtJPVPH7OKM2VLSAijFcTg+2Pq6zwTQ7UC6yC+Kpc59EvHqnCvfOuwu8w0gATNq9qTSmISpCp5Ji0UAsx3UwOScU0YgMdRpRZFb4TDqJvavCiyGuml/pjIoxKIrZ30MCcU/xBUD51URhuIboQaQuQY8l3ZSdZ+sRL8Q8a4jI+FxOoPV1112nIpYhUSFpqK6kn4g5AHEoAhBx0Ht1oiKEB5LdAWTGY+3ajor96q5RTIUnGoASY4QxyM8T3bLVaw2BSGtrG/I32dzcttHRks0eOiQPuuefe95OnzplK1eW7cYzZ9SBwOc99tiX7f4H3qox8MILLw6Lm+jKvPfeu+VzAXCxv1ezyui4nb+4qG6H2fkZEXtPPP6YvfObvsmatbpiGubAzuamFXIZ172u1+TP12zUbWy0ojzppXMXJGEn36VOxw4fOSwdePkzbG7ZqdOngm+XS5YgOzc5PS7Ndzw8SqWK7e5VbXtnT9fa7vZEQGxtbSmH4LPocMymB1Yp5O2mG05bo7or6SfmAdWiL567YIt0ZXQBnXKK8QD35ufmJfHKeUUgjU4T1ixfz1g/+gKGFH9DSOVzVsznVfSxubZq2XTKZqcnbe7QrF26cF5EDd03jz/5lFWmpu3Zl87ZIJuzucPHbWllQzK6c4fmbWV5SXsjpMN1119ny6sbIt7bnZY8DzUm+14QMTFaUUcxOaT+lk3ZpStL6iqk6+XC+Qt27NgJrcNcW6vr8lhUwhZLo+rsZZw3mhQ1ONCjjgkVlDmgx9pDPEweIfAySAlLlrVVtUG7anfddoPNVYp2ZHrCtlaXJfFbo+hqZMQqU5M2e/io7e7V7PMPf0H5yV133W2FsYq9/xNnX5m8fZWl8rV+Pf0rf8fyD9ymlyW7HKjUT00fgH7xOI2PflbSTxFMv1YuChmm8vf/kauO93rIkCSgn+wQoKtj+kN/S8eFFNj8wZ+2IUh/DaHwSq/9akRFsvOC4ye7FL5aV0VSOioSCrx/5t/+A8vddUbnunTD9+nfeL9eiVBYeObXRYzEexnfH7tHkrJP8Tls/vm/JwIlvvfaa3it5/61/v2mi79rOdbLbNHmpmZttDSqCnHWR7q+KsWsjfQaVq/u2s7+tu3ut2x2ftL2q3VbXt02S+UsUxi3UmXGnnvpvFkma+0B5C5kcE57k/YYSENA2CZd7sRNDRU4gEeAN2CmLQk+wl55vTiRwJdiWLqi3RhKBXn5dEZSUhyTfZscD+yEIlCIRcgGctQ6Ekv5nBsydzresRg6IVmnmPte4OVSVRwv+iF4J3xe2AWSTLFA16UMnVhwTMJ9LRQiQGaCoyiWcoUIkSJaH4m7yTm8+NXzGeHeLq+oa3G5bfXxdhy3oig0dhzENWmIMw299zxvo8ODoj/OXfX08gjxGEfyjJIDcm8GiB0wMAooVSCAzFYoUkQBwpCyyxTsxPHjtrqybsurq9YdSVl5ctL6qllBst1lLoWLqe7JC2DYh8kpYp7Bs4z5Gb9T/B3uY5RqirF+LKQaFuB0XWKT9z387w8k+O57T13PgWNFAki4WJDd8vgSM++u9l8Vb4aYRUXW4E8U+uIBImkmYqqOlcsF29/ZFU7HHj1eGRMRIs/QXMH2q1X17dJNQewBZsDeOTBM1um+y1p9f9eKuYGVISpuO2Ppbsvy+Kxitt5pWwfZ7v6IjWSLdnl9y7b26t6BjdoL3TS8ronPUt4yYbyksyM2f3TeXn75RRst0/VBAQTxQld73SDTF1mh2Nzwk3PlgDeIiq91NXzjdd8wdwCigoUG8oGK/yGo5amQAzuB+UUHFEkfgkEWg2g0BMhIosLCtLK6ZhOTk6oGkgFvjyDc9ftqNZhPtOISsiWSI0JGByMk15GjKaLXadj4aNGOLExbsZCxFm3r6YwtXlm2/kjWRrKjNkgVTNL96r9nwYRMATDnGCyOXnXLxihPB4LbnAO5XAukgACTWG0bjH2iqZLYaDd2CBVKvonKyDCAuIASSuiU1AUd5RQJKW2GdIm4dIrYcIzkaizmLg8jYIrzpEugVBIAyzlxbrTrseiw+EuHnPc2agoG+ByCdoATQGZMlQUO8Jw6XH/HcoW87jMssJhz2P8eHSjeGq+2xSBj5QSVS2UJlhYJlXYtbSqVeCCxSlObVUrXp8rM0AIdqwbb7YZAcTZ7JdHIWtDEJgmojsiK2+91zU5ttIkKf+5jJCo8SXaQ35Oi3lcQFXGD80Spb23a7iEqMNibmbbJyqh9/jN0VNRtbHzCpmdnVRWAjAFm2iTOVIiVyzkbSfVsfHLM9vcatld1QJ7nVpPWL0FNAP8hs4LsRTQdhyiTcfRI2lr1XTv/0tNWh2FXJ5J3VMQgx5ly96jw6g5PipDTKJdLAkx07TL9dpklKgLVvYNcA10buzv2wrPPaQ6WC0Ur0jZJAJjiOJji+v0QARW6oWTOK3AJnxQ303adaZ/nEBVIM+QKBZsYZ/46MAYwSBLa1tikApVELiOvDXVhiZxyCbVYFOZ602lJG8mfQsQfQJdrgvK56ioIpqjoL+uYo2NWLo/Z8dO32Kkzt1kK0DadtTQkHOBqs261Bi36ocJ8xGUbkBcRWNztWKcDUVEPXhR4UtTUUQEo26rti/BkflCpR/VhNNMuFiAq8gI3AV+YD/jtqHLwi4+p20kAoWzHQu1pABEjcJgEsmNHlgCq8BVu9bDymesQYdj3sUtwKzhIFTbewZEE4OLneLVO7KgI9z0CyqFi2HGvayqYhasH49dg9CZCKxidxfOP/w7JmMHARqmM3NlxA3d8R6hcCgbw65vr4d4Ii1P1KgTa1MSk/a2/+XcsPzFpo4dm7AM/84/syS88YiNaizuGa40A+bDHxEBVZz6sEI6+KK65OiTgGMdZ5NkCaIekEccCsQgkXKxk4n5FUNADfq9k9kTDkw0lTAHwHQLBYd1mzsS7qf1RmvH+eVeRF7xfOrvunXTvvffarbfdZqvrayIq8PjhnNZXVu3c2bPak0TkRqmuvstSpJGdkJzXAQAd18t4r5R4BAPsSK4PSXRJU0QA20HdSLByTAh3uikk6+d/9WcQQNw47pLk2FVAsDotAoAbjqAxGbR8I7DlXI6fR/I+DUHSyGgmoqWrCAwlqp5sRdIqnR7Y+9//V+w7v/uPWq1HGz5VSxl78PcftP/wb3/NLl14xur76wKaSYSJadS1GLoRASf/wo/8mOVG2QtK9uwTX7Zf+sDfcY8KOkWRmup7bFMeLYmoILZRsQM+Vp1WkBKcsNOnTksiRVJjvYFMYRlFtWpNySNkHrEIawxrOIa7n3voIZn2Qq69+d571Y14efGi9gIVUSADiWxURG2jtKAAYzcejJ0tiSVXdzBJsiXve7y9EcRW50YgKiJJKTI5dOPlICpCV6V77Pi+oTWNCR60dzud4AGWpVq+IMBWYwbCJ8hqAlyQ2IkUCOuPn0/oRBh2JB308kQjX8Bn9jBV7oWqw8AmOFkRC2nUbXQwzg7W2+BenRhf8ccufkbSLB6RoTYkOeNMnXlaC9x5RufJZwfiL5heDNc7P1cvPGH8UF3vq27Yb0kgQ7cSXIdI1iCB6u0HXq2p0w/zJcpBxPVJ5FnolNMzDxWSHoci2egEKLGVy0l4XMt8Zk+fnJoUoc+cjxJ4cS/yR+HdCv5MfB2IRIXiE4ExrLP+N42TIK02NT1l150+LSBX1yZ5qJQNej27BFGBsWaxYPmim16z1MUO0wje+HqATrOvK95pWtR+A1kR/VKIpet1L5YBSOK4ADsAyshYlOpU7tatXBq1J598Wvv40vKypNrecv9bFAv9zn/6HXvLW95iK1eW7N777hOQTWHCRz/2MXVEEP988dEv6lzo0O132/aOd75N99j35Yw1G207e/aczR8+bPNH5q1QzNmXH0f66a2i0ABDcvmC7W5uWKmQV/drVwUSDVWk0rWJB9jL585bgxwlSLIePrxgX37scTt2/Lg6AW5/05tsb3dXQAlVm8g9lDHCLhZEUMzMzql4a3l1zaamZ9WFe2VpWWQFndkQ9/mMWXrQt1I+Y7ecuc66zbpkdsk7Wp2u7TU6dnl5zdq9lO3s17TGsW7hRUHuASkS1wgKzYj7lE8BbPHYUvjJ5LWHFNT927FDs9O2tb4uI+2pyTGbnZq0C+fOqijt5KnTtrKxaXuNpl24vGytwYiNT81YJltiqVfOsrO97RXNNrD5+TlbvHzFCkj8qgCKtRwACOmOvo2VSuqoIE5VpbL17MLiJXVUIFN79uWX7cYbblIHBZItnmNRGd6yUarB8eCrN9xYV8VU7kfHfIpSaORkE+MTvqarO7onaRlePz6at15z32698YTNlvN2eGrcLl84p8pcSMnNvT1bOHbMxmdmJS34yKNflEH7kZPHbWtnx376yztfZ6Lipyz/gMs6JYmKV5N14jXIP0XSoHdl3boXlg9iVubt3Q7SR+mi/69ERQT548EjMRCJithlAKDfefLlq1bt3L03C/yPXQlfjaiIx0se4NrPeoUtYehRce37k2QL15AkGl7ps64lNpJkz97P/aplbzwheSdIDow5uS7ubefFi0OZqFeT0nql8349v7t/92ErF8qGcH4O1YAORYRg1B0rUTiXzduJw0U7cXTesoW0VaYnLVsZtY1LS7ayvmur6zu2s9ex8al5O39pBXZQPhZIFbvvZUZxsYyNlc+H3J2uBgBrCjHTGTt24rhLYnc7LhMUCEIVAOKxkEdhYl+7UqfZtl6ro/WD17Ef0kWH1yd7SKk4Kv8a5inyd6zTFO0B+rL/sFdFbxy6POi6OHfunJ04cVLzWjhHIBLUdZhDYiqjeEwm1flCiF8POliVhwRyQmVTfScqiBOjQTXEuLZXYvnwkPgc76Jw0kKdwkHtg5xZnkiSCHeP0gNZ6NywEx9sK4L84E8qWsXzVPE8HRJOvnAt7KMiaOp1yS6qsDgUrFJUxp4qUtZ6lh0M7OSxkyrMOfvyedutVm23XrfK1JSN5DIidUUQBEKJ9Zn9ktxGHS2x4zP4rIILxvwsEhicr+5ByNucYGHd9y4U/ubFm6iHdOzRD5eHw/vu79rTz+pCDsoiHvcckCXEURSs0rVPoZc2KGJphSWeu6ckf+ud7Ozv7FG72nOI2ZGiH9XzAUPb26uJrGctRwEBz1IvlihYsVCxbmcQZKP2rZAd2FhhxO6+/Yyle21LQ4wgYRj22nZvYIXKpC1v7NjS+ralcyX5Mw3UserPF9wH43ryFvb6WrPq/qK9gUsSZgrq4sDQm0K/kdyIdVpISrrMmZRN3uioeD1L4huv/Ua4A/M9N2eObWIsAJJ5Up7jIP5BEii3A2dho/lhqLilKilWUwIQbG5v2tjYhCYOADhJLT4TTLJ+D4kEOikcDCUPowrKPQ56VhqlXa+mILC+t24zk6N2y03XK/CmVeri5VV74pmztlcHuPXK96jzHIF8FjOSMxn6qj3QgXfAIhJLqoZkUhsW1yijEQGyCLxHrWgS7aiNF0F0iAcZ9Sl5VArpANuAdsfCEADk2NLiQ7dVYIQnm9HcG5AymwMkxQwwb1vb23otiz9J1n51XwC2M/RU2AP4kyxQJQpTnpEREC1rvI6NBnKIgBySgiSORRCtXTYPETVilj1hUZWtzKKcGeeeqJMigCKc687urhZwLnZne1dBADst2pNa/CURRrIgTlst2lEGCnILM0OXfurabcFM2z/HpVwiKBZlnuI9ZkNLEhVcR2wNTG52Q6ICX4x+z+bnDsmj4tHPP+xExdiETc1S/UalBETFvOUKRUkWoEOcSrdtbILqkpbt7gPIQ1R05R3CdhcrWmMXAueHVwKGq70RzLezlhvJWbdZs8ULz9jOyhVVgbjXhwdrjEk6U/hcxnGsOEhKWBHccG95jpIayBcU7KlyAF3LQVfm4BgOoqtYyrFh0omQUdUDARb3B/KLcYkUmEuTYG3oIANeKYBnDtUijUD1eU1VjIVy2SbGp0L1BM/FOzHYrAkmCLoyqaySYaTBKJGEtPJD+TiIHTrIVqFHypfWlCBvwusb1ZrWBjSnV1aWDd8QJDgOHVqwm+96mx09eaPGNpu8CKxW2/0oqKrLekcIa5Mb5QaiosNrGqqOQ2eZ80NyAMNvgrZmbU/BCMdB9onvOIYiUcHzmZ2d1T0DhLz+huvtiaeetS8+9lgAS6MElAfjHoh+JUiWXPvj2OZ3sZvFJVu824U1Q2tDCAD99Q7yqnovIeOkAPkaWScRTsGoMoLS/jgCAB1OhuBdgBD6p2BfPE8ITD1jD1ivJSni59G9BQhEpeD4xIQ0tVU5lc3axvaGP/thtW1K44494Yd/8Ift5K23W79UtM986v9l7z2ALM/O677v5djhdfd0T0/eMLM5YLEIi7TAIoqkKFCpLFbZli3JlERBJCRLlsyibYmSLFl2lcxi2bRZFmnKlkuUVAIJAiSRsYuwi815ZndST+4cX06u3/nuff2fxuwiFGgFb9duTU9Pv/f+4f7v/e455zvnMfud/+dfWLZPqGvb1HsVAdlAEuiaBkAzKoQ5hmj35jZ+uySfA39OZjJONDdEcJdiF8/ZcG15bbwmtJKPxmxQNqsvIkH4RBVTEqRPXqM4b8Xfi/c8FtFvf/vb7V3vfrcyZRh/2OZxDJcvXJSdBgU1HqSeKQK4C1HBc+/2SSHMaQT2J1XQ8bOZI3x92w23dkAx2DSFMGRXWmUFwNabZLdsO6gG8RoOnOuKYn7UfZGYl5NknAC7lCvFA82htTXaeO0FzJPXjI+KxxotYN7oWaE7T2q7ABBynfBB/2N/7MftZz/1V2yng7qpb83GwD7/O5+zL/7eb9vVy69Zc2dFaxdjgeeZz+F5ZhwcPHTY/tJf/bQVxufNMhU7c/Jl+5/+3i9Yut9UGDRDhzWKJ5o65ud/7udtsjapeZgfIn6AWGVjeOL4bVYjRweSXxkDDuju1Ot6nhkH3G+6D2klX11ZtRdffNG+8tWvqDa5/777tCk+c+qUQFfmuGhNp/lNgcaI+XdJyzh+IxERn3NtNhNdFz6z+5wcfyfOdRIohDDteA/ixleb9CJEWewm8Hkk1kfYsVA3MAdR06ECUycqvswiyT3AnA+Xt3O/rzlaysFQH8X5LHnfk2PbgfyBLHD0zOLOkrA+G81rIsFY2wJBssfSLnY7xM9Jfi7kOvUUl2dmdlY1pAAO77cYeUc7WImK20lSXkDmdrz+EXTn7yI+tNTyXPg8xmv9OYnTTcgyC+R9zNnyYEfvTExeCz136Tgvh46KULdqww9Q0abWcgDVA799wy+BRTZr4xNuwcgzfx0ZG7pBnJhEAUuXs485v6Za3XTg8Vrxu16XFGx8vGoTk1W7+eZblElDGQDxLNus/sAuLyzIToGxTZ4aYytJVCTHbpwXeNZ5b2pfBBnKiyC7IZsLlpF1zXdJooIuTNaniW5Vnuidds+efuYZO3jokMDpmZlZu/POO3Qtvv7Vr9o73/EOW11ZsXvvvddefvklq9Wm7PHHv2MfePhheZ0//u0nrFDETjMrC6OPfORD6uBYW10TGEYnw/rGhkHSyHqqlLVnn33aPvjhR2CBpfylq6HXadvhozfZwpnTtnTlqkQT5CQcPXrY7nrnu+zMiy8pg29+/37NTYgkzp07Z2Nj47a2umpHjx11GycJmrzrtd1pyoYC4c3Y+Lh1On17/fQZmztwQPZz7WAh2ey0bWdrS2RBuZi1Ui5tD9xzp6UGXbBRdfVub+7YteV1+84zL9j+Q0dsY6shYQjAF0SFyNNe31479ZrmQO4d+xOyY5inTp163Wo1wsU37Pitt9j62or1IWAfuF8kFWAQXc0d6kSEXSnT/NseDG0HW4xU2pq9geynqMlLxbItLy4ruNtzqDyoe5UOkUxe+x3AS3YYZGGU8PYeDmX/xH6OjDb4QQLGsb2FhMQa69ZbT+i+bW9hrUuunHcIIVhCJLJJZyEgq2xaHWz0pnu3S2Hs19iHbW9rDKlel39+24o5nJ827N7bb7G58ZLdeuSwXT572hr42NOJUa3YzXfcYcN8wZaXluzLX33MLDOw97z3fVaslO2vfe1i0PeEh3E0U9yAxf8+/i0JikdLJV4GeJ6Zm/Z6tZAbdVcAiPNVDbkWyTl57/cRlP/DIiq+V0aE5qEQEP7DEhW9s1ds6eN/9Yan+UZkxl6iInn+e3MreOO9v8/P4nvT0ZG96aCCuumaSGEZdMcx47h65y7LUguLqqt3/Zk3uxU/9L/dt/h1m56YsonyuB0+cMTymbydfv2sHT58UATm+dOnLD3s2P59k9bqNqxYLWmepNt0ZXWLZFFrd7O20xzYlaUN28G+Ws4J4Ds4EWDvzXrp4DzzMV877NOoOyAb8kUrV8vqhMB6eW19TV1R2AmJiGQvA1EAaIwAlg7+Ykl7FuYfhJQQuHRzMQciEuGLmqQcSFpyTYVlURuHTIIOQr9eX5aC0zMz1mcfFDIOOFbECnyBnTie4cIQjps6pFKGLPasSNVSKY6H1/i+ygUmbhXF+fP7EL2jtTN0Mnit5ZbksXOC2o8v1kheA+GgbsEw3zB/cV1lQ6y8VAf4vePR12i5cbBflJ0dNol1P3eJHbtWyJckKiQ4GlKKtRkynm5HVv5BuyWrzqmZGc2T242m1ekyKJVsrDZpDYD8IJKjWwGyOu5f3XapGrob/Nij3apcVUQW7To5SHgUKdogguW9qBX5inPwk7+9S1S845N1v8+EVRdx9WiP6kLmbQmS6JJBFIxoeIBg1q04gyEjHAAAIABJREFU2wisg9CNbbDcTen+SQ+UK3Tl8hUJ7KjTsVlkXFHnb27uSLSJQJIOvZ3GtrW7kPcpy6TyVsiVrdNsWK/TtFKOjoqh3XvHzZYZdKyYS1lFxNiOXr9db1kqU7B1upNWtq3dM5Eh2WLJKtVxK5f9+nHcV69ctp1m00rVooQNEIlYcnc7fWt1e1Yam8AFytK4mSBuboPPkAX7VkbFDz05vvXCf3evwEzwR+O59U4Htiq+EVMWhWxdvD1P4AchqEFdJSW+LCVSAlYpsJdXlqVU1wQWQAlaprSRFRmBershX7U4wUbrYjaA6oyAvcyn1FY7VjC7+85b7P5771CexTCTs+dfeNWefPYV61rGmh3UfrnQmu6TmDon6CQghClsEiMARsGvLoegzIkgY2yZ86583xBGxayDBg5C8P5xI8WEyKLp18xBRVegBd/y0CbHe3sA0mBElHB9FHANu5sBYCtpQhRwlPHNGhO81FYo+AORwHtht8PGzD2Nh2oLY1E4OD/vIUyplGyaWNRo9ZOSQWFTKYUaUhBwjBA/sPcO4A0ErmBXFUF1foeAHwp+FihNiMEHng2d2igVah2CMglmElFAkUDR4h01fN8buOUWm+ho/eSdPIByu0BDJCb2EhUO+LR1HnuJChFkhtqVIC5vQ52bnbVKIWfPPvm0FuaJiZrC7QB02RTtn5+3XLEoooLrkMl2bKIGUdFNEBUeuBfDy1UoB7ukSFSkMtAyZFrkRVSk+h27fOFVW7p03grBjoYCIpIyKBIK+FsSgB3OPQnYMR4prlC28Bz5/XD7Dd6j2SUIesteP/WatRtNERUshoyHPrY7RZSLHgTFmARYVncMwYCo3gjgDgUBNj4MBOyRuD8UkGyepianRT7QeePEnXdAUNjJciaDx3FFBICsr1A9u7dUsCXz+8r7e/ig+2dqtAZwhUITuzbmmK2tDdvZblo+X7b984ftgYc+bNNzR0YK30geoszFBk4YkKxhBnpGIlGBeqHTRgVITkVDfskE6SpUu74jOy5UjdH2iT8jMFQsuH0dwCa2Ljx/FMl33nWXNdpd+4MvfNEuXbo0Clh1H/5de50IviZBpjjrx/F9PdjmKuXYJSAyKxRVXsh68XmjjgoK8iRwfD1R4dhkBIeTr99LVGjexZ4K+Dp2CoS5T6B1UL2wAOBFvbKyrHkKoGJzdU3jsVyp2OrGihTj6poJxyxFSj5vf+wnP2kPfOBhW9zZsdXFNfut3/gN62yv26Df8jmbaxi+IikTSRN+HMkaFa4qxp20i78b1Tn8yZhjbqBY49ryd86BeUP2GmQvhfOLICZXWU6uAIQB3N8LtPP3vUROvK5JEimeR1Tw33ffffbwBz9ol69cVisxSnuOZeHsWVtaXHKiIqj4te706fhz5THAKK3K8Rr4erwLZvj33u0WuyuuA4BHhIvbMGm8sr4oN4WcFmzQOgrmjeu9nk8C0cM6FpXgyfE7AsqDpU0kKtSFGMDk70VUxM1Z8j4njz3WBV5/uJIbwJfaIJdL2YMPvs3+u1/6u9YeFK1e79vqyo599jO/Y48/9hW7fPGkteprrozN5ZRzEI+Ha88G9VOf/puWH99v6fy4XTrzuv0Pf/dvW7+9pbVD/UXMZ9jBlUr2qU99yvbtmwnrs/vpkzHBhuH48eO2b99csPYB/PJuB8gM5iDGAXM3a//Wxqau98mTJ+3zv/d5jUXu24EDB2zQ7WqTyyaN/+PY0rhjRt3TXTWqmxJjIpIJyUozSRCpJgm1ipSAbGxCmHacXwUIQzRE24OwsUs+hz7l+fMHKsjaxvnKFzgIHNQBGgMUu93QUfHmRMXesc3rmX+5Hqpp9mS06Br80ESFPzvqBByaFOxkL0MwoWjDx9hzHxyDoAsYUc1oLg1B53HuGakbIQoy1ECx28iJCrea8Dk7ec09T83vWMYX+NHvxHnqexEV6iDGU1+kEJtyN66KRAVvL2Up9V3XbSa8S8SBUP/TM0jysvAK1nGBLI4qx3h/uAbMT6j6JybGbHwCouJmdZCweYd4VvUsouKCcqN4jvKlnMQ48qgOdXSsB+J7+3rqIIWsRre3Re5xPalFqD/rdFTsISpkP5bL2kRvTGA6qnlAdPYjKyursvm8+547VIc88fjjdt+99+p5u/X4cTt7+rQ+68tf+Zq9933vU/fIs889p/terZRt0O/afffepTyCKATCOnTh/AWb3jdtc/tnpTx++qnv2Afe915bXly08YkxO3XylCyfAPzXV9cEdNd3tm3f/nl74Zln7B3veKeU/KyncV1CbKQwWe4VApnBUOsrBBPHg1AF642lxUV724MP2jPPPC+ykPWODuFMvmAXrl6x6hg2UA5CAT5WAaIyQ7vnjltt0MZWxJQDSJjn2mbdXjp51mozc7a+Wdfr2DcA1sjuMliyaN7b3LQD8wcEgPG5iGpUG/Y6NjE2Jj9u7J5q42MK0iaQZKJasY2VVR0He67jd99jL7/0qhXGxuzchUsK0251GbMAbGb9jneEM4YBFucPHJD9l6L16O5GuY2PfCFvBeaIclmkRey0QYX68slTApXI8lhaWpL1007YcyL6wbecvRZ2HCqBMlnZolGvtJpuUSMbvtA9zjyDuAfSjLEssCzsM7IpLFPq9o777rCJfMYOTI1bFaV4s2lXry3ZIJOx4ljVanNzllKId9uFITyr6Yz93JfP/Ug7KpI5D29kH7SXaOidu2KT//1f1nlBBCQ7KpLrCZkPW//4/7I/LKIiaafU2dNREY9jsLJh63/9f37TMO3/LzsqbmQldSOiYvYPflnkBNc3mWFBhgbWWpAT/UvL+p03I1OS9+OH+f7ea1+zHLVUL2MH2COXq9ZudpS9sH9u2qYnK1Ytpq3XwWanbWtbmzY+NWk7m3VbWtmyZotupJR1B9QJYwoJbrQ71h0yzyP+DDUpIgs6/4YmUpiJPQuoynPT69vs/v2aJ1Hp0+VAlz+1KAQluAYYEB2VYDCIzcbLFQmsqKtYp6mdICUkElIQMZ39Zr1gkQjpAMZULhfdKSKBMVy6dNnGx8asUh1TfQahINV8z0VQrCXUx3QG8vla3zmfUH+7I4eTF4jt+ILIdoGS73N5ve9R3I7HawC30XUxsAtnWJu115K9twsDUc7HWjreYxeDgA34npz3jySBr6MuKIyWzd5l4Q4psZbANhzMim5H8BKQKnUWQM40GjYzMWHLyysBkG/a+taWtQg5L5WsOkEWCeHRZHiUJcrg86mpWT/Zm7P3ivssfkbtxrgCJ4r1oFtlRUIFfGiX7JCTRyB6vJNkaM99rjYa5g/80U2RLrwf9YecQ/J0IjjJzHthLSZcQwIsz9RVJ4XssFT1WXqYUuYJ6xOZLJD4fN7mxrpIAeZ5SBewCzKNGLcQ9lzbdrdpzU5DdV2n2bex8pjq90592/Lpno1XsnbP7TfpfVl3jxw7YuSXprBIoyO02bWNrR3b2Kpbvdmyra2GwbOBVUIOHZzfb7XJcds3M2WIDRiXq+vrEquur5JJm7PeICXbKMvlrS2SJxfExm4P/1ZHxQ8zM771mn+nr8As6fG0uSpTzHdNahmWBY1yknwyHg7EvPIAa+KmvVtWSnl5wY1Vx1TgMdGhJqJd2TMUAFLwcyNcuiulPSHTse0tgjpMlq66c+gop4Cflo2XhjZeytnb33aHHmBUKtdWNuz0+cu2ulm39a2WDYa0HbJY4KOOut0ndCYwAFIWKp+0HYTxbgIPY2Zl8MnOg6+jWplfdj9CB1/ZHGnCC5t7KQcyWbXCsYixWeS91FbH7wXQi9fHwG35/KurAkWxbxLVRo96SLZMnifBNQE0jUFPTLa0OUYlo1j+Pn55viiK3Q7ABxZQLHRi1VEI0rpY8s0Qtg0sdlwPVwhyWwdSRaJOcLDMQWaBBAQly8ol7+11wXeR68r9BHiR3VYgsQjSBbiGnED9pA6ZFCA9RQDXh8KlZ3fc/zZdKzbZSeunCI5GMoBrw/dcj0hU8GeSqGAhdrAXMRtEBRunrs3vn7NiNmPPP/2sNh8TE1NWm5kKREXO5ubn1dmwb2aflArZfFdERX2nb9t17LzowOlqzLJhiwttVD+PiIp033qpjmVSBctb3lKDji1ePW2Xz75medSB6oRxRS/HKluDStVyheJ3nXssKuJ4ARCAqFBmhXzgsaUYyMbo9GunrYklQK4gX2AICorA6ji/7yA+zwGtsvpsT8x1ZfrQdE1iMDL+1fyzwp1zOavVZtTaHi212JZxz71YQt1YUD4BYe4A3THo1n3V3StUGTQDCioPukqqfXnuyDXIZnlOKc6k/bRMmvOdsHvf8bBVa3N6hvlCPcFvEOZYLBc1H3GtGPOjjgrAt27HWs0da2P91GpYq9EQURE7KtqoIdotdVKwgY1AvBQq2bRNTGA9VZFlBOMSW7A777pTQZOvvX7aPve5zymsk2shBaoAXSdqIxgaW3UjuJdUuscx5ECN230lQd34Wi+sfdkQ8ZkgJvSMJMgEFamyGuL68bvX2+y8GVGhopBNQSAqknNbErzUHBOKXgAePW9C8czGJydsc3tDBCw/pwCMaiqu4Uc/9gl73x/5I7bcbNilhSv2hc98xlYvLthw0JYCHRI0+RUBtBiCnRw7IndD54eeh0AaxusaAXvNLZqz/ZmLRKAU7oGsQFml65ogKiIgLOI5bFCS3yc/O0mUxHsdzyMqpU6cOGGPfPjDtrK6ouIX8pi5/PVTp6TOVRdYh5ybQC4NaGum443A+5AHkLCj2ltI7ALGzNHXX5to0cL70CYfbUuUbwLRNxwKAIM8URZGDIvXGhHuYRiESaJC5yqgkznJQU657rv03En7ACrHcZsEzDVeg5VPnO/j78XzSxIVThxEKx3mz6wdOXLI/skv/xMb5iZsp963yxeX7fd+93P21OOP2aWFk9ZurGq94n1QRsUNG11m5eqYffpv/m0r1w5arlizy+fP2P/4S79gncZ6yF9g7fQWejaRP/uX/7LN7Z+T9Upcb6ltAC0PHDhoBw8e1rXQc4olCQKC4VD328ldwr57AsI4CzrhPvu7n9Vmi98T8Z/IC4rPnQPx7gucvK5JkiKSV0kQOTlG4nvF6x8B9b1EBa+JXUEKq8dfOufWYnGc676K/Nvt3BkOY7eX11Jc32gRSX0BkMk1UPBhoqPiuwtiXzfiF8cronh8XMrJkYAmYRP3wxAVu+OKEehZWtRdR44ds7HxSbt48bI6LlFKq0MXRFHPn+djxHkm1m4uigmiFupKyA3VQLu2aE5w7BIVUYihOTVk7CjvLQAIcd75/okKckDo3nHrmiRRIe9rnoPQlaenNXSseQOHH7syZbI52Q34WMbiywEa7luc9+KzjaVOJCqmpibswMFDyp5gYulzHozZ3sAuLSzgg+TiCSxkIJvfkKhw6x6Oi+vCOowIgbWa6yklLV7ndVTtTlyUylhEYZOR03NX640rtBUI5tTJ15TjAIBFN+29995lw2HXnnrqKbvnnrtsZXnJ7rjtdjtP8HKpbI8+9g378Ic/qrnsiSe+I9sgaqetzQ173/vfYzkCsOkClZVnSq+bnZu1Q4fmVeO+9NLz9t73vNu21tZ0vuur6/bqK6+qK6tUKKle4vkojU/a+tKijY+N65qzDlB3yDIl65Za3gnuJBm1tdu/FkWi0jnAOgIBm8nlBeKnALuGKSlgVzYQgBRl2+Hd3kMr5FI2VinYiZsOWzbU4xAgdcCSVs9eee2cFcrjtri8boVySYremZlpnSsh0+zpqtUxHRDXhevFPm5hYUG1EhZ5EAdZwLx+zybHxmxjbcVS/Z5VyBGhcxbrTBvaTTffYt968hnbd/CQvXLqdRsw1kQOAtD1rVou26BHl8OWFM4zs/tsbXVdVrg7zbquLXsJnhf+n6lN6jWMe+YtituLVy7reSbIlzrv5puPW6NBxqHbn9D1g5WHTNeCxSvzM3MO54uYRx3HslB0cQ9rCOMxzpOpbEpiGLpVCNO++8Qxm5+s2lS5aDmGf7stFW0aMdTBQzbM50T0DCAEqcH7PWv1++qo8HV0b0fFd8+S3+9PRoD/G4RH34hoeKN8Bj6TjAjyE+LXHxZREe2pYpbD3vNNHscP0lHxvaya4ud8vx0V/P6bXa94HsnOiGRYuR7tRNfE3k6SG3VpfL/3/nv93jvWv2UT1XGbKI9ZMV+UMmV1Zd0yqayNjxesUsjY1HhJ47pcKdrkzLRVJ6dsc23dWu2+ra43bGmlbu1uWhbJDQDWbkeer5GIFx5BRoHEaSl1RKnGQKZIJmk2K1s7/oR4ZF6kuxv8yS3psBd3y2StWQOzHvsLcmo6beElW9t1dQryJXIinDjdFfy79uedjr6PndSsK+xftra3NJ8xpwoTCpZLzMnMEXTsy6ZY62cU7fpaypwq67uenx97MWEvek3MtvFsL+/yDh2JYd8ShQGyc07T7eDZf07qILCF/PUO6+R+A3KHekq4kwgCrAh93uDfWA85z9gVpjxK2VD5caoDtt0RtgeQDzHBcpuHCKrvWDmXtwOzc1pLyQd57fQZ2yCLgT04tRzzWqFo241tK1WrqnXAmmKnslte7WaMRByJayZrL2pJOtkiARywnXiOyT0Hr417tuc/v0tUvP0nt0ZEDVhPFFxEbEH7iWBiyXjBphhyXPtMkV8+9uj1odyU1GbQttmpCbty5VII327ZvpkZ/R6169Wri5qvEZExZsiE2Kpvqvu03+7ZWKlqtbExKxcylh20bWdjyQ4fnLHaeFXvf+ToYctXSgJS6WJkTZLwCsIJEYDyVehOJtycjh/2qA3PE5UdKTkmA+WMbKxv26WLV63ZGVirm7JGd2jZ4pjuj7C+kAn7FlHxvWbBt/7937srMNOFnc4JdK6UKtownrj1uDz+Zf8jD8Ed6/exIipqE8MDTPEN0EVRixKIyZYCFjAUoO2ll1+11bVVAQMsKoCXTHCsPEziLqZNaSNBActmDUaVRa7d7luBAO523Y4cqNmw17C777jFxqtV22TDn85bp59Sq/Kla8u2vdOxeoMJ2fMn8BIVAKVNRU+Ts9p98cGDzc1mBBgJxPNufv+9MNmyIQVIlOdpyHWIf46Aw+DhHEkFFhhvbQd8ghQgZ8CzHQSohc6OCLxLWTdwZjmG0iqsTZ/nZAdgmr/MFzv8YQEEUZoVCQ+cqils7tGvPyrwWbZNBDqRb0C3R1A5Y4Ukz+3xqi0uLYmUiJZWHMfBgwelemAMsKhxjrS2Q5ZEZSrv22p73gDgO4QEijCx2+WirLt6IiewoRmqoICw4BJ3+7TjQyih+uvabfffr3PkmooACoAYP+N6JlXTcWMfmXqpEEIgNN/z5W2FIcMh5f6501M1m6xU7KnHnxCwPDm5S1RgMzQ7v9+y+YLNzc25PVK+a5O1qm3XCf8EKAbcd7uyeJ/4rKgG4Bqx6RmkejbMkCGRtwIdFcOuLV6GqDhlqZ5bW0mlAYiLrzwZKaimCyWp5SKoNwIK2eTI3sZBZ4BLdXLKfz9FpqAImfNnz9nq0rIVs3TFoMLOCSSh00GFsIgKt36CNEC9pXyKQkFFIc+be4nSfbMpYAalRKFcthIepiIknADi2ZDqr0+hllMLqdo0aXk0b62MoGm0O6lWKjYIqpN4bhrXAZQjQJ7xUShkbXV12bLZoo2P1Wx27qCduPtdVhqj+8XbWlFlSP0NqJfHZsU7VCgQFezYISujK4Ki3SILgND1pkgKuiqwtSIEt99uyqaAzSubxjjOOMd8LqMgbQAS7BaYC+isoKMCSwVUeL/5z35TrczR8obq2ME7B7EiYKgnNgK/iRVBYyZ0KfA65tL4FUGv+D6oIfe+T3zPWJSP/p5Q2vv77YL/Ecz0CTGoaIP1kzqrUPcF9WwENDV+wnv6POVKII2x0GILSEDhiTVDp98WeMLcEa3GpOTN5+2Rj33cPvrJT9qF1TVbXlq1L/ybz9jCyZctk+qHgHInfN4I1I7g2N5rEa+jiN4A0kvtCxjmiNxoXkkuyvyuxmi7o02L7K/i+QbLqBtd1zhHJe9X/D5et+Q95/sjR47YJz7xCSliyESBGMDP9dSrJ/U9cyXzoSZvR6VHZLUC/PZ0VCSPITlvJMmoMGh0Td3/NRTlWgudKMY+TjaKdDdubanjTGskBb34zN128nhOyc+Q8kvkhNuXeeiwbwbi78cNSQRe95JtybGWvD+jLh6RdNquefaTlOk8b0MbH6/Y//Kr/6uVJvZbozm0hXPX7Ctf/JKIirOnX5D1U2wrZ3zGawX4xPj49N/4r23m0HHr9PO2vbZi/+Tv/6LtbC/q2YTI4TMjePSzP/tXbG5uVvYwvi4TlNi1tdUN2TLeestxbRp9Q5fS/A65vL6+JpUZX7v2dEM7f+6ciAoA2FhLDEMtEjf6kbDUtaM2SlzXkTJtT34NnxNfl3xm4kbwOtICklGWJrv/x3UU0YW6DiErwnzNn/F/UIM4PlDQx7HgVgaelRDvLeOPz4C0AUhXzae8Bu/QTBIHu3MOG3EyCPICY5euXRPwHO9hnN+8EQBSjA67N7Z+So6z3ecHlSFr/FAiE8DTW0+csKefesYarVbIUXLRDHUgADyikXjtk89C3FDrvdOAJtQ/HJeTpDFMO75mL1Ghew4goyD13dDvSCL48xw6VsODwn0ekX/Mz13vpmANV16FOpF8lYh2bHwfARAJFETm7q4UABReN2KVkdE8oHMTELJrXcl9KRbLNjZG7WJ27KYj6rbzsPGMQfFpHugP7cqFC9brtq2A9VMhp8yqjALaff3mHKiLqTH5O/WGvM2zGa3BrO0Cd9Vh6CQGVpHU5cpBCmHaiAcgMsY7Vdverms+OnXytI1PTtr62oZCr++9907Dk/uxRx+1Bx98wJqtut16+x12/tQpXaPHH3/SPvjBDynLAKICmwXy3ra3NuyRRx5WBgJ2kp5rl5al0P75OTt60xHLF3P20vPP2Dvffr+IDayoymNVZRG1sNDY9nwi5hC6sQD7sTrhmC9dvGS33Xab6hLmY5F9Zra2uuJdwZWKamx90TUYAs65c9TfWEC9fvqsTU7PWKFUsdfOnrMSe66dHZucnrZ6fcsyqaFNjhXt0Py01SaqhqCohU1sqWyb2y178ZXTlslXbLvRVvAn1398HGICZXBbezfAeu4H/zY7M6v5FbuMsfGqjhVwh9kK//Kbjh2xa5cv2Tj17bBv25sbdujAvEKy77r7HvvqNx63mfl5O3XmrBUqFRumMra6tinv/B7WFu0QeGtmh8hyWFnXWoNIBytb6pBxQrzpPBYRj10VAeNldWJcunrVbUyLruqdmZnTc0xIOhZl+ORDVqhTPHQYuV2pd4jFTpFIH0QRGPMbeyw9e5pvAcPMUt2mPXDPCTtQG7fJUt5Wr121makp29xpWHswsPmjR2yzXrcKpHmlLNvTFoK9btf+1reWksvfj+T7JChO5sTGL/7qdURDUvEfsxCSGRbJfATIgdo//qs22Kzb5t/7P/Q+3z9RkbLp//O/GWVmfK+MiuRxtb/5gq3+2b87uh4EbWdma7bz65+1nf/tM2/aUTFY3bT1v/HLo3OO3Qy8GRkRvP5GXz8IURGDv/e+ZzK4O+Zp8Dt7A7ST/5Y8Pn43GTr+IxkQiTe59dwfWClftKmxqh2YO6B1anlxxe66+y4br5Ss367b8tXLduXiupUradt/qCahBgTA6tq2NVpD7ZEbTbPtZl8ALOQ0qCz7+d19IHsyX6fAY7T3ke0T3W85O3L0qJ69UgVBZkZrGOsg2AL1FfVBoVSSXWq/3bHa2ITs1MCZRBIoRwJcx23Eo90r7h08nNHyp8I5CfdxfAcbbfaSgM5a27DRKZVFTDIVYFdLDgG1itZL7fFcnBE7tON+BcwHTIR5gt/VPmToQkLqBdYnFwu4w4ZsIxO1tab00BHiGQ3+eb5WO26kLnERqBDwvl47AeEiGGrj3do62FcmOvLZt/HvyknVHmOgfB/EDcVcRnXg1ua6HZ6ft6II/5Itrq2K6EbpXyiWbYu9+mBg47UJ29jetvJ4RYJGcD7uHfUB+4coDtorJotkCXjcqFMt7PmSIhvGThT3KMg6l7Nv/yvvpOfr/h9f19zs4kcX0ng4umeUgWOS+UTnSJnjkU2Xd8NIc4JINxBiuUzOOnSlDHt2cG7aLixcEOkD+cUaR32O2wYZUKwJjGHI8manaa1OU/e3jAtKb2CTlZLdfutR67W2rZAl96Jls9PTuleM9Wa/a9WJMa3ldJUOOS4Jff08ZGkrIiMjGymy3px2YI3xICjWLepgMjGGlrP1rbY9/vRLdmlxzQZ0SFE75dISDr5FVPyoZ8233u/f+hXYP2xLzUPIM62ytAGi6Hn7A/dZbXJCCkYUZun0QJYxUlsRcIStAUD6MGVTk1Nqk2LTSltdbWpKICxZC8+/8JLYQyY2JnXYTcgJNsKuKPT30WSTcmIgmwNMpeuhb+16044enrUPfuBBK5XydvnSFVnU5AoVa3cHdvHSNbt0ZUmt+3iQMomhugGAkm80fnSZjApudUgw+WtSdfCNr7iBHXVQBOIiMrVJEDIJSql7gfazgneV0MLoLWh9zwhI0xmCL3hwKZBCClAX7NODtb2NraQFmk0m3/PvLJ5sClH4MGkDbNIGP9q0pVJSGNEGOTc7p0WDzVDc0EmZBtiQzmrRFuiQQQWxrfBAPpdj39rasUlaMBsNKerBzMTyd2gHHRPoz3hgMxDbDnkflLgA3VL/ZlxRSYC27JlT+DriuY8ysaMAUvQUhAGymb7tvvsD8+9ETdzE8yfv82ZEhY4FVUBgvLl/AlFUsJChQtBdJCrK9tQTTwrQpqNiamZa7YupNB0VTlSwGOncchAVFdvacaKCdjpUlw08uBMdFZGoENGyh6jIDjMKUFpbPm8Lr79qw7Z7UMbiLVrTZOnD8pvIAAAgAElEQVSAKFW0cHE/4zUYgXyoTgRie+i6L1auRGZNYmFbvHrNLi1csKyl9VwyBlO5tBR8AglDUcMY5T7BugMUyHe43fHgpdAhtL3tHRVsziu0xFbGPKNC9h0O6kD2OGiTsmKhrOvPhpJWUMYZ8wLPVAS/KoQ/BrsdVz7s5jOoOJGCpGfLy4u2uHjN8vmSHTp41I4fv8OOnLjfskXUMu4TKhIsjmEAlBAaKnXM1pZ12ExjP9LCbqUplTrFKJZPbAohKmiV3dlcs9XVFY1nB8+8JZhzLBUBxjw0l7ZVOscg8O64807NM6gb/umv/7qAB+YSB5b9nFDZREJKKqA3AMkjECkgUeNi17s8EhURvJQSJKl0T5AfsSBMzl27oN93LykjEkAf5x7rBIopozUQFfHzk0CzfjuGWicKdxVgjE82GoAD6YG6XZjraOF2JRVzWMk+9OGP2ns/9nFbrO/Y8tKaPfb7v2/nXnnJep16yDZxEJKvEXCbIF4iKJr8t2RxG8HD+BwpoF7KSidr4vHH6zO6B1hpkAnQdLJCc3wAPJPX9Y0W6CQptffaxXM5eOig/diP/bitb0BUbEgdDiF8+rXXNFerE41yNBAVlKdu5eTrrEDPRMv6dUSFvOudIBiR54kOCEhyV2yHAHh12vAaHj1AWOp2V/QQsivSUiD1d5MUSeDbr833R1TE+3ojIide1+SmJt6v+G9qmR6RONghshEkqDZj//uv/ZpNzh6xre2enT97xR7/5rfsiW98zV4/+bS1m+uhW2fom4Ngdafcp3LFPvXX/ys7dMs9yqjYWl2yX/lHf8dWli46iaNuCu9GY77983/uzxv3cQYgEM/gPLYALVtaWrFqGdubWx30DVZEvAaAnS+UyNxj5gs2TdwLskl+57O/Y+fPnx+tDfi6cy/4EjEYshP8ff0ZjePgexEVyfES3y9e/xFpcQOigtcJKGZTHkQWce3Sv0EWMUZCBoMTUB4IqRFG14DAZweg3VbI6yNEDwp6DERFfHaSREXMmuGYeYaZhwHAFxcXpSbj8+K5x/nMu4YKuj7xGUg+r74x3wX/k8/1cNiRDSW5YLfdfruCkS9evGhnzp131T9rQ8hrcMtn5ilfy6NdqMZr6CwbERVo+rRxdtsHmYLqtd6hEIkKziHmp/A9gceaj8Px/uBEhQs8ID6TRIWrVF0sMVpPApkAWDt61ugY0fl5pxS/2yVbLNhV8We8L9SmytLKZ+34iVuCn7QTFYBW2loPhrJ+gqigrswVsgJYqEcjUaFaVoIMt2sddQjnclo7AJkheOPczrUWUYH1Uy476qiAGKDmr/XHrdej83doTz39jGzZVtc2pPq/667bbbI2Zo89+nW7++47JY44fvxWu3TxopS1Tzz+pL33/R9Q9xOkBWSjOoZ7HfvYRz8sEQ4gPMdLBsbi4pLNzu2z/QfmrN6q28mXnreHP/Q+a5HZNhhYaWLCLp4+Z5cuX7YjR47p2q6tbWg+2ghr5cb6mn7OzxgsCCU8q6pjF86ft3vvudc2NtZtZ6dulUpZGXF0DyycP6/bRiA39iVnz563fXMHpCbd2N5RlwJ2SoD6EK8QFfumqnbs0H4b9pqWz7qPPHZL7J3OLlyzdK5im9t1G6TpzNhWQLrvA3p2+szrNlWbUrA51wyPd8Y2JBL3DuXqgfk51VZkYhw6eMAWr1ySSOTQgTlbXrymrt/b7rhdz8vzL5+08ekZO/naac018wePWK02bc89/ZwdPnxE+yJ1wg/7InyK+bK9+uopgaGs7cwl2bTi6m1uekokCuRLrpC39c1V2bViB8xzuHht0Y4evVnHu7S0rFw5iFg6KlD9QCUiuPFnz58GzTPq8Ioq55zEXWtrECbYD6JyxYWgZ/nM0Ibduj1w1wmbn6ra7NSkXTp7xnqtjjV7PQXR7jt4wMq1mm2srGj9kYUKHcqZtP3cl/xe/qi/9oZnQ1hozd83qfBmzV2drm3+t79mjX/1FQHpE3/nL4z+be/v87vbv/wvBPIn7aXofhhu1a35uW/KFmrv141skOLv3IgYiIHaWrtWN23Y6lhqvGLpsbJeFrsN3qyjIp7bYHnDUsX8KI8j5lu80bX+QYiKN7pemYP7Rtd27S/+w+sIotjpwi8k80OS5AbnfO3df+5HPRxG7/e2lUctPUhL4FYulq2+3XYL4mHa5uen7cDsjO2fmbBClk7rvk3UpoQZQOAuLq7aylrdmm1Eoh1bXtsyAoKBXSGjqZ0klMzlbGJ8fOSEwNrHMwZQDZkP/nL8xHErgRFtrEngCqok8SjrQVS/K+dCSjntcxHmYTt75do1m9k341ZSZDIFa2HvNA+WtfyMHDUIZnCnYGEs6/HtHc25rGceNO322IgCEd7m8r4GOrkQ7Xd9cuDftdcO9ZITHUXvGlV+UVnXwTsw09pr+rzic4lqn2CTCmaEjZ7q61RGaxjXzzEiX7dZ+8BqxscnVHeCl0WBm++pfT1VF3eo4fWcU3uJ0CmE9dWFAIhfBYLjTIEdX6ctInmiXLViriCLp3VcCFptYR8cD3tzPpeAczKQsqWCSBjspaPLCPVass6PAg6JSOkSDM4KFAccF1/xHGONMdrXJcQLz/7uxGjsvvdPt7XmUBfKEpRMEzJYQ2g38zY1ugS+kGbquPf9/XajrvGm7m8ElwjccHsZEtLel4CMdWXf7D5bWl7SGoDoc2enqc44aoRioWQbO5vWaDfVlZJH/MlramN2aG7a0tax8UrBlq9ds3YTLA7BRcVShYyVIeSyOdlJurV7XpZjYDLcC/Y51JWqYwdufYh4BBtLOgzBqKiDJTDOFK3VTds3n3jBLlxdsxbXVN0kfZubn3uLqPhDmz3feuN/a1fgYMptgHjoG9sN70pIp1UYQ1Ts37/PSqWclM9MsNiprCwtCfQY40HeRuGE0hbywm1+qAFRE+ITCgPbC1ZFeAaicGTjyiIj9QpWKrQ/0bInltbDeVOpvuEy0O+17NjRA8phWFq8ovYnhfkVyzY9XVOLbx3wkPZ3BXY3tRHAh4+JQdZSQalPQatNEgyzQq937UG4Aep8CO17/D0qdaM6NIIA2vAl7lgkB7xF2BW7/K4WjpBZIfvqsMmNm1AHK7UUayFgk8IxsLgBmo5PTGihYFEAIOVnkD9sXngdi4aAZ7oQuq56kjpBfofkE7iHILZcLCj1VlNFAAsFwC4LM5OzyJvQheEN0QHcNs8pYALl/Tw4k8BtVP6eA6LNt4B1Z7UhI7AV6vRYVDvKPmBM8JkeUtmzE/fGjgq3RIqAxY2ICt4/qvRjRgX3hdfFVkNda3W/7BIVU7VJm6xW7JnvPCUwLmZUwKSwicH6CQIthmlncl2bmICoICw1EhV9KSwjUREX4giaMOaTHRWZQdpy6aFtb1y1c6++JJ/amHNCrcLmUDYIxZKVq+Mj//QkIK1rgd1WACsZwxAVCl8n84OFFdXN+oadOfWaNs+QAhRI6XxGGSS7RIWPQUicgWVUTEqFwEZQP4eh78o7OZPznBS6nuioYDOnAlZYD4WQK2VZfMulqka/CsCBhxgnu9c9kJDQNQ/A3gWmfIxwjqhEsJLb2FhzP880c0zF5ueP2OyR2y2dpzPEF24KBnWkZOiWampMMRYoDgmMjMQLftKEaXtofVvZG5wrodp8xurSVf2JMpCupN3jgsxMqYMIxRxAI/8fPXrUbr/jdmu0CQQt22/91m/pOly7ds3DUnmmQ3Ghgiz4svsz7fcx+ZUcPyo2o7/TCKD0+cfvXyxqd2Wvcf7R/JEgQ+LP42uTDRaxSNZxBFwK2yb+B8QaERUhwDZekzjnacMYPi/OewLWgl+Rh+/mBMKrUMxyHwuahyjEPvbxj9vd73qPbfZ6trqyYd/4whfs1HPPWLu1pXl+EKyf4jMVr5EONxHmHK9jkiCI/x5V+NH6SVYnMbg3XL74u6N7EMLnKGrxA5e/KZ+3114mfHDyc/cu1hGAjMU3f3It6Mj58Z/4CXUBQgbwzF68cEEgFMWne8mT/eQEIJsVnnf3uQWk3g1Dj0T+6LMT4PVozMRcigDq8vxGsFQZTClyFPA0d696tWITLrixru9F1gSG0591Jy20kbou9NxDtPnlN+qoCMYavmmPFjThvUZAc4JIutH9RcWcJncnz7rKxqhhvYGT4X/vH/x9O3DsDuv3c3b1ypo9+e0n7IlvftVeffkpa9VXHUwO4CqbUjZ5bEaw9vkrn/4bdvTEfZbOTVhjY81+7Zf/kV1cOBXECz1tXCJR8Wf+zE8LnJuZ2edeyiVvcac7iLUZ6yfmTe4miqi4NjGPMM+4XYjnD5ARQKDq5z//eXvp5ZdG1xeFVezq0Vhi8x2fuT2dKm9GVESSVNQB5x9JxgT4rXuxh6iIz7oIcym7PBNLxEUYAzEIkW7J3WeVTZXfOd88O9onsiJQZGyypYoPwF9yHMXvI9EX6yKuIUA1CnSIijZg1Z78mFiTZDLFkNX13SU0fsx+SA4yxHHnm1fglZ5NT8/YrYSiz0zp/jz11NPWJb9DNZSTDepEUhi913O7RMVu11YkKsiJ2iUq+PAEURE6WCRkwZJoDFWnK+UJBVbrZDjOZGfRm3VUSIkZ1JVOgjgB4x6AvgQl72Ps7OUh8syi+OXkoy8SKM2dVIn3iPdgXmdc08HAM0iYNkSFzj10VMj6SYvG0K4sXBDQD3hA18GNiIrRuAcADqIe7j/1DM/syspKqDvcapZOiGRGhcKsledVsEqzJAEN3ZnPPPuciIrtnbrNTM/a4SMHrVYbt2994zG79767Ffz8wINvt4Vz5wQaP/3Us/ahRz4CJmbf+ta3lQ8GuIKV5Ec/8ogNITG7hLNmrdnsqBPi6NEjVqqWrDRWtNdeecHe+c4HrLG+oQtanZi0yxcu2rVrSwIrIBQ2N7flvQ5Jja0kikpEHqViQfU4IpOLWErNzurPW2+5RUCMREf5nK4H9Th1j0jXUkVzD3kZ+w8esma7Z1cWl0VSpLEHIUC1lLdCNm3lQtoeuPd2Sw2xTdKgtpW1TWt3zU6fu2KZPN3ELduob1qxXBAQCNHK+3MdGBOM2bm5/TomrhnP9Qx5VRsbduzoERF9tYlJm5+bVkd8uVSwzbVVdR4gGDl65LCA+hdfOWXjU9N26eo122nRkT1mt912h738wku+9g1N5CG13tmFBWvUUWTnpHSGvCCnrEcQb21CeRA854hT1C2cpqPimvae2GxcvXrVbr/9LtupO+kFX0w9LyvUVEYWp8w7PPNx/WZ8yc5UUSvezQMxRrhqrDE0p9AxTg9Rr2Vvu/u4HZget7namK0tLSkf5dTp05YrV2zmwEGtG3SKVcbGBdoSPNxPp+2//NqlH6Hp0/VzIAHa+bfd9t0TY8iiqP/z37+uu4BOicpPf9xSVc/hGK3JCZIi/mwvEZLswki+9gclKiAAxj71p0c5Dv5eXkjvWiIN37SjAlIlkjHxWPZ2WdzoovwgRIWe8Z/5pI39xT/x3ddrp2nbv/qvv6tzI3k/kt0ldK1M/9Nf1CHdKF/jhjfwh/zh29e/aZPVCasUyHapSZi6tgr4O2UTY2XbWF22dL+h/QEdQMeOH7ba9JRwnu0dgOmSXVlct/XNtu00exLAqQsLAQfdBaGudCGfP1uNZl3tsTwzCNsma1NygpBTAaJR1hlEXwhVw/PmXdx91VgY2OXTWbt0fsFm9u2zlbU1dclpWCg3wcUByknDjiiA94hEcJOgCz8S5OBS4AkA/2AGELFRvBoJ9HgMu12bu/kU3kns2QrRUpTzjDiGuki094gWp15Q81nUEBKLSMTh2FPMKvN607/AsWL+QuziiK+NIjBJQWQd684gWrnD/pN1AvwAwgRFv2oJuQbQ4doTME6YdLfdsm6zoVyhPlkMXDvyZcsl22w0rN0GV8JS2fEkPnN8ZsqypbxqXZwMZPEcXBKSIr0o7k3WMZwjmJsyK0MWRdwbxNrMBZrMuz52nvvc5Gikk1ERr6M7PXgXHAeG5TuYQ7/bFoHdJ7eC4aHjHlipUlagO9034GGswakB4wosgrXVySpEt0sryxpDErxO75NtIDWb7P9ajPu6sLU8Np+9th3aP23lLLQ/1yNjrUbbep2Ujoef9oddy0J+aXw6caIaVNZZTlCB9Ulcls2qHtB9H3i+CyJA2T4WCnb48GHhVxvbXfv6N5+xlc2GtQZp60loZza7f/YtouKHnBvfetm/w1fgpjyFN10IRRt0nUFuwxozAdnAKhUCkvC+Y8ODArNl5aJ7XmNfAYFQm6i5t13KFeBLKyseSjs/LyazMFbRIvbscy+oZQqwADso9mVsegY9Jmfsc9xqJp2hkByQOGb9PmG8BOxBhvQEtjDhdtrkFuBB6PZEqE+ZnMWSFwpaABSWG3wP6cIYWR0Qai1fv7zAGSb2CDSyQLjS2RcSFjUmTAdtdzemUg+GzSsKLzZm/I7bbXgQt3vMxqBpBy8pVpmg1EkSNqbuIei/xwTG5h7yhvdlUvWOClcnAvBubm3Z6uqaFul0NijO+7T99xSIyLE16k0p7UVY5PJqadxs1K3VdYYf9RrnJgsvvGzDsbrywAOmkBaiOObe8bmAtVogpMZ3/1tf1FOhO2PLw7RlP+Ae0IBikBcAcspYgKi472267nx+3EQL/ExYP43IAAE8rhYEnI4dFSqEwibDQTy3KIo+fWyYJser9syTT4WOikmrTU8rvFcExf79lskVFJTKeM7kBk5U1AHA6YbJa2GBTWdxvV657YpJqUAZp4AT+FhbRl7GzfqGnXn1BWtvb2rR5Njw9FXYsHw589qwTUxOOsEQ1BMxvFZKfbqXZLnhwV2uWjXr4q0NEbi9ba+8+JK8kPEBRm2XLxWlMhTIGMBFt+IBoExp881C32o4gaLOqE5Hi3S+iIq1aJVq1XJ42tOBAYkk/3zPnXDwMqtnnnMHFFEovZ5ZLCMclKGg4TNRi1AsRnBM9zQAXzyjbL6xlVN3Vh9LMScqSrUD1k8F25rhUCoHOo54LraCTRXHjGIvgsReLNENRldFW+RFq15Xt0Wn3RRIubXhlk/a6Ac/zVg4MNcBAtBJQccR4OZNN91kJ267TaohlHyPPfYNW7q2KDU1BI+K0UBA7gJ7XAdXGEfSKRIWI4JSZBmbYd+AqYALSmpIQg8MiqBf8BkPiu1oRxD3b5EUceDOO9Li/Y8gmEt6KIxUQutZd0jKiQr+lTEuCxIdUPRn3QX4YhHN74jgDcFvEBVOOG2qYGa8MaZ5psbHKvbn//P/zB547/utmc5LvfnPf/037DuPfdX6nYaKUXlFq3PEn6lYrUdgMgKSSeJERXMinDYCkSKzgq/+rmutL74RZIzgm6BK2sT5Cnkn3oE3uqmjVVtF5Z7sDwfn3AKC50N2huFz4nqB+uuTP/VTIs4ZdyvLywpvRXHjoKB3nu0SFd6hpiJfYLPfCxEFXO+QQeII5I0IBAfn1eUjYo/3YTjFdSvtXWeIAERE5mWPthMUvrrvCXIkEsgx2M+tnuJ7OVEh4FPAr4Pj8TXx/uwFieO982HmmwjGeyTX/DrGzAy/tiioUDhvKFSupd//j376p+2W2++3mX0HrbHTticff9ye/s637dWXn7WdrRWfk1mHsyiWPVerXt/RvPVn/8J/YXc9+B7LFqessbFtv/mrv2JnTj5nQ/OMo7hl5Ng/+cmfsjvvvEOANuA58zbHTYcMyl8AqcmJmvVIekm7h7vynlDjS7DR8E6DXle2BVsbG/aFL31Rob5cVw2/kM3lynL/34kKVlAnPHfJfOaV3fEcr6M2d8FWbnRtw3iOm8HrCAFABFld+XwRyX6tQYGgiDWRdyz6fMb10bOk1n0Hj6nJmPNYe/1+OmfBzwAGRNboHvtGLVlH6fxH5+zPE2uEMgdqU8o7c0cE70SNG/r4HuqoSNTX1wlImO+CmlHvEMUieiOe/b4dODhvt9563CanppSR9OyzL0iF7XMoaxm1jStFd8mROLeHcR+6jHS/JMbc7XLSMxMId06E92XtQcWJlae6nkKHoT8Hfg10L8P3TlToSrkyNMzx/DudHwMRFd4N5OtaeJ58mtAG2LOUIvHoYwhvb//yZzn0F/v9Q9wQQCOudewG9ZrZQz/37Zu2Yzcd884TrWVoNX1NEVFx8YL1Ot5RgfUTaz71w/UdFT6XMw7x+ebLlYcVgTBLi4iisOjyaRLQy8Fi982mNi7kiqptar2KQIVCoWTPPvu8lcpV29rcVkcDofV0gDz+7W/aQw+9y1ZXFu32O26zU1g/pdL23LMvyvqpP0jZY499U52CEKXNxrZ99KOPKBATwIA1U8GW6xvquMSKrjY9YS+98Iw99O6329bqqhTDpbEJO3vqdXvm2RfslltuscnatNYBF0/1bGJ8wp579gVrNTbtj/7kTwgIZH7BjgJw4triNXvgvvvt5MmTqjUefMeDtra+Zlmp4Yeyr8xnC9ofvP76GTt20y2202zbuYuXlKkFEE8NuVPftqnJMRsv5+yO48eM8GcEYJ6r17OrSxt26vUFq0zsM6D5ZrdlGzsbqvc1btirhPmJ+4b6mbFElwdf1IjYiDBHy5rPUlYpFezCwjk7NL9fmTY7W5uy48QSanZuv7386mnrDIb22unTdue996qrG7X1wtkF2Q8zhj/4yCN26cplO/X665ZJ521yctouX73s3esFgkxbNj+7TzYmLD+EaZNpQ8F98vXTNjU9o7kYcRWETjabt9Ovn7ZSpSoAjvq2x1637VaynVYn2NHS5U3XDA4B3j1ISDBEBd3tEpLhf07obyAqStmh3X/3cds3XrYDMzVbOH1a4O7y6po1+j07cutx2ZDxjFLD6qljbmy17BceX9Pc9of1BfBf/Mg7LFUq+gzSbBkh229kfwRoXnj3PZa7+xb9bu/M5Rt2SvBedAKkZyb1e/X/+/ev6x6I58PnZ286oL/u7biAGOGLMG+6OpJf/Fv2loM6bkK824+/eN37T/7Sz1iqVLD+yoZt/cPf1EuTREP7W8+LpImvv1G3x95r/kbH82bnkLxevF8M+77R/Yy/O9ja+a7rD+mRHq9+13n+qMfFiYU/sHy6YIVMwSbHJjSHdDsDm5+fF9k4PVG1xvaaCEaU45v1De2L1jca1mgBiues289aE4/8ZtfShaJ1sQ2ulN0aOtg/udgKsLag9V+ZR8OBLHQma5N28623CHPitRLzIVCVbdPQA+vT3r3Ao1HK5UVWLF9d9MDmQV+1QUc5nTlrK4fAn1VlRpDLgI0RwHLDs1LBDVjmEHwy9yHS9G6I0shmOwoS1S0VyAjHbHKqI/mCUJYtlTJrGgKZ2ZtizaT3K+M24BbWet5k/Y063vdmvqZqgRwtvXLuGPr5MudgWRdxGJGo3a6vDWSuBtzD3yNWO76/k3VW0bEvWSqGegOyxkUoaWFo/E82RZ15uVG3CnZ2dFpgmUWIOYJYOvMCdJUeen0nIqqQs/HpmhUrZcfThJeFbtzgiDEiLtQxuZvfGI9JjgDh2sRrpPfg3JL1aDptT/62iyL5euCPbug8mLNjLRRtu5T3gbPDoMNNEqi/tbYuwWIRYns4sIlaTfUcomg6HhBAIWjGsSEUrHZ18arXwsof6dvMvjm5lmAhyXrCurGxs21FRLqdpqX7HfvoB99lc9PjtrW+ZC11yGRta7NlFxYQRmI55rbJYDOMDXA0xi3YHbZavD9h3aEPWZZSCkXv9pVhBT5ZzqdtamrMHnjgPisUyra507YvfO0p22l2rZchVFusjI1NjL9FVPyoJ8233u/f/hU4EiyX1GXQxRPP1bBkDDS2tyyfdz/Ygwfm7Kabj1oFNX0P8sDb45iwKVphw/HzZ/NFIa6AoKHZxPSkrW5vaEPPRPzKKydtaWVNn9PvpazV7Kh4z2X5O975gM1dKScdTB1IQaM2MxYKfOoFojpTLAuablvsO5tpjv3mm2+2Y0eOalJbX1uVSk4Atjz9UgoFKhaqAteocpnAea3soVChhgUpqSZTEFQAEKLCFLZWwcGQEzEcOyi/5Tmn0NBo8+J+x/IlD6QGk1YECSBdOI7YVcACyYIDq1sqAECXBA7g7U/QFJvVeqthjeBfKxVisaSFlAWL7gpuANfJQQY8JRuaaFk0WfwAY+UJ2IsLWcY3KLRqNrClYtJ1FT2bYMghJnSRNmK9ITx8UWbDTNBfu0ObJSGMeFKzuR9aqw2T7R0VEBbfD1ERFz+pBMk66HW1QQDwjwRTbC/0++EZFQqTHABuTdj0xLg9+eSTOj66gyZq0/KmzWTyNjO3XxZiU9M1q5axfsrYxOS4bdcbyj5Jp2grNYUys+BHG7C4eZeKOSpHR2AiCxx+m107++qLtr22aFnri7Vvd/AZBvjwzTyEBYHlsQUVcFekDRtMgB8xg24rhLozo9CvtDWHrrCjawWve9T9PIO8ns07QHu8LhGcjSQLRSMv5jkXwBiAMVQEFHOQhh7eTSHn3RfKxOh7PoQUDBmC1icCedQRCeXWVVh/AKRQ2HmwIv7IEXCOVlOyEAGMoCUSz0i6bbo9azUJSR+zA/NHrTQ5Z+k8qi4ULx0bG+OcBurgEMDS6cg+zsPd3Wed57/daVirs6O5oosdVKujnIxOq2XNRt1WVy7b0tKiCme+4vPNeJXjSSYt79JabXLUUXH8+HEb6Hnp2cVLl+zZp54WyATZwedzP7U91xiEaHXAnecuYDdeBIWvOK7JzOlLhcqrPddHREFQXFjavxe4yM8TivaA2F33nvxFvy+iEbV8COEGrAof70qfNwALA0EZ3zSpdInFpDZioR06Xj/GbJXw0I0t9zxPpW2sUrKJasnmpmv285/6i/a2d7/HOukxO3dlyX7lV37FHn/sKzbs1L17DtBNxxUV+jGombkj1PI3sNKK1ya5go6AVYXH7/5LJDni8xDPx0lpL7K5/ny5KsPVnH0AACAASURBVLkXrqP7ysoCR1kP0dYmXmvfjLGJwF5ENjfr6yPiG8LrT/zJP2mb+DtvbdqVS5fstVdfFXDDxgvVMvYqcb8Rj2VkuaP4h9CdE4Bv78IJawr2F8pT2g0ijkW2iAqIxpBR4SQH88/AhqjildGctu3NrRAS62sRQbUCgcN406e5n5/UQUmiIv6bQOoEmevj0AHrJDFx42qHY/cxwH9sDnws+1qo7oKownLfKj2n2IXcftf9dvttd+oenXr1FXv1lZfttddO2c7muqXSLjBQCzft1umMhAusvx/7sY/bR37ypyxTmrbWRs9+6zd+w15+5huWSresj0JWmzwn9T7x8U/YbbedkLIKdXGxVHG1d7stooLnqTY5ZT3rWj/lSj3UiVgKsWEB0GT+SfXpYmxrc/v1r3/NvvIVB2a0kdU6QqdDsKMMIboieeLYD9cmzrVcg2R3Be8VM5uS1zn5HMfvRbLKXspFCXHuiPNhWqHKbvUThQQQ5k4s7YamQ85Ts0m0wDUT+B+6Tbmd/YEIddUYuo+7c0889xExqEdt9/ni38kmqlOzKJA6dKcGy07Nt3oW3MYknkOSqFC3UgQE9gw+AOZUemC3Hr/ZTpw4LmvIQT9jC+ev2ksvv6J6JY5dnutIVHC8WTpOBPwjlhClKEEBz+ogs6uMTD6XVLJ0TfCeXA/qK0AXBCHOjQaSIjB2EWTQPYNwkZIkkLpRAINYoNuyYa8dBDUoMV3ROfpSx58LHmTZRn0hG6+MNse7X8kr53ZjcY7n9932yUkK6jiuAUD9/PwB5XD4YXPuYtFUW1y6cEFjvkxHBURFnvwgBwDi+cV1SupaEHRIEdmoVrQ+LC0uO2mXdkCLQGvAcUD4fLkocUYhQydkwWq9om2sbwlMO3XqtPIbCGI+cOiQuhM4/se+/jW7//77bGnpmj30wYft8tkzVt9p2FNPPWPvf//Dqvme+M5TesYR25B19eEPvV91MJ89SafE5St2/tx5dVodO3rY2h0EEx2rTZQl7KE7lPV9cXHZLl0k2HlCHeAIHKiNmu22ze/fr2cDocdNNx3zuXh7S+cKqMb7jFfHBHDwnGNziXUp6wW2U6BI+/bNas3ZxL61Nm1XFpdsbWPbBqmM7I/a3Z6sJvrths1MVezEzYcsn+lbnjHKieaKdu4civ6inblw1XbqLavNTttOY0uq56tXrkhMA0BPXcl8x5rGekdWl6yeihA67BvyqqEmxqvWbTfVpcgcw3hrteo2MT5mhw8f0lqyur5tlbFJO3P2rGxcGId0rF2+dNlyaQQ6aXvkkQ/b+uaGvXzyVQWGA+60yFEkXw9bSTJsqhWbqGJXjFVUxgYpQrixqekKVGo2PM/v8OGjAt2uXlvygY2tIrYhCrxlXgIkxN6D8FXPqKDbJdpbQg6xH6b+hLRQVxGhv8265dIDm6wW7M7jR62aTdnM5JhdvXRJ9+3q0rKVJybs0E03C1zlkcKrnH0kGSI4Dfz1r1+98bL41k/f5ApcJ9cJgO3wOqJi9T/9O29dwRtcgYfqT1khk7dqsWobK5tmA4Rr9BZmrFbJ2+zMhM1Mjdn01IRNTU/a3K3H9IxcPXfeLly8YgsXr1k2X7WllS3bosMCZwy6L6ouRhUY3e+pVgLT8Holre76WOtQI2G9nAdLkj8/rxlI/R4z5MhwgXgEQG/VG1bK5m19Zc3xknTaquPj6gjUCpZm/+qECPtT5irmUJ5lb3z3OofaK67J4FFgBrh8MOeSP8DfAYXBWSAfIjnBfkDCUQiOQsGajZbmAH7Ougj+hbCXc1WW4wDRm9dQ7naBot67pL0+d4trr4E8KBnRnpM7vgYy31BXcY1Ea/Tpnoj25eQuUHv1NFdKLKLuEM/eiHhMDAQXxkW4uPaYhGADzfSt18aStGuDTtcKyoHDTrxp+UrFtltNWXv2Oj0PM+/2RZJjDTh7cL+uuYQ1QVjk2BoiXHLacOrw/SsWfTgduPjGMTC5EHDcoUwRdhDO0WvEXfeRp3/bs5L4evAnN73C0N4lJTKZccb1RahAvkPW6KQY2CMffNgK2ayspVnHVtZXRbhjbwh2yXlBBvS6zMUN7RFiDiP4nMLC2UcO6Ryd0JpCrbu+RVfkwIr5rA3aDavk0vZHPvI+a+ys2v59UyLCW4yP6pRq03Q2b88/+YSIdO4PxAO1DnUaNQxZs7jMYF+GFTlf7Sb1uWm9o/OTGq+Uzyigm65NxFLtftp+/0vfsjXyr4aYTqWUL1oZK79FVLw18/+HdwVuRU1PYdvBz46uBQfkXXGK1Q/WULSNZW16etJuOXrEJseqo00xExKKfVhoBzhRuBGm7Oxvs9OyeruuwlHdD32zq1eX7PLla1ImEUKJwgXwj+8FpFg3hAw5SCOGtueKNk20UvQ5g8yB0k0B0JxGvTYY2li5YtMTNZucADQgwJsJat0arbpNTk3Y3NwBu3JxxR5//Bl/XdZBPQKjmJzZnHNMeA8qHwCmeNhXyA0TLosYYCiESVSMagMYVIdi5lOoCbxdPgJibFJYvAXCADBRKOt8AKRz4Ro6QAAwz+fgl8ekHBdo+YrDsANMowpgESW4OoRRjdS0YfKXJVTR1QPu5RgAKW04XU0s1VBYeLVJUqu3LwZR1SvRHdeoywSfFxvNflS+iaEgERmRcjKG+4i6nfsEUcECIxuoIRkVux0VsZARSHaDjooIHHLOfBaTfZKoiCBktH4aBkAEYmJqRFR0NBacqOBa521mdr+yUCjGqpW8CAEyOUZERZqW1JTVmx6IGkEhgWYBNNlLVEQCCxDw0pnXbOnSWUsPe1ZUYYJCC2sVuhsgOWDZ3Ys7/i+lIBYL2aL8IDMEUOK5r0GOz9TQ2mkCooYiKs6ePmOLEBUhV0GBksEbNIJQSQuiCDxhYaDxFIAqbYbzqBQLQV1Aweh5FsgsICpcBQlIk7Ox6oQKQQV6yYoldFJIEgCx6ZZRqBHlbRlaUiEz+Z7nt1AdVzEAACDVSGdohULV5mYPW2l8ynp9Vy76+PAMFDbNWFvFceAh324rBhi4tbNhOzsb1qYjqdW2+va2usModJvNhq2uXR2p4uK9isUi1k98TuyoYENOm+VNN9+sYrzVbOk9Hv3a11UYoa50Wxdv4YxEBYWN2+hAVADq6RM0hkYEp9Qt+LV6hsBIGUvQ1x6iwhU5Ebx19CgJwscVyQmO0BkBmCaPdCxFXLvvRxGkzuHv8TV+DXZBy/j3CGzqfWXHtwtmObDmtiJjpZJt7dQ91I7gQECjsbLN75u2v/bzf8keeNd77Mp6x779zAv2e7/3+/b0E4/ZoLXtJNOoU8FDnx0IBxCnoE0qyXf91OO1TAKB/OxGREU8r5FtS+IcpHoSMOaZGkkVE99r06E1Br/b621k4jVhfAKozs3NCXzEqgbQg/NgDP3xP/4nrN5oi8AAuHv9tZPW2N4W8Sh7FVk/+Q2JREUEh+U1H9X0IrWiOgmzblfaJ4mKeH+ifZXyOpQpFSxrUviSy/zJr6+l9Iw0dtzyETI/WrPFLop4XLtEReI+BLLDbYZ2jyUeR5wr47WNYzWumf53SQBG1z85nrln4q+k2md8BMsyNr7tjuVyJdu/f17rNKDf6sqSra6uCmSCII+f7yRuToHvEO533nOH/Sc/87OWreyzxkbPPv8v/6U9+Y0vWird1LXxLhRIm4xU1jfffJMsTwDL6MaTtZm6Ld2mUUGCXNPsUIAhHRZTtRlRkCtsrkHJeuTmtDU2vvOd79gXv/glAV+aVwOTGDse4tiKRM911084sNt0uarOCVdee51dUBjPcUwnn28RrAmiYrRuRXKKYPBgfSk1YSCinahwd6D4nFIvxvHFNWC9iMQo68zO1rZvnEVAxU6ZMI+NOpg0wVw3Bjgf7htCDYDF6+drfx/VJwmiIo6d3T/9M7/7i3l5qPy1d73rHXbzzYDYbHhTtrS0bs8+95zU6/E+xA6ASFxIOR7Af2286aQMHZDdQLrtJYHUb6DfdUKJuYIxxHod33fvfKv77jDLiMjTPIzyEWUnRH23JeEQNVcE/0fPme6Vk45OVHjXI2uTaq2QfXWDC+RXLcwvsn0qImCKwZ1uv4M1IgAzAISPUe/oAqRnMsfmrtuhA7ukbgbq1SRRwWsiUdEb0l1L2wQqfTqAy6qPl64tebdapqcuProoNc/nc1YoY8VWlEIYYc7UoGTpVM6WV1bt3LkLynBYXVsXmXLbiVulrPzSF75oDz30blu4cN4eete77RrWYu2OPfnk0/bwwx8UcPWtbz2hmlnK3Fza3ve+hzSfEJQ9MTFuOxvbtr62bocPHLRCEZkBa2HXatOTsqdDsFAsVmSdhBCL7oZ6vWkEvfqziqd7QTljjCP83BFxkXlx7sw5CTPoqiBkm88BAKxN1tQpOlmbkNUT+xbANhSlFy9csv0HD9pOo2lnz1+w8dqURGMKoB4OrVLM2ng5Y8dvmrfaeNFS1F2ZnDUbXbt8bc3OXVw0yxVskGa/UtTYn56asdW1FdnNCgCUR3ZX4poYrk6eBzUwoMvc3D6rb63b/ffdLesKxDbNelMWR1jVYvkys29KIrFstmydvlvrokA9feaMFemYbXknOaTHux96j+ZHOl7WNtdtYnrKLl68bK02YqSUVNZYPxXowqFbmyB5RFSlokikfdMzyhshTwOiAjJkcWlFnbt6DjJYSXn3vPZhQ/YmA8uyv2p1ZO3BXiKvruKUvL+x5kIZ7t3RZjO1CWvXt6yaz9igXbdCqqf98bUr5DTWbOHSJQWWj0HuTExqrPdZY9kTddqqfT79tSs3evze+tkPcQXeyLrph3ir/2BfcteVr9hYecz2kZ1Sm7Xmdsu2NsiSOaR9y8rymkR1nQ5ivaHdfscxm5qZsbW1LdtpNiSuQq+4udOyVhtZB39nPSjZzvaWxHISvbI2AeiibKeTVd17dL33RECwdrA2sR9knmV9IcuNTomYW0r2jSx8cC9AzLbjVpqQIpPT09bACk5iHoReLlAcqzhQrz1lBPIt5XiNMj/BJJyIiF0JqsNxd8DtwtzimvmO9UjdV75F83WUzwqWQwgnEfh5qHRWOBifzXqCAAExHYQ+n1kqe1aErLdl15TVHMnaLmvQIA6KNZxErWENJlNBed6hy8OzD4qjUOnYpUFdwXqgOrJHZgX75r6ye1jPY9Yo8+UQy2fylOhKMfIpy56bxz6Ke7G5JWs8xKmscGBXgPWsu9XJcc/pQLqU8UwQdYHz++B00bpWpEgfHyZZTZkhIAtCBWy91CkJucF1dlwP0grXDazfcRx4/nPTo2fx7T+x4u9DF7r2tt59CenA8SkbKpdWBtOD736n1cbJAO3JLYI9QbPdsgbk9U7DlheX7cLCJesN09Zod7W/J8+E/T/XMZIufDjkFBeQ+mVza1uY3bDbtuyga9Vc2j7x0ffblYWzNjMzpTXlxVdPWSZfsnShIotviPTUcCCrT407Zfx2dL3BLrACrJOTgg5LY4G1dmjlasnWVldEfExNFm2sXLb3PPSQxFJLa5v25ce+bfV2x3qpnHWGaWGCEB9vhWn/Bzt9///3xO4ZGxNBweYFm5vlpWVN6ChHKBQhBvB95+GiSE/3BzY7U7MTt53QwsYkxSThvu0pwwefTb5a7WyoXISt+rb7OA9TasXGi34Z79kBatSKOgzk1ycwGg96Nl7J9nVfHNiXu9rUQ7hZ/ERa5DyQj8oPMDSH13cAl7KZoR08PKcgvemZSavNTKoNmABO2rKlAB4nRLiqxWOn7kG7q6vrrg4YwtYXER6I3aZY57whBwRw0Y7eaOhPVOhRGUcXikiVTEYb7pFCFTuBEMAo4CVYtvhCvgtmAsayRY2bQ66nK32D6pBJGn94ulGUFdHXZicSGfwpS6lwbeNGv0PAEqG3eW8RFHjA5gmvY0CB0IKn9sHQrukgnyt3I+MNy8wCzbnLwENZFWzEUgrPBmRD0dhhE62AR7cm8I4Kz6gYBSQHIuZ7ERV7rZ8isOPH50XQGxEVbAYnpqa1KEJQzMzOyfqpNjVpY1UnKiYnxwW4rm/syPoJoqLVabrSOOSJvBlRIVyArhhL2fq1i3bx9Ekb9FpWKdD9A0HFpicrX89oDxE9zRn/+hyIlFRWG/BcsaCFp1zw1kw8IXs5t35gYcVfmeeO+wnRRMYCG0kBfAmFc5zdon0D7yPyLNhQQPKkc9jF5NXazzMRiQo8ybmvbikEYYlPdVnPtzxAsWYTYOYb8EhUME4adQLG2Oyz6fNnlaKTMVtAecBin41+9zzXqPIgOgmR8m4pFIHRhgLLqYps5HxuoZjgGQG8WFlds6tXL9vlSwsqmJ2scEsM2RURONanq2WXNNgFVAeWk5Kcgq0igBmFPIrRo8eOWaGCpQSFRNq+9IUviCSi2MTOh41zsqNi5GUOKKyOIrdc8mfbAWOOG7VGKkuxB+HqyhTaUF3VjIKWThEHNrh20bIoyEmuW7BEOgXltbp1RxkSbsWQoBdG2Q1xrhm9UULN7qCTA70RVI6dRBG8iz9nfqqWiiL4mMd5TvLY0RVy6qj4mT/3H9uBozfb068uWHlyn0DAL/7e71h7Z01FtDpAJK1hDvKC3S3ExP+MziuqvePxcr4/CFHBcamYTpwT80+0mIvvG7uR+Dvfx01PvI7Xg+x+fLxvzDNyGzMHDRlHn/zkJ63R7El9emHhvJ0/c8Za9R3dFxE1gLsJMXPshFA3QQi9lhI6EcorJXso9OM5JYkYEftB1SXiOuOEhTq6UtARnoHCFx165LhEv13GqsZSIGN3Bxo/C+Hcgezh2XNLKhcU8FlxoxXnsuS5xfdK3jf3049dNbugssjPYFWjsRcAJWgXng/Wnfq2d0apM1E2RgDw4f1CBgznEolgNrnMR/vmZuzn/tYvWGXqkG2vte0rn/2cPfblz5qlGrLF0jwG4VYu2/ve936bnp6y+QMHtQlEBeXAr9shRREC94q5cmZm1mb3zQmopF2ccF8U5cN+23Nzmk175ZWX7Utf+nIICh5KCazW/QA26/4F+4Hoiaz1O9H278Dzbr2gsZTorNEJBPIxvld8hvcSFXHsRGsgyPw4rpP2T1H5FomKTIr6IuymRaC6Zd2IqOg4oev2mbukW5LIis8TL1UNF+Ye/pTNA6RKIjQ++fy/OVEhjd4bEhVoSAF9f+zHfswOHDjo6sHeUIr8F1982V4/8/qIuByR/qNgae8ydXs/wP+Q5wHoohyuYNGUsDHwjgq3C+V6MH55X0jO2K2ZnJu8w8bHoT+xgA/ePQgBRH2GKh5bVoCAaBt2HZmsgmSXqIiZMqzzelZ3G7GuW0/8M3cDPd1qyckN7iPBxZVqWZ3L1IHU8dExj0lbXtmRqGg31ekLUaENfyrr2URBcTkiKsi6QumPl7aIipLmvGtXFn3spPuq6bFwVM2ExWvsqEi7BdRYBy/yvOrgV0++ru5QrNcOHTpsR48e0nE/+uij9o4HH1SI9jvf8U67cOGCZsIXn3/Z3v+BD4hs//qjj4mYXFlZleXte9/7bkul++o+q01O2sbahjIXJsbGJHIBREqn+zY9NyM7DerLQmXMFi9dFQBRr7esUCqpVsDSived3jetPA3qilIRW56UuqYvLFyw2dl9soIix4J6CSADwIh9GAC48qByHn5OvUcHEDkreLWj4hfAJGvbgqWw5xt2rJjv2+23HLbpCcRi5JwRcNu31c2GnUMlXazYteUVq46Ny1p238ysBEgQhXR9sCdkTzI7s8+2sb4olGTLpg6H4UAdBtVK0W6//VaN06l983bp3IKdOb1g5xcWPF8Ny5RiUSQJQxviFls9xixdG4hNotKYe8G/nzp10q4tXZPVyNLKusJFi/mSFdVRUbYS3vjNHXXyG6AgVqYNt/KF7KIjq4BAbmAiKhCjMf4Z+9S0CNEAFLtD6vOh5Xiu2VeyQgK6odru9+3IMbzBM3b05mPq0oB84bPXl6/ZkflZmxkvW6rT1N6YMcBe8eq1RRuv1WxsYsKGAGnci1zaA371mUP7a28RFd819/ywP3iLqPjeV+6+pa9bxrLq6K2WqjboEAyfsenxSblmsAfOF7Pa17UbLSsV09oTX766JIsaYq2L5aptbjdtbRtFe1EdXDxTYCIO6g9k3+SW2hlrtL3rnvWN+YQ58PCRIwLpIZg9H85zC/iePYXAYmQICAJSadtYXdMemLmPOWpiuqbuRXAZ5mxIDXVm9IZaI1D/C3MJdk/LK8s2Mz2juZSuA4gRqdrBIfoA3Z4BBBEp6++wL/Ha2wVgkCES5mKDXfAAbYBtzov5S53Zwc3CRXZYuUJS19VRiM0rBDPrW7PuYlDey+chOgq9pqDm0TFgJRkEYszBo+xRrOo6HQlkuG76vlDUtVetF+yl2Eki5JNwIIpaqC27bQHnWL6aRH5tvYYQcaQUY5M1W9vcdKJbSjLEsV6/5Yp5BW5jMcQXDhpYLimkm32+jtuxPI6dTgA6PiHHs5mCQtm5Ju1eR9daxDGkTTqn+R57eRv2rNdrCmt46nc9nJ6v+z+8YGlwpX7XHrjvPpHRdENyfKwLciWQIBTL+rKVK5A5dR9nWMh1uXfgJFVbXV63Z555ztp9U5eEYya+l6C2iAJp7in3A6GrcjF3dlw40WtZrt+18ULOPvbIu+3iudM2f/CANTtde+6lU5YpV63e6isvCteTEsQOVoMtssmqsg5EwFGtlrUnBzeCSJEgdoC7C9bvCDO2RLJXihl1D95z973K4Frf3rEvP/pNZYk0ugPrDsAxuS9jbxEV33safOs3/n27AjfZUAsQHRUUtq709f0dEx8bgBIBbtubHoJDv0OnbQdo3cszETQVTI1akQmb93HgzMFjilMVZu2eWFh5r5FJocBdNjAoabyVzhWsPWv3Wok2OECBENoYNrKo8zg2ujz43idF1C955TLAtJJpkVN2Qksbibm5KZvbP22VclFtzbQrQpqMT4xbbXpGaklapdOFkr303PP22mtn1P3BRgJ1EikBTCZaWLXAuY+pMtVCeLUvFO51L2V0Cqa+L6aT8yQPgOsiUFqtx25jxRdh4GwP1bZIYE8IfTp46KCuLWFB/BzVEccgnV0QSNN2SKEuUiPYS/G70ctXxArth+RSKAzbz4FFW2GEIZCb44j2EQCxEDgsrmrvE3jSE8hM5wSgMYMESxNURw6y4DnfU+gdBT4gFN60WqCz3p3Bz266864RqDUCRwKwzkYlhpFHwD12VUQlfTIvJIIvaqEMeQl8CkHvdFQ89dRTDhpOTtj45JQNZPVSsKl9s7J+wiKqWmVc5gRcbGxtq30e0JwNOOfC6yOYENUDCnUKgVlOAnlGgIAX1Ng763b+1Es26LYtJ69sCgYnKtioUURJqSjf5jAmgsVJapBWR0WxUtIGF+sv2jPVUZHybggIs8sXLtnChQUVLN5V4WHQyesTryHH6PZSOVlT6T5HFW5qqI0vzyNEBUUThadUonQRBcUzAB4b1OgzLSumdCTYYrCqWz9JLdxzxXCEsgQs6dksWA6yo+fBuMw1LL7LS+v2/HOvSIUnFYeeI7+mABgUuAqYD+MUkOTw4SO2trZiCwsXbHnpmrWaIRdDNyeppmVC21XYRmB/RAyEUHCeP9mGTU/L1/rgoUNSxDEPcDzf+PqjIigAixiPGxvbmvP8fUKRq2BkLzSZ+xxwDzZPo0DWjGVyRc8dEODkHS4ONEEOAXhTsLpymOdXKhI+R/Ka3a+Rkp5nNL6H7J8cwI1Flzdv7KJT8dmJoP91APIeouJGn8fPKKyK2axUKtxM7wpKWzGbsqmxqn344Yds/+Fjdu+7PmTl2qx95t98xv71v/hnVt9YVgHogdq71k/+OZyfWz9FoFRjKHY1BK/2eEwR7IzdWdqgqL0YwCyorxOgdwSC4xjgfXiPSBbGOTCSfbKuYW1IkCNJwiICvbxPVDXzJ4reP/Wn/pRtbTeNjdLrp07axYXzarlOyfIKl/zrAdxIqGgDNfC1VPc8hPJGazHPA9glcq5TxYfjjKQYz6zfY65JKtgbcYnSOi8AuKjqFlERx+iePAHI2+jzH8dKsiMukkkRcE1elyQBdD0J5tZPsWMvvq/ey72lvCkpzB2s7e6Rvm07W1uuxJeXv2dLOO2JBc8uqaLsqAIAZlNrRL6QtU//7V+02SO32//L3psAWX6d133f29fufr0v07PPAAOAWAiAWEhC1ELStCVZRdmWKcuWY0dy7HJZZSmWXF4Sx0okV9Elq8rlJVZSlk0lppNoMRVLImXGkERxA0ViGwADzGC27ul979dv7fc69Tvfva/fNAYSmRRpm5ougjPTy+v/u//7v/e753znnNr2vn3u05+23/y1X7SuVQW2CyBGIZJO27vf/bRIy+GRUY3LxuamDpeTExMim5i7PJtYBNKJePzYCbvvvndoLb365jXrHCTs2My0Dmx0dXFouXVr3j75yU+KZNbjmAoBr6EJIc4h30vCLA+kRHxmnTj3Bo04j4+SaP3j3LOVinOUg29/xlO45+r47inEAiET7BtUG4qQCPWd1jSn8HQtsijq9IgK1GzMLTUU9Ev6+1RNej0sjUQwBWs58z2Ca6FeYdWO8zvO0976fQdFhX+NqXFo/cT+LF9q2QXS8NG2k6dP2B/9o99lE+NTIinohMTWgQ7v5194Xuu79tqeTYPn+Dgv74Qz+6ly16J9QdKVUrGJokc+YPcpRbCTzoDpzEX2ZPac/o9IjDj5FP6DmOwjKrSvKqSd8He35IzrT2+tZBxYA2nwSbqNgds/OWnby0jqe87j+Eaion89OlxfqSFz9uCDD6rBySV+4b+QpSPrp7m5nqICcAKQABBdQanB8i9mVjFmqiUUtEkQc0n17ML8gpP0GRnPyQIJdRshrGRUyPopXVQNNJUesr2qKxcuXbqsQGU66qemZuzChfOyrnDPfAAAIABJREFUMv385z5r73nPe2xjfd0efPxdNnf5sixgX33tdfvgB/+Ins9f/uVPaO/XTpQ8sKeeepc6PLFmGh0esfmbWPi9bh/8wHdYwvZtv1m3fCFjA0Ml1T28z0wqZ/PzC1bdI6STxgTApbZAKzqKWYsgxMj4UF1fr6n5680rV0WMMgeo88keY/9BncIzAYnB3N7c2lItzmuhAkGpsLFJOPa+zitYUOzs7FqB+j51YPlM104cG5FNEeem/GDF1hZWbW1rz77wpRds9uQZq7e9IQXQjQ5rbunWNvkSXgMDPrIHzh4/bmura1qD1aGcICC8Zvfcc9aeePxx7SsrKxu2ubFjly9ft42tbSuWy+oeBajjjOC5F1hFDdmFe+/V87ZX3Q2KUrPv+Z7v0XP3wgvPixgBbNvcqVqpPGjVal35hSdmZ6xMp/I+4d5NnbNomFhaXbF8saSfp+ns9OlzArLICIk7BOHaqG8031F7JyBTye9I2tTEpO0rkNaDTfkO8tZuzN2w4yeOi6DBEpSxLeVShp4um+xYtruvIPG1lWXVqVhbTc7MKPOHzBJ+dwLbuHTStna31X38tz63Fp7cOym/blsW7v7jDxgBgrv5INPiq8mk+HoPaDSourNRla+Y3+i7/q6tz7vbBPkUqZwtL6xYp8VZIatA+b36vmUzCRsbL9r05Lg9/NCDVqpUbH113Ta2d2xtc9t29xq2tr5jKxtblskVRYrihuF5BDgoNLWnRWeGrd0dP4uFXAUaeE6fOe17dKfjBEdoJIrna4hIXDZ0Rm20bWZqyo7PHrdP/vqvK2tgdGLMGp19a2AJrabRjM5PSdSNNGLmc1q7wE1Q6FFr9dZ07X3gT54tAV6jOjtNjUZmHE2nWZGJVJ+cI3SvWJPzBf0M+wSgNuuHcJxMxnNe5aaRtD3WRdXtEJ0o0dySmcwMKqZ8BuC87dmOaiI60Bgoq0A1v7cSRSyN/RTLPcgR1leAd64jZmGwH7N206nPGZ41PtYDnLG80dCdUhgnapH11VVZM+VQU+OG0e3Y9u6u5ctl29oGA0lJRYAdH2MRz1WlwQEbGhlWngV7MQgBqoGYv0D+K02ZbUgTaq19bNzJNUyJFHGXDkR82PzRxEhdBI5GtsaBtZs1NY9S+33x1471HtMf/KvYRh/IOvfk8eNSc8rGqd21ubl5KWHIsCwWaXBxPI2aHFKKObm4sGTtVkfnMopuCLhsHnUfe/uu7jn4Cc0FZHV646s3ndD0wD1iTqv5K9GxYqpr5cyBPfbgBXvxy1+2s+fOWKPVtS88/5olwDPRqqBU7IJN7StPCrwP3LDRqMkeEeUODQv5Yk7Wi7jWDA0MWSHrdpkoVmiWSNAw0GY8uyLcCT1f2dy2odFx2WTnIEb29mxrZ+suUfH1Xtjvvv43fgTO0eFB9xqerJ0Dq7GQ0IWID2c2axtra1r4eWghKNiMADpdpp0Q+C6/2OBL5x7aTnLIvzd4BHKgcQAU5prQW5cRsyCw6HPgpyDGboHOIS3QjvQ5Gw8A3wvh8U45it64McCmAizQiSXQnCyLdNIKLIa2b4MDBLzSoV3QosumCajngAj+fm3b3YN06Vqj4ZYgZBlwnUgbO/Lhdc/sQ9VC8BoEAFRQEt1mXK8flBVGF+w63B/QvQuj3zNFvitFuAasgNwLmG55xoHFbXBgUASDQIUQxqRNFA/G4EWvxTOd0gIXvQpZDHuBSiEUkUIe4oh7BjnFmNLFxVhzAFQQOXYhwWtRskwC47ALUNeqg34ssiz2bIbrmxs6QMLsC1ijA6nrYECtXpX8kH2YALzq7ra+du7Bh3p2Ff2d0lFlETffCBxG8oL36XJ8P2DEjdjBeCcq+H3MDQKmJ0ZHZLNBMaTcgcqIGH863obHxkVUDI8MqSsOIIu8io3NLdvY3JX87gD/zla9J/UUiBPGUh3PdEz22Vn03guAU2PPrr1+0dqNquXo/Oh6EJn8tlHBkAUSQm95LzGIXV7YAIrZtKFO4rlEFr/fpGgyayBwD1kpBDtfu3pVY8F9Qw4aO7L7X9sP3EkP7sarErkg4EsEDBJdERX5XMjJQNUhogJSBTzE7W+oNXm+eA74gKQEXHBgyMPjVdxkXGILURHDtF1z4d396iDkPcl+xDuYE5ZW+NQLL1wUCUPxE+3RDi1vvN6Nxb2A0KDMiTZwR8E6R9b8/wAb+o8Gh0Aq3aveXU8QLnYcExMTKmwJ8h4aG1MIG/fo+S9/WbYMEHnyh94mDKvmv0ZhwxEqpSPcQcgIsnnRGcJkFazugZUebi130vABiRlInuDJKvAy2qOE7pgISPVeM2QF6F4pwI1uFicq9IyEjIr+XeZOJEXvKvrUB0d/JgLomm8iu+lGcmUBdgyFTMpGBkv25/7099qHvvvDlh6YtOWtPfulX/ol+3f/18ettr1iTQizEM4dMyp6gJfAa88jiMHk/UB4//XEex7ng8Yl5P3E7+snpiIQrO6VANzGzqV+ZQTPSCRK6PbkEOPgv6/N/a/duzYOBYEAHB8ft+/7vj8tddDC4qK99PzzNj93w7qQTli5cZ+Sh4RDfL347EIQxnGO/q69Tm4ZzR4GE0fFjQDsaOGjPQxJulsVQVS4ooJ9ysk0wE/+gxj3jZvuntutdnqEDmvikdyJ+Azx+/m+CGZGtUo/2Rznq4p/PS/+/iLZ6dYAfQe1QFA6BCpNiZ4V3gsHiz15urMgONnhmVCib6zbp/7gmqIFIzVGMtm1H/ihv2yPv+cDtrPZst/+5Cfttz79q9aBqOgS6BiGIpGQDzxrAkorDoaLiwu69/wbkpR7zF6rw1C7aYODFXv44XfazMysVXf3bHurqkPT8FBJlomMB2P9qU99ym5cv9GzfopgfgSp4xw9On99//GaSOMZ/q9HNPU9GDH7oH+ORwAdj2L+HudNnNdOhB76KWueBLs+EX+6GYfh7L5qxfUFawO3JuIDpQ5EhcD6GIZ9h7wZEU1Bsafu7EC8c23UakqCCT7Lb3mejxAVh2tsJGVvV6pG8D+V6trDjzxk73//H7PBgYq1WtR92FnUbXl5yZ5/4UWBG/GQGesN6jXZpoVni32y93xBasRI8TC2up8Ky+6qizUGh7t1oq8v2OvEWife/0iSaOxoeJE9RQhAD9aNyhlAyUMTRBiYuI71yGtZMvi+7Kost9bz/cB3nB4JFJRR/E4RB+F5jmRFXAvJYwDoefjhh9R4hGIrrtsi3kXUm8D1/RZduQWdFzhTUFAAQERCMtpCohDDXkkEUCIlsAUCqJ+oYPwcGE/ogJ9VI0feMigqslmr7OcUho1nOCThxOSMra6u2vT0MTt3/rRVa7v20gsv2FNPPWVLi4v2jvsfECmFRdHK6ro99e6nbWtrx5577suyY6IOT6a69sSTj8uOAiB9fGzMqttVKdGoL7e3NqxSKZkdtG10fFh1Oc9nNluw9fUtWb9BHAjoUDB1R8BEZaQiYIW8ChqNGFvWpt3dqk1NTdr62rqdOHFcJAogFOsN18O4MyY0TUxOTAoQu3r1ut1z4V5b29iy9c0tWXBwDagF2CbKhbQNDuTs9OyoFQtpgfFkTAxVxmx+YdXmFlas3u7YHtYf5P5lMrIuAfzj9Zl3nO+4NrqSIU5oLuNsAri0trooe+AOtrZmdt99D1irBajTsflbK9ZooWbtWDqXs2YbgO/AygMldT6rbs27jQnzDtCQs9sHPvQhBb1evPiK5hH3cGF51TqJhJXKA8ocm52ZtAJWM+2mrP+keEun7ebCohWHaKRKKKPk1OnTOnMuLaM2ceszzqI03HAuQ2Xe7nLudWvB977n3Zbj7NNqKtyc8QcAq+5VRZpAWshytNmyd1y4x3LJrs1ODFuy3bDxsWG79uZlOz47azdvLXj398ioJWnIa+5babAspSTnKoC+u4qK/krum+/v/WRFr64Of3krUfH1py7uvfEpy2dyNjo0YmPYU3YTVq+27MTsSWUPbm9v2vbuhvIc6tWmjY2igktada9tuWLJkmp2TEgNXmt1ZHUjZz6yd7A8jYr1JNk0rmxC1aSzHIBttyMLHMhOrTUptzGqEuoMmcmZQJ31aTlkYPdHcPHG6rqA3eXVVRsfH7ORiXFrYcfNeiEFOWcd9kLUxKgauyKsAfdZZ7e3tkSegHsQHA6B4bUmLggoYz1PgzoDvIt1nHUQq56d3d1edkZUzGPzpDUWsqTdlA2hHCL0uY5nqCoDiuYGd5rgve4DxqseAIKKuXDBGYDaNME+mdN6KWxIqgNv4gCjYN3ysyzYE/t+yMUM2BBrKHttbARQ3U8Nwe+jwU2NPb4vLC0scDzVfsA6XioUZO9VGhy0ag1rOsY/LQKLM73GtLtvg5UhrWdYWKNcaNeryuph3da+TpA5jYjgZig1hIMhiiS4mrW+5rbPnN/TaTWHYLUH6ZHPpiyTwjFiR8q23/r3J3uLwt/+qSk1DlqzJQKatR21ImsxChYaAiBWyJXiveJqwu9hnrGPLS2tqPYplwZtZ6eqbCeC2MkKYlwhBiqVijcih0B07nNUKk+Mj9vq6orlwGZSXZsaHrCJoYKdO3nMvvg7v21nz52z3XrbvnzxDdvPFK1hadsXYeOB6OAv4JTMY7cQ62guM7/kXhIaelp7bivvtVzXSsWslQo5PQvY9C6u7lh5oGh7zbblBspWR03SYV8syRr7rvXTN98+8of+HT1zfNoT7juEHns4DQ+mWPFS2TbXN1QEskjpIRNDDdjqB2UWZDYkFjJ1adFjhC2TusEOrFiAGGgEe6eMinZf5D00yO1bHKwHxBbJEPyTneVw6boWXnnaeTA0QHjsOJbjABYQSJ1TTh4o8JAOv/2WZTgA7TdFWnTbIC0tS+V8k6CYRyYojzsOcsJb3WdXwccE1bS7trbJRjokRUMkGpytx3YJ2Rlh3g7UsAvxPSxOjC2dUbD+vgAS3Iq3NYyvM/fyHqTTM7DgkheGMCbJ/0L3GWOkzwe5H5sVpIN71TrbLgIpyBTVES9A3+WBjDnjw71xkPjAwxdZIOkEkCUUAD3+3L5QiisK8scYzoQMkUOnB6jXHUDlOhWiDbBAPgWbhbZpbc4CkjjMdNp28sJ9PaIiHqgZi/8vREUEJvhN/UQFPrfHZ6btC5//vObs8MiIDQ2P9KyfKqNjIiroXiuXveN2dGzU1tbXbW1jW0FIEBX1pgdwRQBOYLzUEwkVJD4+DhNEsIFCoF3dcqJCgUsQFH4wkn1KsP7pgaAt/NYzOozKSkWBf6gqMlL6cJDriKhIyPopBvsCAr2JlUy9rp8H8HCQ0/01I9AQgQjmCO9FUs8AngjgB5sSUYFawg+5PaJCHaJeVIiowAOTuklzhy6LQ6LCaQi66jOeBRG8swW2hNwb5kypWLIOVmLMCTIqJH01u/TaFbty+VogL5w48A6bGLzlFkFud+pKAwdyeZZ9DpPDcojgHUHt+ixv+Eo/UYFvJ7+He0BBSzGL9RMdi8wV99NM2ptvXBbAyHPH843PN+AG6yVEr7wtI+2g5cu7Y/oJOc0X7nPK10xl2zhGHD6wSSAMzp9R77rxdU0kVT9RoaZz1joHruP7B8TS7wRYi0CigmhvD17WNFCHcVRzhOELY3sn4kf3MyigZMMhoqIuL3n+zTpbzKVtbGjAfvjP/4B98I99t7VSA7a6U7eP/cLH7JOf+GXb2161FuT376OoOLTMOgTA+9eLo5u3QLhgeyYLtiA3j/e6nzDqFfRSoB12QMccF9bLSEYwjux5ABMKx5M0u8+vKao9+rI81IGaz9t7n/kWSyazsop44/XXbX1lWV1GkahQWEUAbyNIqX0Vq5VMIEYV7ixIMZA2vo7HdYiv9K9RDkIGC7C3ISqY676O+GGQbAffAxzMjA0Hcew0p5PsdW+dJ3Gd6QeR4/VEIuy2e9XrnHf/fWcG/HXjvYiksJZCdW25UTB7fSQqRK4otNt/nv0+qpKwI9A1q8svKaKCtYSQWor/x9/9Pvuzf+mv2+Zazf7dxz9uL33lM2ZprC6xxPN7G9ctX08CUaJoEAfvhwYGtUawBtNVB7nM83/q1Fn7ru/6bhsfn5JlC/vn3u6G/fpv/JrWxvvuu2DXrl2zN954Q28d3/IYGn47UaGrCL/e30skyiNR4ZfmXzv6rPYTFbKPi+C5cg58zr8dUdGvlInezKq9ZGUXm1Fc6cOIsIaJWItExYGJpKB2jCRptKp6yzPcIyp8XYlWXTxnXwtREdelmN1x1Popjo9+Rz5hz7zvffbe93ybpZJ0NxKc3FQH3ubmul167bK9ceWyZ3DJIi6MP4ScN0r29knADO4rdwqigunTv6bEeURGhfbbYCsXySjGo7/5Is6BeL2A+By4I1EBsahgbW3EENHoff3jsB4KhFLIeflqiArVh2GO9RMV8fPeyIKFBdaLXXv00Uf1vpMJ3/O8GHLLNuV0zc0pcBjSAdAAH/N+okLrRiBVeX/uTudERSFX0LNEF6Rqh7QTPXckKhKuCh5PlEUQrK6sKauBnIVbCwt24vhJmz1xTLXpxZdftnc+8ojWuwcfeMCuXHlTtfj8rUV79LHHbLe6J6WDnnGdT8yefOpxqTFre1VZH5ERsbG6Zg8+cL/tQFQMlqzTadjo+IjWF+o8rmNhYdGuXL1u42OTNjo+bjfnbkk9QXPQ2PiYzd9akC4OooIaaGp6yi6+fNHuveceqTbpykdNTT1C0wjrHmQ5lnI8n3TponJYWV218sCQra1vSl0BQIRymKU1Tz3fISckYefPHLPKYEHdtCgMkqmczc0v2/rWrtUBPajtQsMPyhGatNaxXMGfO5MVeDk8VNGKDclA7mB1Z1MNYKl0wvLYm7Tatrmxbd0uyR1Z26u1LFssKxi0QLZhm/NCSzYtsi9Tx7FbsOgMhV1KKmXf9ce/W8rDF198yRbmb9nU5DFb29qy1sGB1CIbW+t2fGbKBoo56wDwYRiaJr+sZfOLizYwPiqgDxCIjBLAVMgfznXYj8gDXt2yfm5pdrCnocGjY08+/rjAUc4tNCgArkFUAGR5JmDbdqq7shylLk8f7Nv952dtIJO06ekJW1latOHhId3vwcqwTc8et529huGeMlAZ1L6Omh1LnL/52dWQHXa0mrn772/GEXg7lcU36r2+a/OzlqdBKpGxZDdpnRbd8F0bGqxYoVi2gXLOpmfGLZtNqdueoF9A3RvXF21lfUNZM6jha422La3vCBgF52FXE65jCSmnWNudmE6IhHDA3PMYAINPnDwRiAqX1PMa5LaAOammCXmYrPmQh41a3fMYITbLJStXhmSziFqpdwaEfAw1LfiUFBEhv4L1lPWcZk2uS3tKcEEgA4hzn5PnB06UZMHEXF2rPIaYkxrqScgPaifV6bm0dZQ9gRrDG/aU6SDiAeID0oKQ7Y7s9HgPSjYiIBuChGYvWQx1PKA7h/IzhFGzDvFz+6gYCz5WqDI5g6DQFDbhWBN7sxMY3mxDda2G19AMyx5CEyC1Qy6TVpYO9ibsP5xJOItzDYlMWjgdw5FOpvUfJBRNAagzyigqRkestU+DSdva9R0r0vWvpokDS2Xztn+QsHqTXNesyAjGMUcYOY3I7ZYr6pRx2hTugMXhfqtup47P2MMPXrCXX/ySlfI5+5f/nCYI//hrf93zQ8DTOHdj5bS5tWM7O8wvMJy8lQYGdJbN5T2cHKUi84omo+3tXdWruXxRY6iG6f22XDOoORk3zmx+hndFruodspnKA2pgnJu7YSkwj3bDTk6N2vGJip2dnbLnPvd5u/8dD9j80rq9fHnOutmSNZJZqzZQg1Ibe9lM7SYcJuAazCtZjsm63DMCk2R+qZENlQ0knNlAqaTnsVnHmn5XCopdlI6yCPamWYi+ocpd66dv1Fp69/d8A0fg8dEhsY08nEx2WEkx1Km08ipY6GNQkIAzLZQsQO7PzAEhAvAs0kif1VHEg6/wOFcXcBiQoiLDYceD6lyCz0IbAUfvOBMAGcABQAO64CliY/e01AqppDZErikL+CsrvYR8/txPBlAce5u25RJmp2an7JEH7rPP/Nbv2LuefNhmTk6qe5KFW4HFoUMRgbn80tUKnVaOQWvf7LNfeNG+8sJF2SEhsRIJEABS95L3wFUWNxYiFj4sIVh8RBIoyNoXPR3UCURsQ/xAZqQkMaZ4j8w+1x/zKaKKgD/j4VWerAESVUBxCKXSvdNB0b3tuVa3rMrpntABxyaBgoLNm44ivsYH78e9Gutif+macpLI7bUo3j2/IO1dCAqLgniBlXamH1AbYJ3g8uHhQXUf0UWFJx+h2rX6np2498IhUaEeDAdj4nuIQKA6wkOYMJ/rt36KwG8EbgCq/T74kZnN9+TsTCAq2vKLJ2RQYGoup2DtTCZvY2OjNjDo6iHkpMz51bVNSRfZqBV6F8KiYnewA0PBrqOvIzFeL+DZzuqS3bj8qnXbDSvn2WyZ1ykFTdF9gjSV54B7B8jN/YrWYliYYe8jpRLWaxRWIsKS1uiG7kksR5otu/rmm7a9veV5DuWSZwQEZUzshIwduApV56CFaspRjR4JBvgNCcH9ZwTpZkTJQ93lHdhuNaIiAQlikLTKkzxYf3iBifomLaKiC2mlcHMnKiiQeA/FUslDlOle4XmVpUPbXvjKyzY3vxAsmijUfA6rI1VduYptdUBEYHm0Awo+ddJh9H3chiV753Wv4yeAbYeAn2diQKzSTUjYG7ZrPMfl4SEPAjWT3RYe81EpBdnAIfj69esK9XLVVwBW1TF/aD0UAR89wwJ08Jl3kE9kRQBkpQ7qkEnjPp9cI/fFbUtC2G94m6KGesG6QnU1PMhEWSMZaF2NAo/p7r3d+ikCnEdBzn7g860A6GFQMXONjpyd3aruB/8mTLuYz9p4ZdB+8CPfa9/6HR+0mhWkqPjYL/yC/e5//E1r17E+cKLCiVJfzfx/rjA7RN+cHJSyS2PmVV9PWRPc6DUWKtycpFEHUXhNydJlT+Ov5eofL/T5Oe9mCRkbGTqX3Aee8eLnOFz4nPOQ7bgWCxjsm3LRn55Pcfh55JF3WrXaUMj28tKitZsN2VbwhkUuSRnh1+Lcoa+j8koNwYT6Gich3WsHBbGP6FdU+MHLM1AE8gfbMwXv5Yv6GSl+khwqux5wH5Q8DDX2adrXpQaMQPThn27tw3p8SMxGO7M4jsxhxlyHcZQPrB8hb8H3FydeDuecHwxjrlOUu/uBETm496drbewjKzj4Qcqzt7nEyu9hzNeQRZfefwy5d9sfbxDAG7hjU7On7Mf+u//Rtjcb9kv/5uP2xitftkSStZ6u4LC+i+TzD70acyhOOgHVDqpxyOYb92Ub5ffovgv32x//ng/b2Oi4OvQ/8YlftqtX31SdgGWdOqgVxJ2z9oF3okWgvZ+siFOrR0QGQvFrJSrifXBlJvPP/ZZ9/3QCrEfcqhvNlZ/x2Y/Pk3sn+3rCc6o5pQYPJVXpXurx6h6oixH7Bp9Pbv3gj+7tJF+0fvL377WdGjgA/ml4Caqyo2SvSCjVa+EeaZuIqjU+FxSPoVLSFAmkTr6Ytve//zvs0UefNDtgbaW5oql8LTKObi0t2csvvWRrqOdEyAcCL5Bi/lrUXZ73xXjpNzIOIioOCVBXQMoj1K2jQn2q7w/3nYHpZfOImIzrIl2obe8MlPUTn8eHOgSQi6joVwr2jbH2n7AbacwPFRVuXXm7okIdpaEei00Y+lwgwdwaASVkS+HJ7JGRAPE7ENZbhY4mbHFhwWp73ulOEw61J7V8JHH0E2EuEKbNOYA5QvYJ38t6srK06vUX1k8Jt37iGvGRzhVzls2j6MhZDnXsftay6YKaTSAeUMqgZDt96qyNT45KgX3x5RftsUcfFYh1/NisvfzSy7o3ly5fkfUT+9hzX/yS24SheMkk7Ol3P2HJhIMek+Pjdvn1K7a6tCw7qRIqgWbVstmkTc5MCLyWlcdByhYWl5V1hwUVuV4A1+MTY6EmTwvA4+xxbOaYzjLkUkA+LC+v6FwDSAjZJ/V0IO3OnzsvNRmACp3Ju1WCatnXE+oQvXrtug2PjrtKvL1v+Qwe79hOZOz8mVkrFTKqkvLlQVtdWLH1zV27PrcgkuJdTz6pIGu6RqWMTWdFtly7ekP3gzMcKlNlc9UbNjo2Ztsb63pNSOKRUc+tY44uLq7Zbq1lzVbXMgTtor5Ns1501LnLOKnDlC7bUlHr+cjwsIAhzj1Pfev7rLm9bS+88KLdvH5T3d6QzxvVXdl+sdZMTY5ZpVy02vaWZVIpKxUGpKZZ396xwdFRZW3w79NnztjS8oqeScApzl2QZhAOUmvrPIu9JiHaaRsaKNvu9rYdP3bMxkZHQgYJNsL8LOqYkurMvb2qJbC17bas09ix07OTNj0+KgBwcmrS3rj8po1NTlm+ULbS0LDtW0qNAHv1qttfHZj9+GeW7hIVffXTf+l/vX1n69dvv/Wdff31E2/9nQ8tPWsjgxWbJEtrZMK2N6u2tVG1kQrA874tLy5Yu43tHHVj2h54x3kbn5iSFRBd9nuNlu3VW1JJbVX3tJ5Deu6HOpm1medJmQeZjBRjItpRA4aOcdwYsFAT/iMAPqdmUUor6mrhHrINwsciqeDv7n7XVpaWZHkHcD85O2MHKTJpXH3hNqZtK2QLatwjQJk1EOIUi1CAdl4fpwXICtQSrFVYK1Mz8HV3qmiolisW8t7Y0mhqnZLCAoXZ3p5bF9Np38GmumMkPNcaDTmEYAPMuqnspY7XFBQ1GWoqYWYtkTF8nfHhP3A3NUkEvEjYWKjnZbmt8xEkgjfv8XvYA1w15+B6bDiJKnD+DWaD8k4q0JAPyXhTqaWTSbs1f9PaNBnT1AWhQt1VKEhhwH3jKKIasO2kiZoXUikbmxy3NiHVmZxlEl2bGhmQ1fXe1rpqdmzVO4mMZQsDlinQ8Y/1U8bK4VypQPeJAAAgAElEQVTNuP0/zz5r6SxB4w2bnT5m+62mddstmxgdtHc+fJ+9+JUvKuvwV3/ldG8S/w8/OWKrq9g8zwubw1a11epYruAkk0jo/bYAe9WhuHyo3mLcweU8f7Pd9vMFNcDi8rJVa1Wd6cDgIP4hqljjwb8GUIy028qG2tokc65p2bRZe2/bTk6P2fHxYTszOynrp3P33Gtzyxt2fXHD6pa3hmVse69pyaxnhEQsC4xBGFdoWInnNYW56yEgjysltT3KQcpF9jdwGwidnV2sosrWpOk0NGoySMVS0QYGy3cVFf+lbyJ3r/+tI3AuZe7PhidwOgQEqus+gJghyFJAJScwgIgARqgjD/UFD5AkgV1tDCyu7jHs6gI2EQ+D9iAifLHdSqarn+NhxKaJrkKXgnuXNIWkg6z+2gIGZNiGbxuMeUMPdi6JvRPkglm93XSwjnyKVtOyqYQlO207c/yYPfTABfuPn/od+94/+QErDuUsxe/L0inr4bx+cKQjAPla2tbXd+z551+y+x58xF66dN3evD4XvH3pQPcuqGhpEAETfjUMPHJ3Fj86idiUXKHgh2hZRxTLLhUEkBIj3lS+BvYQMPwRuERqrK7LAPhyeKLDCjKEhS7aJHHgkQVFlhBoByMZc76X36nNTBuihzixMVPEi/AJsjS/NldbcP9gbjNZJz3wylVXpoIc/X4LNk57N2Adn95cTuw0hwjOn6Vywba2N3SfgMf4OUK1T913f28i9oMW/D12LKv4CN3REVChm86Do3K3dZDKjkzAi3cFyPfYDuzY1KS9+MILet9DlREPgGIOZXLyWMQ3uDIyYpXhiu4rORaEvG9sQFS4jQ+bfQzdikBbP0nSD370FBWEvW6v2fy1y9bkQEbXRQAjOaikcu5nSZA8oBsHQAcRHSRMZyEbIDKcQMHv3OWfHEi9IzN+AJADgnL9RWR/oTtTne6hUyMWRLE7AGBSYZbhRZR/EELf4zMWx99VNd7R7rZlKT84A3LpzfuLsIFyfdHKgUO9K6MiAOdh3LIGyrm0VSFSdGykMra1uWtf+tLzCpjlMCsLmkCS9Wzag20FNjixyI92SIcjcnhUuB0Q49l7a7iqxjudFtGG3DKfztrQQElBobPHjwl7yQ4W1QVEVwYdkV/64nOSqlIQlQYo8Lv2lS9/RV2G6r4NYG4vKyGCXH2kls+bGK4NQBSIiuA73+k6kRstdWLHrVuPeGia5kQg+LQuCoL1PI+ozrgN7w++WbonATiO4Cg/ewjyHQZVq9Oxz6rj6A6iZ5EOyyrZIF2RanTQUvSNVSr2A3/qO+3bP/ghW691bXFj137+5/+VvfClz1u7tuUgZNhDHJjzey6wW+3XPsEcEPUcC5GBIbS+X4ng4HJQlQTbEj2nIoXD6zKfApETnPVjH3Agzp0MZ63kIwZpO4HkRGpco7jeGJwtyiR0YznZ0JXPP+Toww8/og7YW/Pztr626ioZBctDXCd0wOOGufWVg/bcxWQCUj/fZ/PjSiLvTncw1C1dDu2f+tci/V37JfL1vG9P+gEUOZDgAFZOVrA27exsWbNZ05izV8XXiuB1JCMOVQqECDtQLVIhEBCyiwv7PfdRnfZhvvGakVjuB+YPr9tnV/TT1VgAxMpDzVcB5gHr0NbmprWl5rt9PYzj4d30cWwgmvAPJocAi4+Our7+xt/7SWt3kvZ//u8ft7krr1tSneL7Crc+Ss7Fa2Ttce4r5NCEKxPZFcgLEWFmCvFlTwQsxTYkfjCmzCUOQ+q2C3kKR5/F/o77fpK8v2u+//47wXNIBPQrKuLYi+hEtSrrA7cvE+AvojSoBdM8Z+wfebcnUFC6/3d7roHPAc898FwZmhYAAWhiwMs9XpOTcYerx23vNeTzxK/2vw+97+CJRx3oNoFcb5yjt7t837aGhb0yjlEkirmOTDZt73nve+yd73xcRB6HVw6z7PWs83j9vnbpNbt27aqyDTQXg7rHFTxOkshuQNaneVdwkQXBnKDrMex9ccwTWkedqHD7s75rV6aX2rv9nhD2G9TFgBuuNvZ56Xs398L3s56IMJCdPo4+T12xcJR4dGBCzTgaS1cdRRUNf+fAz0d/rUNNgv9zdW/Hzp8/K9DaeRu/QW596L+L1wLQRvUUa5FIPvkz7vsXCksur6tsHP7ze4uik1qC7nwpl7PaIVXTS/GLcjSfFdCfyRT05/g+hGxSWQTYIQ0Pjyq4+syZszZzDLuPhr1y8WWFaNP0MnvsmM3dnNP9fu3S6/be9z4j3+qXXnxZc5h7SP2L9RO1w9LiLTtx/LhdvXLdttbX7bFH32lbG6uWy0CsJW1sfERkBh2bhGbeurVkt24t2PETp1XzzM0vKmMC8B+Fx8VXXlOXKh3/rhr1bl7uMzZLx2Zm9AwxpgL16WYtD9jywqJNTqHWamrOUcfTDb2yuiZVBYoDwEOtxUbQbMJy2QM7MTthlYGi2982aapI2trqhrr9b87N2dPPvNcmTxy3xvqGsj0g76hRr1+7adeuXde9PnPmtL4WyUcAJgi4oYGinbvnjMh49vWXX35VGVzYG+VKJaknW/tNZemVciVrNdpqCuF+02BDg1C0QFPmXhmVyr7sPRhHAFFZXDDPAP2yaRsZHrQBrERqewLTCrmi3jcWvtlSSd2/mxubNjk5rXWfc6pUqcwj2ac5z815h05iqVvSaTt14oRtb24ouBdwsTJUVug9JBINOFwbyhXuWSFrVkgdWKdRtXyibSdnp+3W3E0bqlRse3fPCqUBm5g6ZisbWOrUbbAyaJWZcavv7Fij3baf+N2lw0Xx7t++qUbgayEtvlFv/P65/2DJA845GRvDkuyAdS5p58/dq9zRWm1HCr3tnQ09y5Qye3sdkRTgQ4XykCygFpfXpOPLFcmoAMfwrCLWZmWOggVED/56LSgFsqqZwSSwY5MbRLnUy6jAApyv0Tyqxk6e+WpN+YyAtMrKIS9gsGzFwQHVTU3lP2DTV7fkQcIywSqcYGLhEvWGteoNPctslNT2o+NuX+dNlvsiSfhQ0yiOHB1soJIiqlGJ8D7c+cKbEwXa73dk0SSVIyoMxkA2TQ6YU2/y2iixBXyjRmi1Rcayn0GW0GCI2iA2glKvQ4TwNc/A8EYf9tV2aDyKe3SsBcDIvGmW622rJlAWFHtswIxkLa4Dg5/7lBvR7tj62rIap9iyOb+LZCA7FmJGTbHcT8xIIF9oWiQbKiXsROe+TttGynl775PvtIHsge1tb1h1e9s2t7dtZWPX1rdrtltvSV1hSWo3HDjA58iybXgmSKsrYphKpLazYw8/cN6efNdD9ulP/d82OTZq//b/mO09Gj/+42CUWXv+pVdExrfaOA+Y1m4yiVjjqa/UVBbORuBc3HPuSY28KIWVQ6JBSrXs1uItt6GKeYt5CHnH0RwbcwwNjG5PTQH7VsynbGt1w86fHLNjoxWbnRy157/0e/bgIw/b5WvzdnN52zq5AUuXhm17ryH7cBrAZC3aaGgv554pWJ4slxpzNdi7UxfuO/6piBNDYZzRc8LcZq9fXFiUooI5Qa6Uz4mEztzFcvEuUfGNWkzv/p5v3AicUyfcQQ9s5jdTpPNgy05J0m4Ca9wHjlUNllYd9oWCHrqFxSVXTwSLFgFw8lzDtsQ3nChli4cUgbo9cMf94SKwCWAI2M0BktfYV9YFDLQH0xBQy4MZpVJZDofesG27tT2rohDB+gaworsv+6fRwQF74MI9NlQq2uh4ReFyHADrezuev4EcTeFGHu4DS7tTrdtLL12y4fFxe+XNBXVxwZgXSiVJxN22ysET1BAAPuq+Y+FPpa1YxpfaQ5PYGAE5HYQ5kGyazkqRPWLK1fOqzUUkR7ulDiv+LZBBhyb3TPQwQu+iAwjiHvA6bNbR4gJigetjARQbH5QcKBxY2LgehcQGtQDXxSLP67FqT05O2sTkhDUZI4KEycCgC2tlWeOEb6EAmZSTC6lsWh1GEBWST7bwp0zq37DQAOwKKj3o2MzZc70JfpSoiHkUR4kKl+p5eFQ88PZ3e0ZFRSQqAEyGyiV1ujMfsfApDgw4yZXNC2ROZrJioZnHfPC6kCHePeFFAjJxL2CCr3OfRQ6/Px7k49/5GUDI/eauzV19wzqNluUBXoM9Fp3Q2CyhqICsQs7pvpMOziqoFAY948HzgAMQFYfAjoNREZBZXFy0mzdv6mcL+extGRVuF+CEBSRFJBl4UATehO5Qni8KJgK6+omO+N5ipzYbPp9js9W8BTQJGoYMwFEgKvgahNh+2w/d/aBUL3RMNkSHIcqrqwRpv6yON/ygFfwVpK23AXAHboMTwaceEBbhmH7s57bOXdiDtyEqIFnpABJRkdG8OXvurB2bnRGAki7mbHxiQs8Bxc1nP/c5rWmjo2PWOUjJ33ruBn7z/lxGosKtmBzs8YIzAuYO7kYQWFZyIYibTkaen3a77kBVKIz7iaP4Wocd0d6dwwfA99sRFXHeSH2m8Y0A0yEIHJ/HeM+4RvdyvR0QFBQWCGnmVVXAxr6C3yFRASGGBwfsIx/+I/YnPvL91kgU7er8sv3Mz/yMvfril629t+UkBXMoWC9FUkbAabBu8snuXbg8Iw7UewZFvNZoTRfJjfhsvHXcISpcjSECJ9r5hENKPIREIrT/fUfLlkhGRnWL7qFym1APHZIXKLcoQgHD1lfWdCjhYObKACeb2MNaB8i0HfBXDoXAVcB5FD5O9kc1Ezf2qyEqYsYE4yI1DgotrRmoIhxwBQjEskWkSYJmhW3Z3sQsgH4API5jJMZioHc/URHHPJI5URUXu4XiwUF7Wbjf/evCIcHgVhzqQOcI2GUsfLuI84N1enNj3TpNX4f6P/qJCv+7A7Wso9QITgq3LZHO2J/9b/6yHTt+1n7hX/4rW75xTUQFIcskUt1xvkvpcwg/6P2HX+4qkkOrqfh8AILpeT1S0jEuEBXs55BnUXnWT07EsYqv1b8OHs79PoIurBXx+78aouIt9znk6lAHpZI5zRFZP70NURHVdLEpxWsIP3DTABPXr6NERZxLPjHd6iF+vOV99nJ+IE2dqHC1R0882/vZfqKi10RyRMXBe07nUnbPvffae9/7LerWjqGMgLOABFw7DQAXL74sKyjWYleDOJkY12sUXhB71KbK8VIOlds/xPXbSdiOJWW1FeZDH1EhFYOIilDE8u/YgRpqU4jrHlERmodEUihDpM+yKZDXPiCu1osfR+dM98BVklI9B8Va3JOcN3UFGR98nvoT8oAMufvuv6CQeXWW0hoeVJVxPkWigoyImL8VGyd6+xDgQNiDgFAQi6GKdlWN26htEhCtDDZq3YTs95S/lEYZm/Wsr4zXSVPdkh0c0HG4azeuz9no6Lisn06dPGPTxya1rqKSwbIKW47pY8dscf6WrW9syr/6iSeetO2dXXvp5YuqywCYWvsNe/rpJyxfQGG+YidmZ23+5i1ZP9134V5bmL+hXIJiMWMjIxUnKgoldQJfu3bTbszNK8wbRcXyyqoaubB9AqTh91ZGRxwQyzqIt7a6opBQAJbBgbIyKvDGvnTpkk1MTqorFDtexpn8LH720qXX7fTZs7axQdBtTY04KNcFonXbsmYqFtN2zz0nLZ2kmaxpqXTOWvW2gKOt7arG7Imnn5LXurXbsrfK5xnPhN2aJ5enKwUvNSVnE+YF9T7A/vjoqGUzSRsfH/ZzTNJsfv6Wn5GyObv/4YfkJz8/f8NWVlasudO2yuCw7YSQ3dHRUS0CqJdUm9BApmcKO9MhAW8QMZ9/7vcM+gwVDcTdselxK+Zytr25qfvPWsX7unZz3qZmjtnS8rLORpXKsMioCBSxB9Awx3Pn57KW9oP4zEyOj7nSPoNfOoQbzTOupARoLJKNEhTwBfrm9us2Mpi30XLOcmmz5aUFm5iYtFuLKyIqBoZGrJtMy5ILUKzeqltltGL7iaT9+LPzdxUVR/bGb9Z//qdQUBwdyye2Pm/lQsly6ZwNlSu2sVbVeaVVx8YI+7a8jY8N2uhoyQYGinb67BmrtbpSka2tb0klVa2hqmiLaCOrADUBRB7PGFvYXqNhw5WKztF6bvY9NFpNiJ19rW9nzp6RYpx6mFqRczhZFp516GR8FpcPcKUDztNNW19dE7ibLeRtZGJMtk/NLnmpNN0kLIFMXw22NBy59SsERalQ1NqNwormocqQZ3m6wwROE1nZD9EkqjqTDCY1BpB1CSlJTuW+8BuClkWYKDM11qlkCqJsAEc4DNKmRmDNqAwM+F5Sb9g995x3RV0mpfWJ12FfZf9UtkXI3IBI9UYjlAPgaN6syz7BWYLa0S2f3EKc2oC1Dns+3hdYCWd6GrJExoADKOu1q/2TivQmNS9NG9jwsbaDyZF3SVbFXl1rPnMWskah5mSKZNMiKrAGyyY6NphLKkx6MJewNE1FKBnSGau3D0RUXJtblEMFplwHiYy1OgcK0cZ5AwyG69UYUFe3m3Z8Ztzuv/eULcxdtUI2Zf/4nzg2w8ff/juDtrC8bgtLa5bAWqvdtVyhrJwU9hrqshQZqTRIejtbsCX3+wCmKUsu5qFUIo5PgVGiVkFlAm6mel1nFJ4JP8dVd9zCtFbbtXwmYfuNmp06NmHHJ8fs1OyM/cdP/6498eTDdn1+2a7eWrHddtL2kxlrkBOVNpElXBFYj9eFXltRwwiPSSY1vxhrmsjIjlE9qONLV3VPh8ZtsNQ2dlJkxDSVFaN26W5XRH+xXLhLVHyzbiB/mN/X/Tk6wRIC5Hq+dyw2dK2k3AID2R0yLw4Q6rQK/vw8/GKtQxCaqyR8NB3ASepBpOjj0wo7C4FyeLlKacAi2W5KkkfIzqmTJ210ZNhu3ryhjU9dtHQdKlgoLbmWQDl37xDgpM2Oh5jiFsupTleS6L29XQUXHSAHK2QtnUjYidkZGxuvWLuxa81GTZ2FLLpADgp3wv6lNGCjY5Mqem8tLKnIfPXKdVtZ37V8MW+71breF4d5gEXZNYWwJLwIIS3YJLGL4T3KM5BrDGRPPMyxAHIQ4Z0olCh4tgrcCaADBTGHkeihh0SccaegYKN3psS7R+nAioBmDIX1/BBCUB0k5V7R9Sz5c86Bee/g2vUNT9ZRZBSkbHBo0LK0DB0QjFnVHGjX6woa5F7wmoTC0X3IQZe8Ckk91akJYEpAep2UCjHRkBT7nbZNnT5z2+E5HobVqRA67fqJCoHiBGtKlUOnmL+fePD28fJuxUhUoNKhF5TQJTYniAqCqdmIyTIplsqWyeXVgR6JD14vjnvsqpasVd0STlTo+H+HLmbvSAx+3fy5X7M3L120TqOpECkFaCkbPuFBv+mUiAoIKwee3T5D3xOIikhW0NUWxygG0MZ/03GH3znXDaMu6XxQo0RggD9jkKvCHkNorcAhz/WyBAd/VELdrhdvWSc9/A37e6MQOqqoECgumzKlbutPZTe0W9ZqEpB4SFTE10ZNooAqYX5svF2bm7uljArNKUBfio4+kFzqi9DB7QDVIThz2/odOlLfuqZ/bUTFufNn7dixGQH/iVxG4AL3qVZv2osvXVQXR6k0YLW9ms3PzdvG+kbwylfDSBg31tVgGRPUQbxGnCf9RIVUIupsZswP5OXcCyIPqg/GPj4LERCO//5qFBVxTI6CsJH46H8OI0gVn8k7Abd8zkPcC7azueXrUjbXIyoqA2X7zg+81/6rH/oh208P2sXL1+yjH/2HduPKa9aubbt0OhRsvNZtoHMgKzQmdHUrisABNZktCTN2kiA+lxEM//2ICvVThnwTzb5AWEg9ETYv5n8c6zgObmnR0bMRid64LjDnPVvJCTp51fpqKvJrnzwixiqTltdoHlk6/qnNhm3VsMzy5x81nwhdiIwkSkTvlPJ77WG4Xw1Roe8Pa5XyZih8A5AIsci6DHnB6wv0TRw4UdGs9TII4pjG5yyujb7+ecD5UaIi7jGRMPLOdyxmXJWlEQnEwlECM66ph4c/F0b6eudkRFSVcRDb3tq0ffaWtyEqYuCx7xFYNLltoZPzLR2mnvnQd9oz7/sO+zcf+9/s2muvWgYLJhEVng3z1g9XHvTA8J6RnCssDtUmhwQghxKFlvdRFXptOgNRRuYL6hDuJyr6n9PDdf8QNPZ1IsgM+vajuHfFfVGtD0es3g4VFU4iHyUq9Gil2aOwU3Ay6+2JipAhFsKZUb8IxE8ktO9GQls2VUcUFZF00nsVJ3VIOB0d+2QmkpLUB16ffDWKCu9H84ygeG98O0tYcaBox0+esKeefNoqw6OylNvf55CLH3bDqjtVqQEuvf6a3bhxLShXVWxJHdpP0HhDSM7z09JkiB0S07EBRESFssPcvrNH4PiVaSHS+1Y4/IFsBFkHWHfo8BToHMLneQ9SFLDPqzkIq8BOL9PocN5+NUSFz6X+Wkr/Vi3jZAUfsZZgnqYzSTt2bFqKCrdnjK8RVYH+b/IVVtfcPta9n92itH+fkUUGv6enqPA8Kh/TrDrqqVHhWsn4ACRSrg62GRAV1DtZ9x2ftrIlDtICpC5fuWojI2NSVJw+dcbOnj+tRqjnnvuCPfrIOwUcHT9+0jY3Nuz69RsiKp56+mnbqVbti1/8PRsbH9frVIbLduHCPVDZyluZmZ62q29clXry/gv32uL8TRsaKskqZWS0IpAdS1Hm5+LispoYBgaHVEOR+RDtXscmyM9YtPLQoOeTHKD2alm1ilVWQXXFyVOnbHdnx7tysc8IGTHYLtFwNDUxpXuD+oKAaexZbt6ct8rImDr+aawoFJiPhHYO2dPPPGnNetU2lhctk8rZ7s6ejU/OqL7l905NT6sZC3uQa1evuUookbbt7ap+B8QUFq5rG6si8aanJ2XL9L73f8AK2aS1amTSkJ8Rle8p29rZsbGpSRscGbJOymyHLKQme05WSojyUMUSsuB1G2Blrxx0LItXvWzqgpI+l7NPfOLXrCmgx0nsU6dOyCOdecb+OTw2YZvbVdvY3JZSGqCNGgMVivzh9zu2Sdi4akw/R7F3M1a5PJ3dbZ2NZo7NqOmL+pU1ABsYB2L9zLq1vaWmHhTMIwMFGx8umbVrVkqj4h6zK2+8rnt34+YtG5ucscGhEavzu7d2RYIXBwpSlmB7+WO/dZeouMNGe/dTX6cRuO/mf5A9EvlaM1PHrLbbRERqF+65YHawb1ub61bf27Jabcua7ZQdm61YcaBi1Wrdmm12pIw1Wl3b3WtaFWyB+sUSli8WbG113fLZvOyBnABsqAmQPBflU8jqL6l1hGeMbQ9MhJqa56w8WFbDGJZPNHA06w3VzmSoAa5j4SQHiXTKRicnDH0V5zPWgwINnKgLcNcIdkk8p1jMAfLyPLPHQYqydpL9yF4OBkP2AGsujgsiXXMojcmPcHxlG0LVEra96TUNWIlyDKRYxGGgIScAcCfWGjAGnDTaLciNhpwyAJJpR8P2bqAyJGcS5W/p+j0vjCZYB7P3bXx8XH9XDRVAAbAfbLMgw6PtqtcCruTg7A8JgrWy9gtZYiVEQqgKDuelfTC0dMoWb827wjPcB9W22CrmIJ+afvagCRirZynfUS7kbWR8VA4o2YN9G8gn7L6zJ60MyZVGmZGUBWGuNCj7p6s3FmxhadVtuA5STlTksyKlaNbEuYX6p5TP2+7GmuVZQycrVsiZ9pR/9i+Gek/Cz/zsWbt85aa9+OoblisNWDKVtRYNrChuIJYJ5t7znFZwM/LhqBNQB+Pm4XUZ6ke3wGY8CEJH/SML1v22rSwvyTaccy111UhlSPebn+de12u7lsuk7KDdtNnpCRsZLNmJmWlla549d8puLizZpSvXLZEv28Sx43btxlxoDMNSn9o6pSYE3XPlsHiGHc8AN5wGZ0AD3TtqsOCygQ8XeyTPBA3j3OMmihldU91dXIoQ+neJiq/T0nn3Zf9TjsA9BLriHYqqIktINt5tDgh7yCvdp7EzUa2sYnRZ4F0x4YeT6JXq8QvO4rJ4Fgp5PURsMBS7laGKTU1N2drqqtX3airYKDpZCFiU8QQ9fXJWHbk3bt60ep3F3P3pOcA0Wt4NI29b/PPprgokAQs6xSbe71w7CwzdQ8iT8VDNkIXR9aDtkQobVNmw+t6rblsCEJ3AYgJrGhwYOtbuEN53oGC6TvrACuWs1eocIM3KQ8O2s1cLHWW+2MNMd7UAuod4tL6Q5VKQHbNq4TEImIVckMXSMx3q+jl18/J+0v4e2Bywh6C4hgigIyseTDncx6+xSc3MHNOGLCubfQ964nvZtBg8NnTGOfopo5rY3d3pea47GQBxw/1qaXwzOWSMOW3gB3QssGAiwUb6KNJmV91tzX0O00ioHdjfq+8FCSWqBHwfPb+CMO1+oqJ/7scDvFQe2JAJmD7suOZ9RHAw/lwEbTQmCvFyz3gOGS0C6zjkpjM2PDKqYooiAoJiYGhI+SNsTmwKEbCJIIDkgio4sODB7//Qq/mwU9vxt3gN8fPqmu7W7dobr1mzWjUsH/J0RkCkMGfVdcbmVBDhxPWxmQqEDIoKCiEUFXRpHCUq+oEsCpMrV664tJYOsGD5xGv1Wz8ViwRpe7cBO6aAktAxqd4DulKi9ZQUGE5URPCW988zz5/MQfmQqgvUgRa323IAxTtOulJUBCZN85F76f6eLnvEroFJxvP20kuv2q25RW3m0ac/AugRRPE/fR2In7sd8HFv9P7xOZxfTlRE4O4QzMNTnnH38MwCdmADZXW+TGMXwXilEjYyNq4uxUabud1U+CRFdSGTta8895ysfbT2BPBbII+34L6F2OoHf50Ac+snZ26876rTafaku3FOHp2DEayM9m+Mb7R+cmsjvze9HvBgYdQPfvY/f/3AZQTo+fpRMJjPCTQOFjgQWG26jap7ksxS+DFXUKa87+mH7a/96I9ZrZu3L1+8JEXFysIN69R3PXMjzsEAiMXfq55VcoQAACAASURBVHkX1CjKdgkkld5zUKrEa+89d30A4SEA62tIfE7pXhdwGcguRp6vi5CXXz/WcOFZ7Ls2qVfo8pLViOeFRNVA/6EBoKrVcJCDrizI8bHBQZsYG/PwU702BamTxvNrqwop3NsDOPaMFfVWE0ynYHrvLJXiymeXA319RWz/c9IPPLsS6g6KCv1+fHSxTGTe0x27K0sXiny9Ro/oiETJoR2Yxjv60Yc/+5UAR8HvkE3dAz7751bv72Eu9RNWvpb7IU7zMOSzcA8A8NrYywXFYT+47WRgnPX+FERlqOThBzRbpOzehx+17/3+P2v//lc+YRe/9FwgKnT87SOGfT3x9xTed1jz1f0bvxaetkMCgU5BrCsD4NvnAxHvF88JRLVyDXqErlaOnurkLWsZ87ZPTXSn2rF/PvSPC+Oo/yT9pyva57uIhPChwxG8gnJzQpdyzMCRGsfJ+NvGI6rBSD8J94PO6XjffAycNIjrbo/sCQQWCoL+9xqJMX1/UFR4d0q0qYr78e3WX7e9bvS/O9JcwHucmJ4QUXHh3vvUec/6C5AMUbHf9AwvDpT49b/wwguqk6iT/f0F1Vp4JmnacOuntDqzndjxMY1EspRBwfoprp89wL6fqAhrkZQDYb9mHeF3yvIpvLZbq3oTDB3ucdyP2qS58uOt9nA+yw7rnn6iQvf3SFZNtH1kTnOWPnnyhOr4aP3kpHHIL5HiJSVAFwCHj7jv9+/lIuqDokMZZwmakTwHp0dUbGypc59uX8KgqJuVSwdBkSPrK2+pNGeMnM0mh+ygmxKwhJqBTnrOHNPTx+zs2VOqB1948Xl7z7vfrbMHwDxNBnNz89aoN+0dDz1kG5tb9uyzv2Nnzp0V2VYo5+38+TNWLNKw07XJiQl75aVXbGdr2+45d0aWecVc2kZHB3V2aTS9E5Vg55WVdXvj8hVZwA0MVuz1y1d0/qHzkVp+bv6WFbF+aNSlHCAbi+cG4IyFZWJiQvOOv58+fcreeOOyZfMZ1ficrbBuob7dlOpiSg1WV968ahOT0zZ7/IQtLi3Jsmp+/rrlCyl75pknNcYKoG3t287mtoJyd7Z37P5HHtb7Yx9nj5knK+wgoWYall+UKSi8scIYqgyquWv2+Ky9cvEVe8cD77ChIRTKZjtrayJrOB90ugmdJ6hJpmenLVfMykc+sZ+0Rs1tOmheo5kJYEnKZUtYdQ/iwdXpdDpTm7EDvPTyqzY4VLGRkVFZldCyQOA1wOdLr15SKHgqV7DNraqIq7iPUdcRhnpz7mbP/o97AlnFfsDchtyg5mBu8UENMDY6ZtMz0/bSSy8JyORrI6OjBtAHsEowbm13y07PTNjsdMWGi2mbnhy1m9eu2syxWfvs537Pzpw7b8dPnrbF1Q0rlgdtcHjQ1jdXba9Rk3rlb3/+bpj2nfawu5/7+ozAIyu/DR8hQD9laSvkStastm1iYtRmJsdtZmrUBsvk7uzaQbJjuRIWRXt27cYtW1zctEabsGTyK2noSFlH2QWuHmTfyGXyAuDp+PesBc9KYF2XFZGZjY6M2PTMjHChra1NkQc07fDMyfaaPaAN7pG2XCZriWApjvoNdcPQcMXGpiasyRkyn3V1A/ljtZpIGAG+mbRUYtSJjWq1tzepmQp7n1ZTexK4VcQU+L25fNaGKwM2PDKkdaUyWHG8pzwQGmdxrnACEwWYW2snRfRi8YkiD5s6Gmbpjmddp7bhOgaKReFeOG1wdlT+Z7ejpjdvvvXaJp59qLWGR0Y8B+3AgrKjY5XKUMhaQGXJmcQtnwXGhzMyeUzUF8o/5Oexuut4Nh1nE3Cc5WVs+sj1IH+R1RTbq64lsWMHC6PeldpVHQs68xVKBRseH1VmU21rw3KJrs1MVGwwn7bJ0RERYLVmy/KlIetY2m7MLdjC4oqsnrF/apFTm0tLjeMW7hkFRHOfu809kb78V8gc2EApZ//wHx3Wpn/iT65aoVyxW8vrlikMKLOIzBTsE7l+9srKEKHTnpVHpoTbVntTLWNOTccZB9wE4J/mVbA59lHslTiXgc/xb85FOATQ9Oo4XNqa+nmT7ez506dFVm9trtmNa4t2/p6TImlQe+w1921iesau3ZyTIwy4mAi1Ek2nTtqRdwvpwLVAzkUFCHuwmlBQ6FK7oWZWbmha2AuNNLznvUbTypVBNXJjT4baEZwnkZ564k5tVl+fFeU/s1c99T99zC7/16ftCx99xp752Ttd3A/Yb77+I/Ztg3e+8Mbc5+ynf/hH7R+8ePTrM/b9P/Ej9mMfedwemR7wLzZ3benS5+yn/+Z/b//8yPf/6C9+2j46+axlnvmp32eE/o69vPhttvj33m8ftH9qq3//cav8geO5a8/y/T/3B37jN9U3PFiEmaTTEMbRg3PpaAG8lTcsXsXIVhvIhT04kA76UqEssJEFgAWNB5EPfEAVyp30QEQKPNhTACwWJV8AQlhgp2v5gneBryDTLeS0CZw7e0JF/+TklL3+BpLDTW0WAIVROsXvivYfFKsiB1J0HkGwuOWNg5YetokCno5WFna6RykyM5mkjQ0PyV/1oNPSQQbSAGBsp1rTYaMLEJNM2V6rYQm89HfI8yi6/IyDqaxaPIJQrgnBF9jBTyRZvsBLWgbolKZrPXT1hnwIwgMJARcABhhGt5hCkDpamOKBlM2/urcnIJB7Q8eRbGNCIG8EmdTFGjsUD0ybKkAyhyNJnhUo1NaGFzMDGE9keHQHAKCxMbFAdg7aCkFifCsDQ3b+zFmB3dxPFv6Lr17Uplxr1LRYMhYcZtUt3Wlbu9MSYcE9Qq6NhUG/9VN8mCIwEX3h+62WIsASraoiMBmBVe9+pmMKoNiX6HarYY29ai8EKxIVoISRqOC+RiBeZANdilgOpD2Pgd9Tb7ilSz+Y0w9CRBBAh+4AlEKcddt7dv3yJXWQ5bD5yHuIeT9RQVdzDC2lI1Nek5BpymfwnArICsAsb8L1brP4O/k3YwJRwYELjCkCm7HjUsVXLqfiLIIZ3rV20CMqGIOkgtIPuytjILfGHksnhXWXvTNGNmH++WDZ7pY26ghIiXDUtTXxhHShQbTR8cBul7Myzm4psG+f/ewXbHeHXAu3vuonEnyOHPpfHwXf9NVoyfIHKCoiINj/+iJoIKIODpRRMTxQtvP33mMzM1NOwCXMRsfGLZnJyW8zXx5QGCWKqt21Vfu1T/w7WUhIJcJY9ikqYmfqncCiCBLyDNO5KPBIqC52d009P7EROxJPR5U9/Ey0gFKnIB1JzJ8wXr1r6QPr4jPXT0BEwLh/bsWv9493/Nloh8b3CMSiUFT3J/Z0Wc2VSrlsTzxy3n7i7/xdqx8U7FO//bv2P//zf2E760t20Kz2gnL7f3f8uwDrXhd6BLQ8t4bis79Dvf8ZjCBtBMGEbUb1lUDPAMLTlZtEGu2+sw4o4rWL5Uh/QK/fTEAKvicSgXHc9fu06vgeIPu+VtNazT3ZYjz8wP324LmzXkCSBbG5aVubGyK2meire7u2sr5l87eWZcGhqLsEQLUTe6xHjO/hPuNB2dr7QtdzXDvv1BnNnuiKCrd+0kOagudACu7ZToxms1kX6ObWHai7HGDvX9fic+bPjhMnITGgZ8vUD0TH+d1PVPAad5p3/UVVbz7o/rv9Gc9/HBPuAXNtv0lGxe3WcofX3P+KAMc8Y+RaQdoT0p2w6VNn7M/8xb9kv/Grv2aXXviKZQ/oWsdT9+2JCs9sCIC7sxROgun6DtV2Atr2XfkIqKiJ1rdO8R55H1gLoKgQkN9HjPH32+yR+n5WhHaf4qMHePfZy93pmZWyU+vFPq2MLpUPXe69e8velQAQT1sqARjuzwP7krR3qncOiRvmzyF5gSrVnxM6rvtBaW9gObRKPKooUHhmeE9xH5LdmsKpewuqKzwiaSTy8qsjKuK8UK2USip/6Oy5c8ox4B5kswVrt1B8dqxBWGi9brX6ng6pl69cltWYFA6htg30leYlcwsrNYENaW806Ve8icQDmMCGNNRlkRgNO5vbYvJqqJZZPxpkMbj9gKtUQj5LyHhiLBUGHLJGONDyvg6bKML86bMjOyTRQsUa9py4fsZr0Z/MyZirFfKp+HnW/YHBoo2NjfQyKqIa8DCs2/Nbtne2lbHAWMScrLi29u+/HkhPcqdbIMQxdUWFExVy5mE8AMBR1QaiAkA6lcpLXTGTGFQ3IsHJ87eWXPFYq9mpE6ft7NmTsvB55eJFe+qJJwRYHJ+dVYYE1wgYd+7cOVl7PPd7X7bK8Ij2/nwha489/k5lBgGqTU1O2vU3ryts+cI9521jfcUySUJas7KXgkiBBOY2o5bmOvKFksD15ZU1kdWLi0s2PTMlL2/8yAHztY9m/HzEmYkQ7enpKY0bX9/Z2bbKsFvF0ghC3Yeyma/RvVvIl7zhJZOz1dV1NXzI6iKbslpj1yYnR+z8+ZO2s7WhGi2bK1gql7fq9q7dePOq/OnpyCSnJYvl7oE3bK2trGmtB3Sj9iOjpN7YU8PR8sqi1Azf+u3frp/tdlq2ubwU5jC1S0pECJ3C91y4x7KlvNWrO5bkVpODAliYzaojlOwH3hPkjJTRnCXJgQCs4VzFmr/r9eHQYEWEB6p89lV8yg/SWXv18pu2tl21ao2fS0vRzj4xMjyi57lEtoTsOxt2/wP3C/BhbikPsd3WfGUdp4GGhjg1l4UcHz7Hv109acoo47xVzCYsZ20r5xN2YmpUHbaX37hsp06dsuXVdUtlCzaBasWStrG1ree8MJC3wZFhZbj8rc+v3LV+6t+q7/796zoCj2181oZKQ7Jeg6xYX922xD6ZP3krZlAz1O34sTGtF8lswmbOnpZibWluyRYW12272rS9esdW1rYUqk0TJzY01CrURure57xbLut55vlhz3Sg1ttwILix0mUPo5FV3fVkbKrR0M95PK9YVEFON/dqNjgwaKvLyyIWxicnlHvT7LQE5HowccKGUGHtow6meTKtNRObvBzNAwmaFz2wOjbVOFCOA8C+iA3wFfW/JqgDPFuUszd7Fn9CMmO/F9WBXOfCrQXVOixYy6trtr6x4cSN/qPKTAjsTgWrZfZ12QChYghBz8KDwt7q+3iwmZZlaVYkrlQrhYLUFMPDI2q2kn0Q2ERoLopnMSm/yHzt0Aib0totRSbZsHIqYG2vyRaLdRwAnn0vCdOMAjubEdnAwivrLeFajimxzmO7xfvdWV8jwMIKmYRlDjo2VOZsn1WDbwI3loOEMp/A5Pw9eiMxrb5YX0HQ8F8qkbJcJm213W07NT1m505Pm+3XrZhL2v/yL0d6z8NHPrJpl6/dsvXdpnWlxEzqvAT95VaR6lx2NUk4J0ZrS9WSyt51WzD+BBdhXHnfEPCcXXFzASek5srnsnZr7pZUiey5rnSsWj6bUbYH7i/FfN6quzu2tERu1KQtL69aktzb/a6dPH3a5heWRNiIqGE2pJ0M8vFO6jUZA+ol5oiUOuCqhKEHCysRFh0aP2kw2hf+UhoYsO29PVcppSGyDkT4/SEnKh63j33un9r3Hzez13/Rzr//H9r1tyynTlRM//qT9uCP9n/xXvujP/IX7B//2LfZqblftQ8+81P2bO/L77aPfuLv2o8+MWDXn3vWPv6rn7XXts1OPfIh+zN/6t12Ibdgv/L3/qp9379e6P3E10xU/IfH7cOPjZrHy/jHh3/sJ+3D9qz94D86vBKzli19+Vl79trXdZ/4z+7F78+VvNu907Z8iWITOw465h1YlxpXvsMOdmhDotvdUF4gR8YnD59AD7mW374O6YQutyTvEhEiIDUp4F3fG4J1I77o6oG2GOBsBvIjYWNjY1qMkOvy4HPgZwPiUKMCVvkVgPV4zLmEKiEwhj89O4HNB/acdct9lkN430HXdrY27cF3XLCpiVF78SsvWPKgbe96/DF13xBaA76wtLwqL9lqrapNmaKYkFP8R5NpJGSAuG6ZY+r0AhgCdOyKfIjAmdu9eIgiGyud8jE0mw0omgpojAl887bxHigAEH361Gmbn58P7LmTMyymjLk67FjoghJDYKfuxYG6tNgcxbqyyHJfBH75Jo8tEJufpNBBZs4iihKi0a5rk4JJHiiVJV0sl8o2NjIi5n1ufl7ADgQK2QsAG14QNDSnCE0SWSGigg6LfTt27rze11FwlLkVyYhIFMSiIn6Nwofx5do1FwNBcDtRgaTOiSc6IznsDUlRUdSYckgrDSLRTGkeselCCrBpxOuKFgVYP70dURF/fyyuYoGhIqJZtSuXXrba9q5lE8gYs5q3KJYoRgBgAArZ2L2D0OWGqJpkDaXOSScGi0X3TeSD7sp+QJKJQ6eYQhcR5gbZYgSguJ/c+xjWpGsVd+f+k3q/gC0Zf37j+3e7KDotHIzjdRkfNssIYEjppMfJ1QgRHFfXo0g2t37qdfIGUFvemxkOkszdrlV3a/aZz3xW3ZAOSN4eZtsPYB1dQOMcip/va6I9Yt9yqKiIwHX80yWWFDkHlkunbWRw0O699x6BCXUUWQcdGx0f16GzdZAUSTE8Oa2i7nc//Zv2e7/7GT0frD8xo0JgIhcVpZtHunr1pdAdqyJLlk8hVJmMin2eHwcWb//efqDQi/o4BoxbGwsirZqhi7aPuLlt3rwNYBzncrwH/c9ovBYRIiG3JV4bhwE6M1njmSvlUsmGSiW7/9y0/f2f/gfWyQzav/74L9q/+fi/tcbuhiX361q7o+FL/z3R74zKAoF8/h5ddYStkRMVEXjrB0R9uh7mf/TmhUsqXIkgviKAvaHYj98XiYr+ORhBY8m3g/oqZoLoa/IT9Z4k9X7uk+uza0889qj9uY/8aTt3bMquXrkiO0M8yLcAPVFZFYu22W7Zyvq2ra5t2cLyqu3uNaxD1yskN03G4dmL1k/Rm1+MeN/civehB0aGMTicW3cmKlzC4QHeW1sbspeJa2pUA0VgPM6ffqIimKgekkFh/CMQ7XVBj28La9jtNj/9oHp/Loic8BKHioo4F7kOACipAgKhcxTkZvwOP1zCztwRUYEVoSWtNDxmf/6H/4p96td/w66+clHdYagt3o6ocLsrJyo0z1xS5M9nz5bOg34jeaiDCN1sfdcT3wdjA0iezLrykY/+5y6OYSR24n05uuYdJS20d/lC3hsCvueQqGhbIhAKUm4GtaDuK/NOocaH1k+671IiObkWnzH3kw5KE6m1nGCjVllfX3+LVSJAf5yf/Xk06iW5A1GhPYqmCz0PUdXrBJlqvT+AqAiX2huD3j6tNSplgwNYwvidvO/eB+z6jTnbUme1qwU5vLIGu+US1859xQYy7Q0sQd3H51mb6GwD/JVKIOzhIhvUZdC1lNShTryxfvbmrI+cgA0uSAAPytlgeUktGetklMbcM7rwvE50ogbrRs+j8ppT+y+/I5BnPncOCdjwQ3330tfY3noZVDRxznk+RVpNCJXKgJUJTz53TsCDi2gOVddafxMJWSdRl/RnVMS6yqenq181npCDSbfpYq2jKYnaaBNFBarYlKSWPibB/pNuWoiKZDqvWuJYAhulgt24cVM2SDR5rKys2flz5+3UyeNWrW7blTcu20MPvkPv4/jscSkq8ArHBunhRx6xlbV1u3zlTTUuoHIulvL22GOPWCp1YHvVXZuemrJLr1yyWrVqD77jAbt546pNjNH1emBT0xP6fLkybJ3mvq2vb+nskC+iGscale79QzJicWlZRAX3crgyrKGn45YufuYA3urMHScrGmoyQqXKfaX5aHxs3Gr1mgg2Mhw4J504ecYWbi261Qa1cgaAqWXH8NM+PmXtdsNJggY1GsBTydbXNowskeHhigjcra0dWYwwJjQvlUqDIhN4DrAuK5ZyVm9QVydtY3PDvuXbv93KAyVrbG8qTDWhMw42XYCCdLpWbWpmysamp2xrfdU6jT0rFwoiBuiuRqEvSyYzO3P2rGoxXgOlBV2tADOoRnifAmmKZdVb2Ewyn1C5WjZv1xeWbWV7x3b2sAT0OckcozPaG74c7MP2BJIEq5rx8TGBb9S/jDnzWQ162A2rEYh6OyFSCbBPYFWtZlnmHONY27WRctZOzIxYpZCxkcGi1fZ2tX4ur2zYxNSspXN56ybStrm7K+IrV8wo06/d6drf+J1bd4mKvp367l+/viNw/vonLZ/JWy4zYOPDFdtvkSZ/YA8/9KBlUbB2m5ZJ7Vu9vmNrW9s2Oj1kA+VhW9/ctZ1q25rthDXbZu1O0vYabUsRSozfP7mMPIdRoRzUr+wfrFXKWcCHv9XU8zg5OeGKeqklaXRt65xKsyBrs8qq0DgGWJ5Jpmx5acmVZONj1qaZlropZqZCkOAYUW+I8AVnYe9hDRGQEyyV2HsBirlO5T+g/hKG5PaEqDzSKc8vZR9nT0UlJ6UDDiIBXGZvon5gTebczuten7vpTbXkp+pXcjbwTAiFUbPA8W+pg/1rqEhY09RsRH2gBj6uy5tIwHDkbsB7lX16wSYmPMPIsQOvqfw85gC7NwN4LpZskgHBqVfkn+uWqnM3b7jzBAA9GY1gRVh4csZCcVBrOM7AtosKgmshh6NYsLHJca2JywsLCtRO8037TctqXYXkcZVNl/PwAbUW53xqETDFlJxEqFf4new3NIzhaJKyro0NFe3U8Qkr51M2UEjZz/2vhy3mH/7eJZtbWLfdRtsslbU2tQ3rNLgCVk80W4e8QZp5GTdIfPYANWlyxFejiZM81FTgD7K171K3J2yMvCTZX7vtvUizGqobb4RFTcfRC3zp/Hnqn6bsm8DYsIuk9gX7hFyCuHjz2g1LpPPK0+D+Ndhbcjh5sK+4LS84IBaw7FGqh3QW8HowWu1jIRw19TgXkNvUxkVEjYnefDc8Mqx5/IdXUfGRn7W5nz1lz/7cun34L2bt57/lB+1H3gLovx1R4QuvKzIG7Fc+8mH7vt/2z/3ov/20ffSplv3GR3/I/vg/OyQj/Kvvtn/86Z+0v3JuwX72237QfiL8vq+ZqLiDQuLnPvNF+wv2q3+AKuPru2H85/LqD8l6yRdVHkSRC+QvsPGwkCA3lwexA4jqrs64XQkfAAD8jFhBwDlvKnYvQUBhlAFBctVlUUsRylzWn2xKWmSVS9BV4UbHTq2+G6xkErZXr1tB8l/f0HwRZiNwoFUZPCTfhy5DeeqFDlp9PnSd0g3E4QmAVPZO5EqkTIxovVqzpcVVm50ZtPvuvdfOnD7p3oatlqTrM8em7Y03L9vK2ppNTh+zweFx+8xnn7Nmi+BFOpuGZXtC8BoSNg5T2VJWKgM2KPe7UwCEByYRUJ6CWcX7zz2TAadZHNnUYc1lMhGUEWxkdB6wEbFBscjKmiiJVVRev7tcLok55x7SqT87O2vr62u2vr6hjV8bhTrnffMBbJG1l4K/3e+YcSVoisW3wy6AXZ6+L2ntZtOl3/i4yg+vZJVhD8RjQZV1WM69GGUh1arp8I2lCIdQbJ94XQ4702fPulwzdDIzj3ivbqfC4Qbve+yQPOw1AoVsAgp0ChkMEcg5VFTgxRggTjbp/X11LckXc2zMiYok1k8FefyhiMkQal0q6T+6JujsYowjYN6EwQ5FQwREfdwOiZIIgMRDvZ6dxrbduHxJBzcoPoLB5AeZ9k5o/gPcYC7029owP1MZJylcHeFERQR4pHbq64Ll74BChIbzfB0lKiLBwHPA+OrZCOoMzxV2NQHAQATg5JkcAFI95HqOs+p+A+hjvsRiqo0tBUQLRR3PcyArIaYolBRSz+8N4aGyI5MtUkJjznM/d/OWvfzyq5QsYdxdiRQ/BNRF+wp++g42Kj3wLvyY+n9v86+/naiIr837FCELmMpzm0zLl/K++y44UdFsaK1g/qRyRcOcoDQ0bKNT03bt2g379L//hK0vL/X8lLkOPFUjUaGumjtYb/SD6brXIjfdnzsqKiIRFt9HvO/8bOxMjeBSfJZQVHCDRR65nKA3jl8rUdEP1se5z4tFoC3mYnANxVxe4LEIaADYUskGSkU7d2Lc/v5P/bQtbOzZP/kXP29fef556zR2LYm1lezDDm9mP+mi4jIAwgqZlp9+IGlATAWcuq1J/LMfrO7/vE9hJyookCnmkQf3lEHa43xMow1cnE+9P8NciuN+SJCyJ0I+MtpOVKQOOlar7trpk8ftyXc+bPefPC6iEv/TpYVbtrODoiIpH+3NdtMWVzdtYXHN1rd3bWtnz+3GOE0ImAOoYj92Yp7ObUAoqRSC8qi3LgXAuZ9gcMVdUD/ElHV1fLuiwpkiJOEAVBs6uPTPzei33xtDjWXwtA/d2lEu4LfSCTLWcD5iA0NcW+L8iZPyKOgewXS/Bh6FqKjwexj3drrB1HkUrIbi2hbvyyFR4aE/7s/r+TkQFQcU/pm8/eAP/2X7zG/9jl15+SXLqqt9X8RknEuHcypaYB2qGfoJMp63cB7WGhifWQ6W7Cc6VAfVROQs1KlHblfOD5xxLOLP9s/BOP7943W4J/hY94Bf1jPIviNrqLrWdfBsG1la/YoKJys8TySV4eADeepKHh12U9596NByn5WQ+9uFOeGKCt7v1uam6rvDeePhk0evOYLaUeXH90cSQ/WKOkwi+cjreVD1V0NUyOItqF3613vVGu2WNWq1YK+WUY4ASgr2o/0ueWf+nn0fcSDD8yD49X4d0k/pwBsUOxw880X3F+7LffB7g6LC62mBJbEZJVyYByz616mxpEwJVlEuvvK5T8cczQs7EHWa/xzW3SKO7Jt4H5nndAHyfvqf5944KNzydtK7n6iI6yv7kvLqqAkANgDQBwqyTT158mTo6lQF52RdWLNjkClgkWqHkO3Tv8bHa+F3yBZTlmNufwGIxbq3vbXj4aNJr/dVX9IBCymTz3gdLDVLzo6nK9bZT9jK8pqy5bBCApiHUDl/5ozduHHdrl2/YY8+9ohsIk6eNndydAAAIABJREFUOGk3r11XDgbd8vfd/w5bWF62S5ffkBqDTIqx8RE7e+akzgqQBeOjY7a8uKRaGHDvlVdeslIJ0Kpox8+csM2VFRsaqFgdD/dqTQpsOo55c/W6W2LSRFXI5WxzZ8dyAOc0iZjpuWFeQF7QYFMZHBIRw7OEZ3m1utPLcgHAYAywYSJDIpcv2O7unhqgsJwid0F76EHbanvbdv7cKTs5O2U7W+s2PDhkg0NDlshmrNVo29VrN21pdV2vwZx+7bVL9q7Hn1CQ+fVrN+3EyZOyQGPyj4+N2sbGqn7v1NSEXXnzDfvAd37IirmMGrU2V1flCc+DR3fx1NS0DR+bsfr6htvUdtu2u70h9fz66qrJfrZatfXNHdn8njp3zoaGh62+s2UdKfo5ezRsZ3tXCgmuQZ72O1WNoasEU9ZJZezGwrItrG1YFSVGrthTuJEvwTNFXoqUwaWi9pZKpaJ5QJCvzoUJGt78HNtotPT7vOvZn/0HH3xQRMfHPvYxo0OH7ujZiREbHyzY+EDWhktZGxkq2/U337TZE8dl9zRQGbXiwLC1ACAzWVtbX7OmwrSHLZ3P2n97N6OiV5/+//uLK5Hvfvz+I/B09YuW6CaslCtZdbthjRp1QspKuYyVC2k7PjVqD1w4o7930x0rzYzZxuKq3bi5ZDt7+7a8um2N1oHyBvZq7AXDWmtkZSR3Pq+dwAcU2hyaSmITn4DdQAwALg9PjFt5cNDDoQkrrtbcTjzYtYqsyOe03m7Q4NPuyBacnAdslsqDA+qoZ6vnfNohNNkObG15RY2SZOrQMMc6x3VCnKYzOdvbq2vv0FlLFtpJy+b/X/beBEay7LoOPLEvGZmR+55VlVWVtXV1V7PZItmkmjJJiRQNS4YwWiFAHg9sDixBY3AwFuSRpYE4Y9ijAUYzNGQbgiVZMgRpbNq0BWpMUhSblKgm1VtVVy+1b1m5L5EZ+x4xOOe+F/Ezu4pbczz2sIJoVi6RP/5///377jvn3nMM96InDcFjPvcC6D22JbzLCp1Iyig2OCUPVrgzb7m3fF+xxPYW9B4d0HG4hjEXpBwRi0JNdcKkDv0+T74JrvDSF5pw/LjmMhaReOYgP/bYY1LH4DEou8uuNuI/jEdcX1gkxvyGcZP7HBIzzAckMV4pa43Z3dkRxqJukqgpS6gYimu9vC54fCcfzmtxhbO8F+x64zHyuW2NN8lkYi0ca/0d8ZtEUn5C3GeYjJQVY7Cw1sgiw/z4Im5G2ep2vYbZqVE89Y5zWiPoefTvPsXqeHv99R/dxv21bdRbIflfRKLs2rBOZN+No8LbuCmT8Jq5zpkPqxERHtuQ7LDzQOL6y/Wf84frBD1F2PlIQm10dETXRNyFXXfMnSvFgrpt2VXKvI74GmXAxsYm9VkcHxL6JOPeuPImalTb5m5c/h1FZIeHde7Kb11OSblgrk0sCKD8FHO/1AA7VKxAnPNH5Dm9WopFPV8qRJFjmqkosMCB8/W7lqj4+//hz/GJgT/C0vdfwydf/SWc/Yufw9LPvnQoIn59ogIXPoEbn30v7nh5pe/7BG784UeAT30cSz///IOj6+JP4/Of/e/wzNV/jsG//jt6zyOi4ju7FJ9OOGCfVdWsLnfAloFURgSoktCxkG0nPaOHnAahzjxQlVUiD0yGRxsXGWk6rXFWrceYGFfwjgsXsJ/LGeNNfV3tZiMywyYwqIWpVJR/hUnJsA3e2GbbDFlOIvaQAKlMd82E17O3Rg4QDLdg4M1QDZiMuGpUqAWOwDt3fJViUezuM888hbHRYbHORB+oVzg4ksHo+BgQimFnr4jPfu6L2NjKIRpLabNIzpradqwMZAAJRckAWNWljL4jEWkBmga/aeXLXMeBSwy01bp1L/jNOzdlWoxSAyY9ontjwJwAIOdlISJD0j6UYSE73EGhUOxp2nEDxGScnTLSHnYpncgdV6EmXwsaW1FjPpnSv5T1YTUjj8/JIKPkuplk+XY1+ZpwYRaTb5V0TMR5LclEDJUqJV6ss4IAKqsUR48f0eLrgUIt1K4CUbObXh3UpnT3mZ/NwM1xZCWCVTV7vWgjOdhP3u4ae857QB8NGpRvrK0JOCDQ7HVrudHxbZ70qkgPDwkA5HVz3DheZpoaQqVZcyCXk5yhmaQzq9U070kr9Ku41R5e2cetq69pAWOywE1Vj0xj1SMXTSftZI+IkXYaQ8qUqeWTm9g4qEco9RAu6NKMccCrGx+O/bVr17SAMfkybwojE720lweIfPToA/veZ8Z+0+8KsTnmpRg4XpojTj5EgIMSUwOfCL7x+bZOCgI+TKqYjJDIIElirY92DNMqJUlEgOGrz7+I7a1dk2uzwsleBa2dZ78C26izvtzHYeCjl+B5kM7JXNmgHazktuoKu06TqLKkJzuUVTJIM23O00qjJmJrfHzCWlVZPRuJ4OLFV/HyKy8bmcvD+04V56Fh5ugHgfjevXPj58kHP+4GeNpz78/HgCrfZSM05wD54SViLN5ZBY+AH6cV7u+5zseBpSJSDlVcB6VmPFgqkoVX54B6A6EpFWTaziKaO221V9dKFb1PyS7194fYeZXFj//YT6hy6Ld/519ia3vbgXDWrh0kAd9yPoHOGv87T956mZE+MO26gdQb4IzrnearwDuC8wLsyRcbAOpJ0OA96d0Hd508P2tr70uP8f3B54mfJ28QzXDiqiGEOE86wNHZaZw4Oo/RwQxCrSb2d7ZlODo1PY7Z+VmsbK5jfXMX97f3UKjWVQ3KCmJ+JhN+I1Cs48aDs4pNzh+Gz7ff6Pjr8ABxnzi1tm0dS1XXpt/t54uuORQSQV6tFGxuufnmY4JCjSsACMq32By19mMD2w1E5iNrcdq0coP31s+h4M8PgKRuwpqWq3UV6V5x4+T8mrjh6jRtY+avI0hMJiJxkWD6j/feVelSMoQ5jGSIIhE89c6ncevmLbXBcyvFzZSXmPI5jDObORh3D80B3ntuGBh29FmMjewAdUbSRsj1yQMaK3P+s3szmmTnmnt2D+RfB8fN34MD8f9h6SDvQ9uRHwHSlmPKmExDcY6Xlx7s+2+Y9xfvp7XT9w2SrWfCvvfkRP85kDOZ5K7MfNDW4uArSHYGv7YSQ9vY+3HQWuhl3lzcNh8E7+VjclkipALEdfDz/Ll5lx6LZVA+QCCYm1IPbj399PdgY2NDlXHsWiThKNBcXRvW8Whmk+pvsMpR92FWMGOEWDSeUC6hggPp6Es4wRU2HJyvfG595415sbBqj3mReXnp+VC8snXLCIcIBtKDyp1qKihpKf/y3jl8D4liHpfAthUaOWLHnXdAh6x33AP3Q+m4rTHBzkxtmmn6XCtjZHRYG2PNCZ+Q+9F0ax7zKObx5jdh4yFvuUMv67IwTycBGiyMcB2XLMKh+amIZWfoyXHxx2QuRylWVsTPx2jymcad2/exvZPD8MgwKpWiCBWC8wSoX7l0CY9feBypVAKDg0PYWFnF1rp1VJw5dxY7uRyu3LypTicCQHNz0zh6bAGxCImEimSEVpbvS5Zofn4We7ltdRYkklGcOLWIfG4PQ+khHY8+D6ywnZlfkJfG6uq6qvKHMhlJ6r555SrmFubVec3rHxkhKFI2+dVqVcVGNANnYdj01IyAJ3ZsMAdjReYwQZRKxXKMUERdCceOncCXvvRlVbYKFOqSsCrh6Xc8of+uvXEZE2OjIh7o9zCzcBT3Vjaws5dHPDmgrg8CLcv3VqzLl2RAx/JCyqBxnnJvRICf3YHRRAjv/9Cz6LCrnjKz+5xzBG+q2Nrdxtr6GpaWTuHk6VNolSoiSKNxku4tFHK78uUg0d9odbG8uoZTp89prLotyp9VRO4R4NtcWUOU3eraQ7JylnOE5xZCIplBvdPFa9euo1ito9ENScOc81xm2OkBFXMRmOP3TIOarToGBwc0Y9V1L1UA5ssk+6Iir3jt1BVXfshK4GYT4+P0Bamq0+L48UVcffWSpJ/On5hDJgakYmHcuX0bC0eO4PbyCmaOLCKaSCNfqkgVYDA7iHQmiWgihnyphF/4i41AJHlYMH/080cj8PZHgF0NFzafw1h2FEOpIYyNTGBna0+k6tFji6iVC9jb2MPcZAKjwyygCOPI0lGEEyns7hSEe+SLTVTqXVRqbZSrTZHd7HSKOsWARqtuHcsymWaFeEjPK6vxrZiqLXkdvmcvv4/BsRHMzS9gd2cXY/SecX4C8nRSZ54VvXI93draRCIcE5g7NTMjFQcW2bFAkmCxZOlKJeEOccarUkl7Pu6l2JnHGBmLshC2Lm+cZpP5Gr10jCRnl6V9vuVtPk/1WFi/yIK5NKXNCYi3dJ3EbyQ5JB8BSl7ZfpfrnuUAkF8Fi0cZYxhXmIf5jlafwxJHYxyybgoW2qpKw+IT1RISCYHnxHN4fibvZPiWOkm6XRVgsDCy5kgJ/owAuqSjKL3uOmR5b9iRx303X9yXq1BL3THMjcIqQrU9muGE6lycndXnba3el2QT7w1VNFRkQQJHnSJx7ZX5b6NJ3IlkRFRECceOeTyvi3sydglyPeAoTU4MYnJsBMlEFEsnj+D/+Me13sR/57NXUKrQG4XdaIzcYdSl/GJ4Hsea+wTOF16jVwjxha0+J/U5jRWssLjTOkVJmFQrlD3vKC/nPpGFrlx/udYI42J+omLaFoaGMyLrOQ9J6tPrrFQoSzo9nYhjcfGIfHY7EXpytoXncM5xHaG0oN8f8POZs1GSi+fB3M17hHKfzRyHEo9+PnL9oaoJu5OUM4e76EbMr5ZdmN+dRMXi38OLf/bDqP2TZ/HsrwEf+Kefxuffdxcfu/BxGHXgX99ER8XfAP6Z68b4qd/9v/F771vDr5z8W/hHXycG6/N+qIhfX/gZ/MIjouLtr1aHjnAube2zVt3vq/oIxNgGxEu39DbHXIQcQSCA3n3tJZ/U7UCm2FWdt5xME1lC6rtlkkmMZLPShy0W8tja2RbTLeiRZAhZ+Ag19AJAmEynDfAwpMnAbNvgWNUpg61V4hkAJ3LCdXXoe1fhpmBKrwDyCGo/ayrAkykdzKS1EeCC16y3pTPOgBSPh/HO77mAdCaNRCqDwaExXLr8Ol5+5TU0mwQTQlr42J7FTaaCfrctgFma+2zZc61dviOA+rG+wpKSTFwwTLjciAyBjM6Ekq13pqfIxcIAI1VtwjoruEhw8eNmzrcASrbHyv9MH5LgJf/n2/9ct4YqAsLW+UJTI9vUGsDK8SWoQxKErXRcVGhOzs+qV2s6Z2OyzbyKCYP+FExkWN1lbZOs0qWMFEEMJgXZ2SkBnVrMPdAlYMykq6QTS78GL6nhwMJGwyrSVH3uKuD5gUogmJB0zKNCbZWStLKqLV7P8NiYOlb4YhUCq9Z4v8hapwYNhKchJhcBGiv6FtZq00gLzTVWXxAYMIF5kVMeBPHG6QLAmJxV8thYuSdd43KxJM1+du9InosbUy2srDQ0IyhqbxuwSLzDNkdc5JkgJJWUhA1kDBgD+0eZY7W5sYl7JNaAHlnhdaFl0O6ASf83HkSyTb8RkR6s8ABnkKjgmPF9QTBQOpuus0lG8NQxJsDq9PxbbVdBSJMuERVGCnChJhhPXWnqQ37lz7+KcokVBbw/fRCM58rzCwLoRjaY1qmPSUHAU5Uheoj0oPS6Ryx2vFVyxoMxTpJfn8d7tbS0JICDn10ol7SZpa4qW0WZNCwv38fVq9dU2eqJFPpB6HMIMPN/7BE9BMz0ACFHVBg5ZSSVlxXyFbf++hUaHXAsgN1VNPuY5sFigXwiFfWXhzpK3M9ch4f/Wz8fPCAf/N6P74OICiZUfl612KFAQpZttmLUwjI65bxNJWL40Ic+pHH5zGc+05M80Tg5YuUwieavW9Ji7j8/74yoMEpAwGOgo0JznLfePHeNXPDjJpCTcmu2jgTB8v7aZrHk8CblQURFENhjHNaMtKmrMYgwZHMdpK53KoaBeAxZdm9FI8ik4jh+8hiy2SGsbK6po2JlK4d8lfq/dRTYKt+hYb0nP01yyPRW7V+uFTJ4cxU3vWtwZKOP337eaE1xcnKRCCvlTYbQ+wbwfdT8ZvWtH1ffTeHvjye3fCzpA7QmQ9UHpllpbgTLW+RmHODqCYb+3HVSRQ7QtzjQlhyM1ginTy8S2AFhHVXnWZeYP56fv4lw3EyqeT88UcF1gR1yNCp3QOxbCRIjRu3nRg5K3869gu+3bhX7hYgK1yrh54bPO/R7WxhdXHJQMSsPkynEnX/JgTj2AO+NYDw4DCz3TtB9oVNxRIXPKfivgePmFcWz9t06ZrrsYgvJcrdZPkxUhMLcDPfvte+qciOgQgSCgVzf33JODyBte4P3QKLCZBlZLGHz++0RFXYQdpB6ooKV3/Z697vfLXD4ypU3jQCR3JLJEPEl43kVRDD+2Lzy98NurXU5cQ1j5TSfyx656AytOeZ+rvp42yMqCJhQdpU5ktZQan33u4g8ucrniQbDPBdLn7q6V1acwK5NO2/+nN2srQa7Q61gJuT8Pb4ZosJ3VHjCSCAJi386HVRqJQyron7aCClHJPoYLR+OQFdRkDB6IFGhqk8jDxWPnCm3pDNcRbtye0clvqV2umsdqu9avIBUYgjXr9/CroDmJPbzOZw5cwaTY6Mal6vXruL8E4/Lk4fdETTFXrl3H9VKHY+df0xyJ69dedMqVfMlzM1NYZ5G0PGICnRYZXn39l3FpKNHF3D3zk0MDCSV6y6dW0J+dwfp+IBixt0797C7l0cmOyxNacpQcV8zkExJt3x1fU1mtQTrfay9ce0mnnzqgsgKyZyMj6kTg0A7x4PVnkyMb926JZkk5lEEyghg0cNhhibOX/lqzwcvxGKRZhWnlxbxPU8+gWtXXhP5sru1rRRp/ugJfO3li5J2GRoZU8EX92NDg9aFwJ0Idee5F6EJeKtB6SlKyJJsYIdwF9/3wWeVl/KAOxubGhsSGQRsSuWSCuDOnDot+Za93A5qtbI6KgbSKQErpUoVL73yqjTv3/mudynPKu7vIZ0kMUYT+g421zbUhcDuM5IiDAmMQ3X6ydRaSGWHcXtlDblCAeVGG82OkQ4ExkjIJOIJ7O3lRDBFo+wQYsEMwR8ClATNzECb9yGdpFwwJaAYIw0wZCLJXFeVyeyCSSTw2PlzWL5+FfFuHcPJiDor0vEo9vd2VfG6trWLiek5DGRHsba5hVQq4zzo2khl0uqc/NgLm8jWD/rsvCVwPvrBoxH4DozAeruGD21+TV3j7XoX2UFWhHPdj+Lk4jEMJGMYzsQxNTqEWmkf23s5xAei4NaNJEWx0kKl1kG5RmA/IUkbL8mtONGk/4J5TXAJIFnRbXedQoEVrtRqFXWH8fljV4D8BWJRKTkQyFeu4lQTBNKSDGBBQSiEjfV183uIUIaYhZc8j7Ak+hjbST6vraxgbGQYk+Nj6qqo1yvaL1LOjnlvNjuq+EaJavn4uJxdHY10GXfFDFSn4MsK8wwjkQyfigCsEIxfq9iNBtXsJsvlemtwkoCx279KmURyQsQXjCiQByy7PxzhQYLCcij7LOZdvH5el+ShLAFSnJqdnZMHhXw9ZKBt3dzUWxKm1WzKC4+dIfRII3FCMF1SV64otEo/Usmgmh8mP1++PvwsSgoJOwub9yVxJ5iUOk3FjxxZEJa3s7ku4F55JHPhMN/TkM8R54N5f5CwsL2HLwJKxCmFZB0NxJXMk4gFdi1kBhKYm5mQFBQNu7/0x0d7M/+9H1nDfoGYUxf1lpEhXAvZAULsh10M7FYkRiPfRF8ELEk/I5FEZjjpYj8eIipYnEriR/sDw9fk6+EK75TrWZmOJP+IZY2ND2N6ekr+FLU6u1sGVYBQKZcxnM1gdnYKV69dQ1udKhxXjnVMpI1UZ6SuYkobHEWanPOcvJS+EVGmIMJ1mfeW94Pdfuwq4lzi7yNci0Nt5WPHFxe/O4kKEQUf3u0TCou/hNee/0Hsv8VU++FExZM/+Qn8q3/8EUx/7ZOY+Mnf18ST/FL99xH7/k9+/RD8o7+O+//kcVxxnRiPOiq+AytW4BBH0VYSx+DkNbgZmEw3z97o9dwYkA3wY9U6NfaMAJDGLE2PZApnIKu2Rgq4NM7lwxZBPBJGrcyqpKwC29TkhI61trGpZJzdFdTiY+LNgKmqe7Xdu8puX7IqIM5AKgLSDNRki1XpT/bWge/82sAVqxwkGK/FR8HaKoXJqAtcVWtcAtM0aorHcP3adQV/LgSxWAjZkZTIj6npWQxmR9EN0aypLE0/6uHSEIgL5VBm0AgGgtuxuEzxeB1WkUt5J461dXoQ5Lxz944qodgGyYoHC4iUqTK5DgZfkxmg+avpBPKlRNsZQ5E44j2UrqEkdQZV1Uhw1Zf9KWmvVU3+SG3mtV67MzfIHDMZBSVp+mrMrqQIqJVHTWAaDY2MquqAx6KpD8+zWCpoHnDjJ9KKhs4RalHS0C6kbgrWG3NTQB1KLigDo8Pu3ppOoAcOdd8kF2Emsr1iSQdE0djbOjdsHnpQ2gAEazsVqOoIGiPHLDFgxYcRbEb48GcCE1T1a2ZWBBZk1k6BRXecdod6mU7qxFU3GshrXQS+jDoIyAliazdQLhessrFQ1OcOsiuB1xU1o3WSa+yAsYpmA0KYpLCjwpIZVj9HkUzTR4a+DjFQQMRLrFhFqcl/sYKN8k+sAOAmm3/nuynMSLuv9e4ffw+6GdjpDGJ7lZt94Jz3l4khx8/fKyOHqEVpoJ6kn9hCqvGzKs5Gky2T1mVlEhQGqJCYE1ko0Af4i6/8pcac5vWG5tl4PwiA5A5VPgAuNvn39QBtB4DbvTGQk/foQUSFB3V6BJEDVzh+NEM8ceKEzmOvkFc3DmUKmODykHfv3sNLL77kDOTtufXG1QLrXReEdTHYKzjPrTLX4meQGPJgcBB4DY75g4gKf2xPknhgyINg/c93AKzI5kOk06Gq96/XUcHjHiYqwrwl7AShzibnLjXNqSEej2GW1U+lkiqWDwPDVvHrPSgCJtZuvPx99X9nyZtpzPpXkLAw8137neJJgMyQVqsq/22uB4FhT3IEiQo//x5EVARXYU01R47wXz4D7KaQrDrBR9SRCIUwOzyM6eEssukklo4vSmJxY28LK5u7WN3eE1FB2YoiDejYadh1xInICSfBI48O8wzwJveH55Z+7yrHffeDjYfFFCXLgev3849EBTsqguOqsbJ2o97fGFl00EdG5BDjAKumuSGIMq5ZFXW/rr5PLvY6IUSc+3vRlwayG8jPdhKBrmuJWrs2/6ryqLDugL5Ukz/3GKKOqGBHhXU5hFnFRs8holyekHfzzI8Bj/fNEhV9kN6WgY4WrD7hGyQqnGT6Qdk9yaTFkBgw4NnfR/4bJHIOzDWXI3w7RAXPxxMVrLS2NdBkxTxRwXWGa/7DiArIgLm/DvTnFwme1gGi4vA5Br8/8LuHdlS8XaLCcgl7+XhhG/O6tP2ZW9nrwoULWi8vXbqkYgHKGQSJin7HYxQkZv1Rg3FJOQEls7hOq8ggZnmcl15jxHe5jCejezFa5JERFSYLRaYzQKg6AtJkAu34XIs0jwPkajBeMierV8vW66Wp6Qsres7uvTh5+F6J6A108VkhhyMqGiZ7QDKfOWd/rlrRkApr3MsXGSj/oISEKk3tpTXGpVryK3KdI3YNJrnln4nDMTv4PQ3dCVi9+8RTQDeG5XurKBTLinWFwh7Onz+HbGZIQDXliGjszAKaUyeXsLWxieXbd9U1cObcOWxsb+PFV14RaEZQe2pqXMB+ZiCpboeJsTGsrW6o6pL+Bpubq+okyg5nsHjiiIpSUvEUQp0wbt68I63veDqtLgESFZJ6C4UllcjujVgqhvxeXkbPvJetZlsyHpQeoRcDi2u4f6BnXjY7qHWX94XrA3MyyiYR9Ekk05JHmp6dwyuvXJJcKHPBZDKKbruOc6dO4ul3nMe9m9dVcUxpEJLiRxdP4gtf+gpKtQbGp2Y1R27cuoW5uQU0Gy1s7+xqrzA/P4eOqnZZVGFWT+lkHPv5XfzAD35A18M9zca9+4iGQxor5nm7+znJaDx2/nGU9/YlT0pAkOcwkM2iVSmhVK7izSvX0OqGcebceUxNz2B9ZRnZwQGUC3nl7tdeex2ZsVEsLp3Eyo1rOPXY47pnrXId91fWkRwcwr31Dazv5pDKZFFt2HNOQ3PulQTuCWBqYm1tVZ9v+u4GrvGJZixmFTALlpLJtMaVHh0EHTnuPA91jDcbJj3JeN+sypticWYcs6ND6DbrksaSHFUojIGhEYxNzWInt49alRr/NdDucWpuTvuVj1xcxdlcnzANxvpHXz8age/kCPxJfQu/3FiWmXYikpRM3vYmVS3YtZREt9nFxEgCR+dHMTk6hImpCQzNTKNeb2P13ip2ckXsFWrY2smjVOUzQBKDqwv3gdaNStCYJKt1E/AzWtqDc4/K9YjPImPdPOd/m0oTYUnyDQxk1CG2t78vI24CsdxvEjgmmE0/msuvXlZOSdWDzOCQuty5VSdBQgCX+AtjFAtOWSPmfVG502IHFPEg5i+McdznSxVCko6WfxKr0HpDmaCoyXIK6xBoHlYc9MWOJDFZAc91irFYZS3yYjWfT19QyjWNuTDXV+/fJSkpkhsiKkLCXMz7yn6mPNpJQlnHRdQZK9uafPrMacV9Lp7c2zN+sYCn3bACwGQ8jnxuV3LdjGlcT3J7e7oXvkODOwRKk5sPB6UXqXbR978kiSGEjAURzusiQ3krdkwwbrIgMhaVvBGvix0xLAzmLJDPj8zTOY4mecpCKx7HOk2oGMHztvFm3kXyOxLqIjOQwrTMuuk3UsHLz53oPQLP/lAee/my1i2XpIkwiEsVhv5JLeFw7IZk3sHCE5P3MvKHn2dF1NbJ73EvzlmC/ty3Kz9xeIG61VstqbzwfumekHxxcqCz89Pqytve2VHIIypfAAAgAElEQVRxbJzrvusSoQH3/OwMrt+4hi6LXIgFlkgWxXUskhRcL3veoaC6S1UkuJ8X/DwZr7OL1Xlt6Dw70DPi/dLY0Vlr1OSLsTC38N1IVPww/ujVX8I7Xv+HWPjpP3ITZhaf/MKn8Xdw2FTbiIoPDD0ktK4/j1/4mx/Hr7/K3z+O33vhX+Cjy5/ExI8acfHw1y/htfUPYP1bISoWP4Ebzwdkpg4d/JFHRX9AnhiyCW9G1baR4UNubVOm2e2DN4OuNm/aHdkeUPXLTu5BlWBtmtOY9h3fzweKJEKpWDCWtt1CuVjE7Mw0BlJJjI2PKYHcy+9hZXVNQD7N0RjgeGBW8zNZ5KIio1qBulYBLtBOVaFGpvA4BBmNPe13LKj9kEyv25iy8p8vvk9arYBYYv7tzRs3tKGh3jpBZQb5iYlRHDs2qRawRHIA27t7yI6MatGjfh0rq7c2twRKUQ+VhntcDJttVkDFjTBwCyAXBQabW7duY2cnJxM6jnG+WEQ81bd8t2BKRp/mPUwImiIqdI+cORAxUFZS2QLX1PjyWswYKYQRVhIlkgIJ+SIDLfmghBlp0+SOf6PrYos3F3SCyM2WtJDZicExt4WkiamJSbCrYXtzU/eUjDPN+tgOSKNBifK0yMwTECPNw/nAjYkRFUwI2K6WGkr3wGwPIGij7L1JSSYIPHFJgwMeO2EzJTVQxzazHqRUpaM6MKzHwVluaqx6BJtLJjgWvc4MLx/heiR0TGeaKp+QkC2mgjmCoKcvwdfP+LlmrimdemoRFovI7e/pGSBZxc/LDg4ay88EJ8z5GtPYqfLYdVQwOePYmeyGtbqLqADvPXs4fKW4PYec/SSpSGDt7e7g/sp93ctgNwW/92Beb7wCMdESK2fo5eSQeJ5W4W9Sa756XhUkvvqfiaTv0HEdQJ4845i02lZVqyTFERU8rjxT+HnhsAwnX730hhZfJi8OeXHJgsmB9EEUg/eDnREPIipkwuoVQb6B9BPPzzoabC7x+pgcUHaBQAzHgEQFn1ESFdzAchN+8ZVLeoaNNQoQFUFteD+n3bwJglqagwGw1I+3kWAHDcX933mTVl8G5O+l/73AG9eF5I/hpboUfyRobjfeKnIfXsl3+Fy9AD+Py2MGpZ+UuPI+yVPNbeJJAsZjAjZ4P3wC7uePv6eqvg2QOMGl2rimPszdP28vE9N/t0gJN3ZdoigOYPdku5EWfcksTwj58/DjJaN3t+b589I5OKD+YXmK76jwXicR00WzGBhqIBkOYTSexER6AItzMzh76qRi604lb9rau/vYL9eQyxdViUqgihWjPRASAaKCsYY7MecBYcRgkJxxhuHOKNlfh4BHSdgYUeHH04PNTJQbdXoLWUeaBz3tGbNOSv2NI4r9uAgAd8+AyF8RFCaPJjDVxfGeCXVgfj+IkHOh1jVXMc6biapiuvO/4ua0Lc8ikxSwv+mTVyIq9DCE1engpZ86TXYVcsPar1b3f2vknRkn27w73FFxsJY7SAJplh7qoOqBqb6bTapKtikWqak5FVZ1rT9W8Fk+MP/cxPPHfNg8VPeJcTwyl/TH8+Msbd4Ox8z8u8yA2e6Xj/W+UtF3evl/Ld8jSeGeIyeN1Ltf9KFq1pXfmM+TvQ6vOW8hWWSmbYbTAvKDXV8iHj1poB5LF25NXuvrST8Fn4l+jDHCjh2hJm9gL8Z2rnHr62tqbGXVtc17J23kJB5FArpiCm9+afmvmGnLHeQv5cgKSrbxuXOdvv6Z8kSF10pmNSHviaSf1JHg5EE9IegKLLgORZk3OCJEOYnrhgyuhTbm1PM36VTeE1Y6mqeGk88KkF7+b/2/HAR+7Ys6gh0b9VYVs/MzeOqppw7EZ821tsl0ekLG5x36nvEwQHD6Oak9B0EMZzTuu02CZJ3fd6igypE9vXPtms/a2clTkn66d29FADs7KqrVkvymRodHlNOz6/TUmdOa+5Sw2FrfwM2r15Ubnzp9RkTFS5cuSYakVCxjemYCx47NI51MSCN9emoaG6vrel5pBH31yhsYyCQwOTWKxdPHUdzdRSKaQCKWwq2bd7Cyto7RiUkz0Gy2sbK8gsVjxyRjd+feHczOz6kqkzGffngkg5hr856RCGEHBvcClKl69dKrej/fxzxa0lvhiLyyZmZnUSrXMDM7hxdffEUgO0GPZqOMdqOGx84s4fEzJ3HnxlUszE2LUKnUGziyeAKf/dM/Q6naxMj4JOjJRnKFOuo0IqX8le9Wpwl1Jp1Cp829VA1H5ueQ29vG93/4/Ygypjfb2FnbVFbKIqx42jweCER+7/ueVWFUdT+PerOKeJwGeG11socHBvDy116SMerps49hdGQMuztbSMQi6lAgYURpPp+/cD+RzxWsIzmewl6+hJHJadzf3ML2Xh7p7Igqb1W1SkCyQZ+OCk6dXsLo2CioB84gsre3q0I0nhcJDJH/baBSrolwpG9NUXJVJmHCMdcaQU30dgNtythm0khG2jg5P4XxoTQyiRhWVpbVxbG2uYPT5x9HG2Fcu34LE+NTAn/ZXc4SsHKthidzTfy1m/sPDeePfvGdGAHf936gvsUOHOSxe/VpB3+odeRgGur+9AE//E6c7v9Lx/jF3dfwH8qbSMXTmB6fxtTEDPb2ikilBjA3PyeptfWVuyjsFlV0lBkKY+n0CSRSg8jtV1TFXqq2UGu09TVhBvqKaj1ldb7Miplf2bjUaw1t1xjHhSfRi6fbwezsjJlLh9htURHGki8U9HwlMwN6xhi7SFCw8CkeiSsfze3sSsaNGBOldkqVshZeSoYzRrLQkl5rRxcWsLmxLtLi9OklKT+srW9o78biAXZSyESZMtkE1kk8ar01OaZ4zDAT6+YzOXRV6HNf4FQ9GBNFpMhnIqTuEJ4Lr5PvZVU/r4Ejwa+90TV/LxJA0tVWdOm7opmfc1/l81mOIY9F8oFjyrjDHIWYGQvnTPXEmZTXqpI35N6UmEc+l5NEET+f+FO5VLKuDno6uT0vSXvrnDBpSxIL7MBIEftpNIX/MH5z/pOYkYcGZZuEI4WF4f3Ahz6kmPqlL34R169fV+7kDdEZe/n3NUqfc9/YaWkdtUJd5lgsRrYczAiWKEZGshgdHVbBK2WlvvCvKeFnryf+yjqK5aqOJ0/NUFcFB4kE9zScWm2pgpCcEWbFbhhKljvJan7Pa/fKBTymFEE4jryP3neU3SDqFLWAQCLDsCbCl211BnIrND45pjyxRLK9UMZgJot2y4y42YE5NzONW3dvodUJKxdh3sg8m5J/MlkPhBl6GErCyu15ef6SKeztR03qnHmcCrvQ1bpoIYz3lR5itjf/7pN++vi/QPEXxmSA/TPOAFsj88Cffx3pp8Wn8Yn/5RP4+PuK+IOP/QQ+9vm32VEx+zyW3vsruPuwgP6x38D2r57GRe+Hceh9j4iK/oCcTrJKyqSSCMwzYfNssN+W28bANh/W4cuvzbuCL1Umq8PBpCnMiJtABwtLrHWW7c1s+6N2HuUwKCFEDdXhLFvIp5BKJxXkb9+5g3LNDKEZWLigMYnnoiJahIC02wxZV4V9hpexYKDlJpnBlYsAgX1WdRozbawo4SP+nhVHPMfssJEVDAyseuIrmeLnWSUmmfow6tJIZUCniRTBfZIUZEY5Lhw7BhcGWy5KrKjhZkFySc0W2GpnY+gZewOhCUhRf1CmSk6yyhuRSuLDl5wJJTCvCLUrs8ItFhUxYBXGYY0nx54Vd7w+GlARCFcAdmAO38vFj0lAs91wUkb8HBp2pxS0SdSQAOH4c6Mutr7dxsjwsHVZsPqA7DSN/5JmPMWKDP4rE0hVMNQkLzEyxr9pqZKImwIu6GNT/Jl17HiygWNtwIOTc+FcciQYu0R4Xu1Q2wxkXZW6ZAR8BaukdKyS2EgK+1fgZQAINULBXkpApafpgGb5UpiMgwcXQpQJCQDKvpvB/rZfIezbj4RXhEJY39rB5s62rpMdFdy8Dw0Ous+kLBAXdM4ZX9Fqc1OAdcyeox5RkcpoQ8rPUEcGvR6oDakEjXJfDeR2d1GvFmSI6+e6N7H0Ova8Zl8x7pMhq6p1YKJWTiY/lkDx761K1NpMLZEzM28t9o4MtMpI1/HjunyUfLTrJl/hOiq8sa9M0Zl0pZK4dPEyNjZ2lQBYRYJVoPIZCAKl/YhFEi7oWWFgdg8A6nVRGHBuuhTu9wFvi/6x2RFmklv+xWulTvOpU6dMUqFUVJU+W5YzmSFV6T3//Fexs71jT6cH/10lhjfLVY1Rz+cn8AGafCYHEwTt/P33IPqDQHp7f2DeuwfHQ7SORu5di5fh0vX2unHs14eP75+JHokQJAmcKSt/J6NWp53JcxXppOy/o80BAWJWZFM7nWaYVsVtcdJXjvtr7N2bQEeHACjnJeGfpyDBYafVNyz21+Fjh2R9NNdNZ7YHkHNuu0phI+dMosuD1p64YVw+ECP8WB0iTXoxxJ2r76pQbOP6qMaPLrrhJtIEeUJhTGcG8T0XnsDi/DxKpTy2Knnc39jG6s4etveLyOULAogI+FpHhZN6crpSXk7JqxH57gY/rr34KVLCJMWC1yIgNWzeInx5s1yOBUFSmp3ya2nOHjCjtw1IcI4ceO4CRIXWra6tu9qgOXzA34cgeB78DH+83mfwMNxAct1kjkIwrMXcwbrz2vXqAQLWX6eS+25EZb98xjgf1eXIiil2fDmiwr/fb0JsLI2osNe3QFTwWWZlXj+M9L7yYUjzzH0js0j3DsZBxhn/TAafy8PP6IOe2eBH9uKaGl/7ZxP0g7L8zRs3MpabsbriLueBkz0SqR4wmTeQ2zoqDscK42uNqGAex45OPV8BAvHw3OkPEDt0+5X5/n1euk3svOsIsu4bIxssTvW7Y3rA9aF74J8JH0N4n2uVqvKXA8+GKzrgdWeHBgxwkJGm6XALcGHeE+poPhE097maO0Ot035DaiSQJ+5IgvXvB8eGcZTxWTFaeTfjJP81MTnlWtzQupxCXZI6HjtBnbQUCQX3LPM6La+ydSWTSeP0mZM6NQLHud195PMFVCo1FQtwzHkeKuoJyPDpvh3yqPAFFlzQGu0aZuaMqDCwxXUDcc12XRJ+HmpDHiCjD5um92IIZTWd0bgRFX2vGD+PrAO6T1T0n1+7H8eHjiIaSWF5eQ2b7F4YyCgfevLJJ2RMvZfblWfCydNLypOnp6awt5PDres3BHifPnsGW7s5vPDyyxgbG1eByczMJI7RoyIakr744uJxvHH5DemuU/rnzq2bSKXjyA4P4MTSMZQKeUkH0aBu5e4yVlbXMTI+gcHhYXlUmCQlMD4yiuXV+xifINhhZBbJCd4X5tTcw3BfwljHuMtzoVSmOp66BvCNjo4JmKJB58TElOQnMkNZvPDiy86rj0BNC7FwF6dOHMW7n34H3rz4EuZmJpHb2UYbEcwfO4E/ee7PUaw2kB2dkOZ8uULwJ6lTJYDIeTuYyaiTlXsMyjkW83uYGBtBuVrEBz/4LGKRENq1BnY3tzQ2hWIBuf0cFk+dwvjwsIBPzUtqqNcrSKaTqFVK2N/ZUZ5wf3VTnRULiyewdPo0avQLZDxt1FUpeumVVzC/MK9cjIVrAynznWhRejccxcTsPK7fu4daq41QLIlwNKF94ubWtp4ZzqmhIVZhp8Qns7pbXSz0JmR3FT0CK1XL18BiLlY5A/t5SnsaYaddliuGYKdfqbCHTCKKdAw4s7iAqZGMznfl/jLmFhawvLqB+aOLGBgewc7OnvOZM5nakYkRSV6VqzX83cs5jHcO5YcPWEce/ejtjkC/kKF/pG+HbPDIiCsOcQezI307x3u71/WN/56yTx/N/SWi9EJsR0SmtppUYKD0TBSTU1MYnxjB4EACw5kkd2zYz5cQScRwf3ULq+sFtIgXCPiJoSpfioSeCa6TBr6bfDdxA+I1ZgxsubRGjNJp7SaOLx6ThB67uggsF4p5K4ZLJVCXh43lp8ROBgcyaDfb2N7YUrcC1wXGA8ZByjdT0sgAXZKMMo1UVb58KptNzM7NaJ29t7wib4fhkTF1p9Ebkc8813aC3ZY7dEyqjmQGJbtd7qJ9nMs/WRBondksLiTAT69QhnXr2LA1mIU1tlcmyM0EVIWdbQLNZb2P18trFBHh5A09Qc/cRt6OTsZZFfaUNndSrwtHFhy54Iy4nbKIinpLZcXojZUVDCQTTr7OinIpc858n8eWlyu9EJxyiTbqTradn0uwPZkacLJ3UHeJr3LjuPkcbXHxmLoqrrzxuvw42UHPe808SfLmql2gXDdNzSktSzPpEetU0ZoQkcwe1zGudYNDGQyPZFV4mYzH8PxnJnuT+50f2UaxVEW1Wpd/HyXDiH2Q9DYSgV0uhgUS9DeSiNLkltdzHVURmsu9lFdxj8D7S9at07XOOal5UDHG+W+6DkZJA/J62DnSbWNudhqJVAy7uzmRcvSSTcQSuv6RkSGMZAdx++5trU/sWuKYcN4ZJmqFmkaOk2AheW8eIx6/sS4h67AwJYeO5noqmXbF2ZabMmeU95P3RYtOv+s/zyj0jePUt/EO1znx2MP/dOOLwU6Lb2CmjffiX7/y6/jofTPG/nY9Kj7wm5/G5z+4i3908m/hVx52ar/6e2h+LIHfmfkJfOwB73lEVPQH5QQ16RwJYe1ZLQOvBUKSDjeAQuwxTXAD7dmykHYG3AZEmVEhgwWDqqSKXBUvW7KYFLKFr8sq+5YDu+JRaXXTYIndBWyzvXHrrpJlvrhRlEmQa+GwBYVyN9S2M4CUmzZtKsmGU0qHLb7tlroZ7Bh2Pdz4ctHyRAWNE7e3t8U489yZnPMB56LLY/NYMtmJsYvBuhVMHt0IEGmoC/yjOZC1xlNuyMAE60zhuauirVyWtJDtsm2T6xl4GuvwemhAzeoAC+ImZaSxlLkOdZWt5Z5jyLZDJtxatJksSI+1qnMUMVKpWidHKKTFi8FQ1Q6U3OkB1gYikhXmfaUGrRhbdDE5NSmd31CEm3XT7WMgJahNjeT8/r6Ox404F8DxiXERP7UGF31eom0ASFjQHUPayzRMioRx5Ph0r2rSb0ItxzMiygNbXBS8Aa7uO02DApXDBx5tQzR7eaK8N5hTuZ953eRequo6L+xkLSkwoMonn7ZwSyM3QFR4uSmdD0FIf0AHSHuQN7dfUHsmv+fGjYsNWzIF1nJjTx3wsM0Zk4YIEhWUd4iaTIs6YFL6mlV5maFRGSmxCoVjz99vb23h5ZdfRCW/qc2dJxlEnCWp6Ukyw5ILT1T4KmxPVAQBMF9BK58QJ0El7UpXDdknKgwIFODjEzmSWz2ZKSZkBC9s2nNec0xlGOXKUL/61RfUEs9KhLdNVLhkWBcqnwj/wJohqeQ03OthRAXvFxOFsbExERWsLqlUq2plHR4extDQsDbKnqgwoswO6j0q+kSF+n564x6cr8IrA8RcD9QjaeIr/y0b7BEKfpNsBG2frPBzzoCAgwsej+uJAhuQAHh5CIjuAf2HZZFchbaukdIHTvOTc4t/c5io0CdEwwIgRLU6QzZ/fD8PPUlhj76RST2SJEAu8md+vvZ+330rUeGvXJ0DDlA4DNTTr4BjoA1GoArfg3xKFD1R4RBsfaYu6q3pn67JdfRJ/khVZSZpQuknLqDhUBuZWBQj1LVePI4L584gHY9pg7ZdzmN1exf31rextZdHXtqx1MeuSxG11yWiuNT3faDMUBBkDI6tTQ3nfeLAZn+tRlQYKM2XJ8f4NeM4z5XHlYdQoOJc9yxAVATvmV2l3TvGCVXmd4xk8eMcnJWenAgSEzpGoNpa13OYqCBU1mo7f6MWOiTDHQHm54WfWyQq1Fnjuk9kOEjNda5lAuLtjPxaw5v49ogK26T7GRI8n29EVMjPxT1Lflz9eB0mi74loiIAjPsYYMC3rWnmS+RI8bDzE+GzJvC/36HUr+rijwk89DuTgufTadOLil0uVvml6q63RVTYRo7rvo2nMpdeB6/97JsjKvinJGt8NR0NJ5nP+pfllXb3uIZSa9s6bCy/azcN0CeQwvnD/E/zxRPjFk3MoYobYnVEcv207goB/Y7g8ffYd1PIaFQEP3M0/su1itWM1tWkIzt5J+aTfH57RIVu5EG5MXvWgcxgBu946glVPHLzTm1jVpYXCiXlarntXRFKBMWD3XWKhe55PtxVY2BTHWPjozh96pRdv+/W8xKLgYfdH7f3rAe6fHokhTsGP9Nfr48FB2KEiqS8j15gHSPkHg7j/ORZhMJJrN5fl5k2fQJopk0Jx5mpSayurqpz++TSkvLYublZrC3fx41r1zE2OoHJqWnsF4v4y5dfUkdFs96Q9NORo/PKtVkMcuzYUbx68TK6rQ6OHD2C+/fuYGQsi2ESFaeOoUBvhUQaoU4E6xub6qKoNprIZLO4deuOOjVJjgymB3D1+jWceeyMADjdxkgYudyejDwJBjF/N3PNDlZXVjA3Py/yNb/PDs8IJsYnzHy70cTgYFYStKmBAbzx5jWT3GWXPB+XZhVnTi7imXc9heuvX8T0xJjl76EwpuaO4nNf+DLaYUoxjaJBCd9G0+RIOl1sbW0r7rPDmpJOLDDLpLiHa2ByfBytdhXvec87Eed+qAOs3rotkJCyTxubGyIGTp85o2KdcqGEhfk5yUVJZjhCkNOkQGuNFq5cu4mJ6Rk8/sST6pYjUMUuv26zgdu3byM7PKz/1tZXsbOVw9TkJLa2ckimM5heOIJXr15DpdlGNJFCp8tn09YU5pZau7odGZYPZwextrain3FfwgIsmgBz/0f5rFKp6iqgw9ja3kV2eFRrDnN4KgSw4IrScZFwB6lICCOZBI7NTmF2fBihdhO3b97E0ulTuH1vBTPzRxBLpbGTy4uUoJn28FgWycE0cjs5hGMJDL10DT9bN0neR6//1CMQJC/+/wvv/YPCFXyhm0MqGsfwQAZD6UF0O2FsbebR6TBXj6NUqCCdimIgkRRhMbcwg6VzZ5EvVrC8sqE5vJ8voxuJYr9QQpcEPvd7zg+PMYuFkXzmvI8cAXutD46oJKg6OjKC0bER7O/v6xmYm5tTtT1BY+VmLEpU7DL552KhhGa9hUQ8LgyEeALXUnZWsAsvLeDWuoCJiwwMpAVaE3NZWjqhfTj3cOzG4FpMnIQSPCysZL7KfbxylTCLVctot7rCU7jP0fqjHMAIGV8Y5CWMCJQzbtPX1Ev2WKyxPY26tUjqKD521KFGjIx/r/27L7qURLkVL/j8wOddHAvuW5QDRKOS4bN9oZG/6higVwUr6unPEItid2tTHRXqAHBdesGiMJ0XC2SZ2xDED/N7KmlYHOK5UOFgfXNDig188bpIhpBI4tpkhuk1sNOOOIm65pkfNEi4V+VnwTWEqiXMWxaPzskvaWpqWuD+9es3MDd/RGseAfgzZ8/h7vJdxVoVM7abeP0rp3oB4ekPr6NcqavLTRJeKtAI6Xp5vuyMicVpqO26QBzJb/mQeb7ymjke/UJq6+bkPeaCIXxQPo/W8eD32Ybz2f5aMsehLsYnR1VUynksx9JwVGM1kEppjaEPE4kKdiA1VQxO4iZsBQecv8L33H1nJw4LjwP7GY/VWOG1nbvJRRmu2S/ANH8PkmHqHP+uIiq+7xO48Ycfwf5v/Qi+5x+svWX1eCvR8I2ICuCAv4Q7fu0Pfw6Pf/ylh6xOdsxnrhq5oZc8K57G3bd4ZPhDOIJl6Dl8+F2/iOcecORHREV/UKbFONpi7R+M4ObAV0NJq47Mr1qnaFzNijyTsRGLqaBJDVADKvmSPpx7EI1sp0l2DTECp5QASiZkQMRkdXxsRMxsOjOA8ckZ3Lp1VxsDsuZ+s2uLhOlgC7hiNThlk6hZmB0S08mHmRqGZIT5XlbgsO2bCSbZcnZccANowbChc1xdW9UixsWMRIl+V2so6beNk8TG5f9AYFbgkYKeGd2o4tNwCo2LtE8jYQVfjgUXPRIRJE5IWngDcg0SvSGqVYGWZN+5AWVgaoigsRY7tRPSqyAZx9TkuMaOGyeSD2R95WOQTPVaFCtlXgfb98wzhIsxNyaFvRwG0tRfNQKGQZXVYqwUI3PrTeY43vys1fVN7O2XZS5NuSxeA6+ZF8oFiwGfrencLHHjpMW420a1VlHVlLQfwRbRhiSg6GfBsZw5OqZL95V8GmO1NvqOCg1MryvCaYxZN41FaKtctC+dla3jFdyxFLBd3unnnp/1vc2/A5k7cBUCYuP1JLiFwAB2v9CJt/CSQqqItwTGa8KLhHD67ZI+EyNPXUPfNmmdRnoPuQq1fbLjhZWr1vHjOzl4P1gdNzw8ogoE6nGmBwYRTgwgFjdpJ5NM6CCf38effP5zKO0uq+WQHTDeo6IHJgdAIwNgLMkxUNeAYP/y4KUREjFV+/J9XkbIy0Bo4XV6j3ymOd4+WdHxwwZ6cqPIcVOrbRe2+WZ7arGAV155FZ02qwosMZKO9rfZUWFrtwO83yL9xAqJfgXtg4gKD/ZybElKiKhIpVCt0+S4ouRseHhUSfSLL76EtbV1V73qpFY8uB7Y73g18yCQbNO2qzHQPHUdBLofrhrWV8ny+yD4acC7I9McWeHnp37nmDP/V0auWgJmpEn/5B4EevrzPACQ8k8ClbqMjzyeT2ol/8UNidP41HHpASQJpX5FbZ9ocZWJgfsVXKb9eASfU191ZISC1zA/KPkTJDs88aAE1XUW6LlTm7F1BflrDYLKPi7xX7/G9O6JR7cDJ/sWooJx2RH8JCpC1KgNtTA+OIgzR47i8VOnMDEyJO34vfw+tgp7WNvZxXqugN1CEfsF+lNQ49UqkjyhQOBfvV4O/NeYO6+Rg/HM7rw2MC6e8Fr9HNHzJVDaKnSCRAW74SIR84Tgc6z250BV/oOICv/MCUB01XXqSBPJ0icq3HZV5+EB7ODz2hvvABF9mKhgfCFR4avDOg4UD11n1SUAACAASURBVBJcit6MaWZM0dOy5RkRDFblPs/1EKPnY+GDOyo8SO4WHPf8+XH1P1UC4F+eCHdPnOO/e2tWsKMiFDWpAz8nD4D/h7xAvlmiQoup88rhKRl4wEp1xnkaEfquCN8FywpBduFE0XZCXsG8S8+QZACd/JLrZrXl1uIKQXaSXZxXjPH87+0RFbY5p6dIL36yU8Z1V1icMNLJ//7rxTT+zq99rGDThtS9+n9vm1TzzTYPJQMrnI+KusVYCWmdEiLiPVivWOs6eb2coyMtPGHhY7fWRddpxjnH6lLmkb6jgmsVQRDXutwDJFgdzmN5osIuvn/9wWeK1YlPv/spAbGmp+07FVmw00a9wupEEhcF7OX21CnIfJlVn35j7mOnxR6TWm23axijX8DiopOpMhLItwhZHDaC2oYm8L0jz4L3ycdtdaT1OusMiOmNLQ9E/wtDgA7EJZEqkRDeOX8BkVASy/fX1D0i37pGFaz6XJibw63btwSenz57VlXtlDKtFku49MpFTE3OysS5UCnjxZdfEaDNjuTJiVGcPXdaMhSUCpqfW8Dli5dFRJ08eULV84lEFMMjAziyOKPOh0wqg2g8idV7K8gXSloa05kMdnJ7iowpFp4ghASLIJgnqzAByOVyJmsbsYIq5n4mbccq4YyKr1jAxXvG7k6CQZVSRfsfkiwbmzuSmbp5+45JanDtY4dUrYzHTp/AOy+cw9XLFzE/OyWAiWJ6IxPT+OPPfRHtcALj03Oo1p2JtDyQgEqNZq0mqzE8NIRIqINENCJ98lqZEhZ1fP9HPwBmo+X9IopOC31jc1NJEfPWpVNLyO/tqcPk7Dsu4Oqrr8rXY+nkccWi+EAaK/eW8dLF1yT9dPToMSuwIbAnEKirsZmZmxVQx/1Ko9bA8NCINPL3CiW0QmEsb2xim6a5CXbmEsiynJoSGfyX0l/jk+PWhd5qqeiLoOb29paed3Z7j49NYHRkAju7OXVBrK6ta59D3z/pwbdb0n5nJIxobe9gciSDqZEhjLMLKxJCbndHz+ebV2/j+KnjGJ2YQrMbwtDIKNY21rC9s4Uji0ckjVks19R188MbNfy1ziOyIpgHPvxrKzb5L+Hl5Xn/vzzX3y3cxT+PbGJ0cEDEWoI5YLuLgdQQtrYKqNa7+PAP/lXsbOewtrqCleV7Kroq17oIE6OOEJtIIRxLKmbQn7Miz5aEyWtKKtGBrPLZsQIFgtRUkmD1DmMac4PJiQlMTU3gypWrwmgGUhlkhgaFGzAmsXjHjJ3Nl43gbyY9iFKpouc4TuPgLgF1SmbHVJBJ7wjiUFwbua5bIZLlYieXTqo7+MbNWyJIFo4cwb6UNEgixBVL5V3gCnDpkUEZSpKWxJm452MMJlZE3Ijv5ZFJWnjFAnqwkvCU6bXvHkdIOBIxEebDktbusrMxr/eZCoaXHTYZKOYDHh/wWIKXX+YelF3qxIhomkz5br6ff2deCk3EVTTaUt63tbGGNrsNaGbNDnjibSp4dHJV4TDKlXLPC5W5vQqMnLQqz40yURzTndyOxsMrqPBY/ByOz/jYmPAkdnHQvJv7HRY1syBIPmfRKHZ2dpEdGsJHfuCvIB7u4N69e7h7dxnb2ztKUa3DJY7/6sd+DM996UvyfGCh4PT0BP7gN/s52plnrkjNhIWblOhjfLfOy763HeuhSXpx/LxHRb9rxCSdiAUa3sQuzhaaJGrcvpnn7e+NgUGWX1lBk31hvopdHF88ImLk/v1ljTEl1Tj3ed9npyawdHIR125cQyiWkqQij9FqdbWGkGQTflavy48lnUzq+fC4DM9d+KGTHaP0Y1+ZwKKJ+QJTupC5OWQIrr3QdxNR8Q07Ht5CZHwjosL8Lj663TfQ/vgffgG/9p4iPv0//Rx+/HcPkyHvxa995hP4+Pld/M7f+Al8rCc99TR+7/nfwE9Fn8PP/MQv4g/uHFwCjv3sb+DFX34CG7//cTz+PzyYAHlEVPTHbM4ZYvMB8W1tVilmhs6+golByVelMTDqAeGmtsNq/7gCgG0gzRDZg9AMCAyuWrwcxGYMsJkGDg2yaqiq6k0a07A9d2h4RKy3/xx1LJDh9gAZyQS1Q9HgqCogkWZMTGD5Pdni0ZFRBUJ+KKujPKBMCSpeK4HI5eX70pDN0qeDBIi8HsisW+WeNxLidSoACBR3xoQStTfSRkRFoBqYQYxbKi5wYs0JrpEppfFUzyhJcJYzh44ikYxLe5bVeFb16GQnnDG4gmbH2uGo+06DOgYuEi++88IHuXgs4XQSCcCbsR3vz1AmjcnxMdy/fx/nzp3G/eX72gxz3PkvdQ2PnziuFj52V3BMNrd2tXhxjFkFwHZ6Vpd7EIr3hAk8JQW4QFXqVcQTMW0Q2Q7p9bBJVGjzzQqm6ayx+E77XPPGV4k7SShfNS7YzeWkxJ60VfU63MGyWIPxdJ+9xII3uzKG3X6vCnjJGxnrIIglRLLO5q422G4em5k5/79vpt27zyIonJ65O0HhsxGSZzFJ3ihX4mdQ/zDKFse6xs727lbxzASQXRxMmhIJkhNDmJicwfj4hNrbaX5OgF9VmSQnWO3tKu5VG0tdxkYDf/5nX8LyzUvaKCUoOSESL6ZkQ2uwiMQ+oGHXasQKz8MbS3nQ1gAm6xxKpNIizDiHZD4uvxOTFyNFx/vIhEhJGg29VBVAgo5ANee8VXzSVIwdUhr1cEwSBexo8smGukucBrqqUwNa1D62SA3fVUx4ctRHM6vING1vw866B3TaWfXRB0L60kem1e41z00Ki/Hh9OnTmtvcrJNMJCmazY4qKXnppZext8dNNMkFm8GKm4fMQg8DvQ+t3+J4+wp/3ihVg9uVMR55jXN+f7hLwAgAb7BsiTGPRZBCYxHqaN4xvtv9cFW6QVD4EAh/GPDzevcexOZ58H7p/BzByM2/ycX126a9TJeAQGm1B0dAji5v2cP5OegNiIPgmxm694bGnl//0Doqxnc06P73EkynOOploVyHnR9PfWagy+oweSFiyWnKBkkn+9p1jThDbdcLTpMWGcQlog2cP34S73r8AhbGpwSSrG1vYHVzAzslGhQWUKrWVaVG4IIarNJTddKK/twCrKm6+rw8i1+vJY/kpSkCfjo9QkakJIkK63oIkjgGunPNMoNDznFWpPnxYVJvY++IwB5QbQm/f5+ID/lS2Gf171Q/9siDwN13/4z74/qNmuZ4SKuokzw0KT9WOZOo4MasRbDNVZUpcXcbFo2H87ES0EqSwpFovqMgOOn8+AiI7dq67ddp9wT2gfJ+v58VeDi/BotXHlDvr0HaNFMvl3JTbjRM/sn3iFIZIKwNcd8bxcmVHQJk/Tn37kHgOfCG5/1K9KAfgAfFbQ2wOdKjP637RqBe1KqMmc+4tcKIbPef38wefmLtAXCEvG22eB+Zi/lxDD4z/HNPjBvRp0W711HTW5dcd6V1QR0E4+359KZW/i7ZbLM8zRncB//OtdVzbrPLkTEteF7BtcEO73aoLu/rSQ/ReJfrddI0rgUyuFzCvI4szolQcH4VIhYilO6xa+nPd+t0ZYcx1w51ngrssHzJXbiedebDJjFqnWzymuDYBEixngcKQkgPJPH4k2exQIBXppjcKPPRjKMlDTzmhzShbKPVYJUN898a8oUt3Lt7S10XzB1ZRMDuELtXXOOaIj+O0WvBrdG2Xth6w/9ZF51bZxxZ7vNav6fw8czGol9o4r/vS7Ax9a07osyeHS9lqrF0xSLvXnyaqxLu319DPl9S8U6pXMDp06dU/U9/CoJUTz39lGR/SNQ0qjW89uplAdQzc3PIFfJ46eIleVE0a3WMjA7h+PGjAl6KxQIWFo7ghef/UuOxdPIEVleWEY2GMDo2hFNnFyX9FOmG0Wp0cfPmbRELU7NzKnDK7eUFmg0ODCpHu7N8D+NTk7qvg4PWzcx7oZw6xRw+gbW1NUmGMh+knBJjLd/DPdP4+Li6pZn/UQ6C68f03DxefPmivBlUaMIuiGoJ50+fxDvOn8Lrl17C8SNzuhaa4Y5OzuJP/+xraHQjyIyMoUEfE+UcYXUAROMEwXissI5Ff4oku761rkUQTYTwnu99NyLMLdpdbK2tY/X+Co4tHkUkmcSNa1dx8uRJxZC97R3MTE+hVCjIPJUEjwxUR4Yl0XT12g2cOvOYZKwqxZKO35QUVgrXrl3TefF8SIAOZ7MoFSuoVJlTd3D05Clcv7uMrb19DGRHRBhy3lq3UEdjyA7vwaFBxKImk8vCNc7Z4eEhVEpFxQ49p6EYxugrEkugVK4oz+Peh9fAIgJWdsdZQFYtIx4CBmJhRNHE3OSYZI3z+3vyFKF3RjSVEkFxf22DSbPixcKxOSQH0iIGEYni8uU3sF8q4b/tDuKHuuZn+K29gsD9fzkg/rd2jQdW7N5a6juWv/1jfSt/2e+e7u1JH0qY9H0x/tOe48HrIUnxib0rODo/i9GBBMYyKYxRAi2WQDSSxtWrd9GkTGdsAKlkxsjRJnX+w+qsrDTr2M0VsLqZ1z6IcYAdYtVmS+C15C4Zv91SzHWQhY0k8rlPpSIC38ecSsV3mQGsrtwXzuPjPHMFSn/T86ZULEp6ulqzIhkWCrA7Cq5oJx6jj0OlV8FuEyEi/IjrKD+Xay8JAskCOVUBgdaplLx38oW8yUZRXo5SRVTacKA/YwsvxsvbqghXxblWeKPl23X2+WIu6wqr9kgBxgniJCRehIN1rJqf+y92MDInUBwnfuM6aZXTqsuCMkbWLc71U0QH/1a4SFg5x+zcnM6bxQ2Wg7KQoq39Prvz+HVue1vdJ9lBw1r4Pq4rljexYyShzjBhXPR/dfLlvjCWRayUXFehpeS+rePapKpNVpYFmMK1SF+RKAoBo8NZ3WMSEwTOuUck/scxT8fCmBgbUoFsPl9UcUSxROyOqg8xnDx9Gm9cuaK4ODI2jg9/5EP45b/7ek+V4ML7b6i7h53mLLpgZ6lwO0q7O9l6xKwQTcFc8vTcy9g4ea8l3hN1wrj9iWF6vB8d7S96ubnLSXp5N7flylVJcDRw8sQxTkvcW74vySuuAoMDA5I/zwykcfTIHC6/dhmVJjMiU5+gGonoDxWLWdEd70OjVhPhozXG+Zx4yW7eN44754cKDiVFaDghnx1+zbnA+6/iuu8eouJBJtqHA7rrXEh/Dh9+76/gOTycqHjyw38T//3f/2n81BnguQO+Ee/FJ7/wCfydxxK4+8Jn8dv/6iX5TgwvfQA/+19/AGcSaw8mMT78S3jtN38YZ+p38el/+W/w6RtFALN45kd+ED/1/mPAtU/hZ77/f8N/fMga9Iio6A/MNGWeAjrWvkpQmwnfpu2wJOuUMHkHmSNFoj3TbT5ABDHlfaDqXWPW0wNp56VgFdv8LLLTBP30sFGfrV5RuzPBB1bpclPGYM7qJyapmcFB6y5w1eqSaGJlFyv3yKg36sjt7YuZ9O8h2MiqdmkmNuwhZlCmKRsXL7WuscqmWFILIIMWq394DWzlYpLKRYGmQmQ/eT2qfFKlvte8t24Fv0kzcN1AKwV3t9HkYq1xdQXNXLAIDFDmiVU8BJPJTFcr1pJPE24jMQz45hixQqDTaihB5qHqdbaNdSVNw+4GVhhIXojash0yrfZ1dihrVUXU826SHKJJOisRyqbl2Olo3Pg926wnxscEUPF8eN081k4uJ7kbkigVZ7YdZlV/JGbkRdr0YimLwHtCYLVaK6s6l4BIo0mSwzberJxID5m5sxZkVzVnm2Dz7wiC5UHAkH+rbgpfSR4oqnHYT29i+79TMiRSxAAE/5+Iit4u1wDc4Gf1/r7toE63wPt2QCO+qIvmwA6nn8w5wuQjlYyr6oo3UdBxNKIq6SrvQdOAOsk5xdNIpTIYHRvH+PgkRifGkUpnnYSZAUc9EInATcxJY0lmxPQweQ/eePN1XHzhTxHptpESUWFdFdQ/VyohWRer9gxepzfL5HE8aOMJLy3usZh1Fh2qhDZdZdP85/tYzaHkqmmm97yvVtSiJ0fPl2TCmtYJ1eqE8MXnvuxaMJ2ep5eNIbHhhMmDlf12fmau6+dOcJ8gosITWdKCNtPaHgDlpJ/89x5Ql4E5OwAciMcxymazMtNmnKhUaW5sRoo0zGKr6quvXraqRdfBc3jsfEwNnr//WXBuHth+eRCf10k5tsAvg4BasJI7CLIq6QTbpWm6znlnup2Mp/VW3SX+B0lV5fmHvDI8kBY8Nz+Onqjg2HmiQrJfruPGe2L0AHPn/xI8z17i16Ou+5/k38dr990ovfcH9NSD53ZQfsU6SPx9kQRYYA4E5baC5+TB2OB4BAkXno/I1UO+Dy6IGEhH2ScHwtLMmUBouNvC9FgS73/PMzh37CSS4ShyuX3cWSWosoO9al0bhXKtjr39vFqbS9WagCaTweuDqZ48MiCJHjFGNvDcgx0nwWt4C3FB/dWQrYX8Wx8PbE5ZVby13vfle3zRwWGiM3hfPElgFdjsMjT9XsYuX3UefEYO/62fc/46RBpwBjiPCsHZ7NiqWTePiIoGfTT6RuIHiApJXBGAN68jyVZ6MDzgVePPw4+TkTX2jDzoOevPO9eR4OKU+TswrhvI52uwVH3FvIVroadtvCydexeLEuRT4Ym/Q9Jr9plufRROa2S9qsAcKeh9m0TIKD8hwcMcxKKIr9jz86Wf8jmDdHX0sVI/gibzFt/Z5QhGjaMnKgLcon9G+C83rt6EXfOHREWw2u0QGdpb53l+3CwHukeCzyOrNg/HqF4O4IFqFyxF9jqiotfF4q6F58i8k/OHILQnWIOxpEcCBc/VF6gYRq67po5FgTHmgeJBl5Dr/uh1PznpJxWsRBM9Pwn/LPt4eZCoIKlswAuv0553W4uZBx8gKrzXkbsIH+uYcxrPWcOJE4s4e/oMBjPDyi0rjY6kPrrgBt7Ny24C7WYU3RA7Yvewu72m+0HgppAvC2AhAEX5qEatjJGRYRw5cqQHqvTXVOvY8c+zX/96BJqfy66gpE9weA6nL2Ole06SnrGABQABgCjYAcopzvc8dewpoBPD3bv3USiUtfcoFPdx9uxZTE6MC/QvlNh9MCmpUubxJCquvnFFko4EgLZ2d3HxtdcwMzUtw/XZ2SkcOTpHZg2lUhHTMzO4+OIlxbczZ07j7u1byAymMDo+hGPHZ1EuWkcFpcKuXrmuzuhMdlhmmrfu3FWeNEIpjEgMKxsbmJmftWKHcBjsQuCeyiRJogK7d3dpIJvG1uaWzLX5Utd4Po9TJ5fsmgpFjI1Polqrq3r/5YuXVFxCgINFTa1aBU+cXcI7zp/G6xdfwPEj8yIqQpEY0kNjeO4rLyCcSiOWzEj7WxIaLDwJhQToVWrm5xKn/AgLUMJ04Oiq22Qnt4n3f+B7tadqVutYvnlbprbbO9s4d+EJeRAydhT29i3/BM2qy+h2WgKomo0aMqMjqqqtMZ3uUN97HLtbW5J2yu/siOBj5TPzMAJpHJ/pyWmRCMViWc/V5MJR/PnX/lKdFaEY9ffbAkgJerEjmONarVQkL5wZoPY6r5GxgIRJHOC6x5wpzKpk7mGo3c8cJyEpLM1TPxdVtNZBiyQKq1nbTTTKeXWtsEBpY3UNg0ND2ON9mZzG5OwcXrl0GZOzs9jP72NoZFC/ZyUvs7Rbt+9hdz+PRDqBMys7+NvJCUwRcXv0+oYj0Ct4eChh8A0P8W2+oU9E2IrQJ/7/c+j2WG1V8ev7N/DvKxvqpjt1/BjG0zGMpBPIptPq3IpH0/Kf6IZTaNKXJTaAQr4gEq/VqiM7MoyRiXGUKzVsbudQrLBgq6lCmjrjcci67HntLG5QZ76TPeUz16ib9BD/Y0cBu5cIynJ8CBSru5EyijLeruHxc2ext7OLne1tpyxRQygWR4gxsdGiJqPyPi7CPF6oyy4NrpGmriDpJ76HpKlf19gZEE/0iEbGUq4d5ZrJZOv9ga5h5UosLHQmxnzuRVLKKJuyQVF9JgHtOOUhieOw48T5PPJ3zDH4XgL9ZhpuRQbMCRjHjJQ3HwpeB1++QMd3G3O9FNHMrnR+tmTXu/rMuVkSFTwPgtRRK46TvjJMRhDAfi6HYiGPTDpjJuWppH5PsohjzxhXb9RM8khqB4ZjMQdkfJWkeNfJNDuShJ0AvB7GRRXhcs8gvKZruJS8U0lM0Y+igQFiUq2OYuLwyBDilO5uEzekhHgcM9Mzkme8cf2GiCnifNVGQx59zDVPLJ3Eb/2fVOGw1+PP3hIxXW+0EJXHCLurm4rzzJ05t6IJYlKmaqKuGCd7zd/1ZGmlMEC59aTGVttFkgD87GrNCp56/rCuYMXnV07imf6rJ04cE2HBNTiVoBw7Se6QFGNGhocwMz2BG7duoNwgVsl7SGn6pPOiNbl6EmgkgLhGkuwghscXfyfSzBW1yFOkZd0aHD91MDnJKnro8vqE0Qk7+G7xqJBZ9iye+/m/ih/+1NeJ485U+z/+5I/gx79sRMUHhh78/lruLj79v/8Kfua3rh16wyx+6lf/Hv7HH30aZ0ad9la9iKsvPYd/+j//Q/yzVx/y+Rd+FL/3v/43+OiZMQzbs45aYRdXP//b+Ns//ylc+jqn/Yio6A/OvNuEBQE1Egw9s1FukFRFbaCybfj7YLEYVW4A2fbW7ahiiJsZPjys9CGzyBeDK9/XbLQEzLNSi5X7kiIiM89gl2C1TFUBXp0YsRgee+y83ssHlR0H9JUg88nWbAYh6s6SXGAr4tzsrABFXgv/xneEeACAP2PCyiB8YvG4zHB3c7s6Vm5vTwwwZXW4IdSGvWFmSwTfyfjK7K/XshfuacpZomK7WAFarFDrUlPRafxLkqWLBk3CaTArrUOabTdRp2lqh5uPOliHygVeqg1O95zvEUjADTA60jYfHRnCkaNHcenipZ53BxdB6rfyBEjK2D2DEnVVMgwMiDBgpbhtYKJo1GsYpJ5js6lxZ/USQX2aTnERotwUz4SbrHyxhDv37kvOhRtzJi/RqCXxAjjYjdJsoVQpqRqsDXqdkLFn9Rsr90jeGFGRSJF8OSi7wOHTptxVMnriIliRy2NYZ4S911cnaoLJtdmqOw6CxvY2MxY1TW67V75LgkfzHhV9BKYH5vf+rl8J6X9HoqgH3jnTKL6L88c8XroIMekxW3BUGzWZkamDQUBkBKNjU5IdWDh6VFUOIc2PAc13fi9wyAH9Gh8B6tTttoEgKCUyaWcTX/jcv0W3WUeSVZwRmq2TCInLHJUahjwHDwD5cbLF2ypcBew5Y00/hrwWdnUwAfXv4fB5ooKfz80jiRGBZAScHFFhI90nKjjnuYHkvVpb38Hl114/cK/sXFy3i+tisaqavsSPERVWwREEtuwZdNIQ8sUwsFomz72qe4tVfPm/tYSUoKbNEz8GmUwGx48f1/PCykKZbImITWN1dQ03bty045DEdABbD3jzJmwPqIj249qbXy4UB+etZdB9ouIwyB8klv1zY0ArJcWikr1h8m8cQVsxxmvJmuycq4IKdFY86HyCS6jjG3qyQEGiot2kZJDJ8b0doiIIRjIO+Er94Hloc3PIW8PfU/8+7yNjxqWWiGs+cF4ckBexOGLgel93PzgW/uf+fPzz49+j++alb5zylrpP2h1kqPWbiOGZpx7HmeMn9D2J8a2dbWzu7qharc4K2mZTxpo7u3solquKrQ1H/ngC1d8zVe73iAqLBZ6ct/HTjOg9V9+IqOgD12YoL3BUy5UZy3Gt6M+3gxXofrx5jGD80JrZsqpzVaG53MHf3yDIGCQN/X307xNdH7aCCV4WnzUCzKbtT11/VqFZ7PbH6cU3dgeIqKAkHfOOZq8j0hPe/vwF+rv7b2TNN0dU6N6ThhaYTMDarwdGVFi1muukiBrRottziKjgys44K0+pwLX4mGDn2V+bemC6Y+ftfV6qyGv4c+P6VqKCR7IxsrnP+2MYnMl0UfqJuYtfWw0sdoSPupAifV8mCz494oSbd14vz8WKJexeBeeJ//oAaeskvWzc7UoZp0xqigRgfz4H50ivO8GblDvRxm+KqOC89jJ5gS4HG/+DqcWD4o3mFivKpXFtq5wRpJ7wt2DgCXqOqwiGQ4UCDyYqKOnZJyp0XG6A4/ScSiEaoa+VRsnGP9BY4g2yY+rk4ImxW7mGTHpARtBHj51AenAEtRZBB+uikrxcN4V2M4J6s4ZrNy+jWS8653fGTuuoYYU6/6MppjqvHDmtggVHDtvc7Od2vuDJT1/e4/588HyyyxP8uKvax0oi+92ETnYhcOz+cawj6H2PvQ9oR3Hn7n1JLhGUopTI+fOPqQL/+o1rGi+akRKwbjVaqBSLWLl3X6TA9OwsNra28Ma1a9qvtBstZLMZTM9MCLzb281Jcun2zbvotrqSNLp29Q0BM2NjQzhz/oQkN8aGWVlPAPquDKLZIR6OxbC9s4u93T2cOXVKkk2bO9uSapJmebOpruRUKikpLo7j2XPncPvWbY0BgbzJyUk0aPwKqDCIQH6pyKKiCYH4uf19DI2O42svvKRj1kk4cL1sVPH46ZN454WzuHr5ZSzMTmNjfR3pzCCy49P4wpe/inR2HMnBLOiXVy6VkEinFf939nKqNqZM79z0JLbX1xAPhzE7OSYD7WKlgA/94AeteKvZxr2bt1GrViTVtHhqCdOzMygXCsoPG9UqMsPDyG9uiaSoVUtIp9y+sdnG9TvLqNebePq934tYN4Q6Pd66kKnrxuqqOuDTgwOSkYlF49jL5bG7u49qo4Wn3vNe3Lx3H1v7+1KwpwZ9ZnBIck98ZtitQplaEmySKHFrHf0Ha9UyQp0WZmam1ZlCKRkWE2kf1u5I9lPzn095yIiidDIlsJJCeSRumpUCzi2dQK1cFCEyP7+AW3fZMTMtM/W1zW2sbWxpD3T63CmMToyJTCMA+drlKyhWaxgYzODOvVsYGR/GM8U2kfzvfgAAIABJREFUngml8Fgsg8kQi54evR6NwMNHgGD7RruGy408vljZwb8prtk66orInjy3hMFoB9lUHKNDWQxJSi6MN67cRK0VQnZ0Cs0OFDMpEz2QomE1UGu2NE9rzY7IAppotzshVDn3md85yWdiPXy/wFOC+9rnhZCMJXXS/Pn46Ch2drcNf5DfpXXwsaivWijhe9/9buxsbuLuzTuodULIpOPIVxqIpRIosao8mXbkIqvebY3Q/5wMNNcmHpNAtUnmtR2Ybusz95cE4b1sEnMM5jxSEnHrsicOCPzansHkmfjMMy5wr2i+ktZ14X9PDx92aPnuLVb6+45BgunKsVxnqoq91AFiHbhWGGPnp891+zJ+b7gaMRQrzGVXCD09SFRw32n5L2VerUqK6wjJHHp/MA5zH+vPUx2u/JsOQfyEOsNMwpy4FL07KnacEAkVSoOzA9Q6Qfg+Xod8WF3XR5e5nqoHOgh1WTgLDKRYRMyvbf3mukySZHdnV6Q5iQzGdEoZcs0dGR1TXKaPCK+RBMR+sYBEMi2ZrEvPn+xN+vd8ZEdFk5zrlGgnOUZ5JBL1JIBIcDBQEv9SMZPHIUIhFdOSnOC1c87QT0WeHspPrePFlE9YYGm5tiSgfNodKFyhpG+708DJpePKrba2t9CoWRdFkhhOt4MJGbcP4srVq2hGWBRinrYkwKWqQYlQGrI7fFUFra47ifeBc8WbaZs3Cv2UWia5FSGpxG4K85zlPeNazb/hnuu7h6h4tCJ814zAeC0o2WRApWmAWzW9f4lldqCO6apRQsmqVviw2MMUErDHIMFAyEWByTXbplkxw+oU6VxzszB/VFVBr712GYlkTK1PrAKkbJOPDSIWolFtDtgO/Oabr0vvfmR0VMGclet8cJlIM9Dx3Pk9AXuyo0z4rT3KKry5CKtKrFrF5PgE9vf3TBqn21WQtuO1VVFEFl6AM6uBCkUiszo+NxIE8GUoK8DffCTUfaJE1qo3KXEUT7JKjcHculCYrPuAw2MRoDI5kaiS5aiMpMJKXqV1HPVVNQz4BF1tYRgZzuL9zz6DVGYI//ZTn0EoRPM6Lhimz5iIJXqbWi02Csg0mWO7c1mJOkHsTDrljJBbApcTJHzKJW1gWWU0PpLF3s6Wrm+Imr3VGvbyBezus22cRlpdd1/duLWaSGUG5FERkkB7R0kIx6JSo0kVu1OaGMrafTgMYAjwcUTFgx5AwhZa/hwAbKZVDtnwf+tIDH98D8rY5tlqWlVl6ogKbfhdpb2+Piz/Evyd+2xPlBg85aR0lIgYiKg5x1oRtlMSPOYCU2ugWKkgNZBCNjtsi2utjvn5Y5iZmcfiiRNqCwwzgYuntdEysy2CQwa66fwknu1JHRsvzu1KtYTP/vH/hVoxL6KCQIWSiljMzI4l0eQIHncdnINmks0Fz6QCVL3ogTu2c8bjSgoIdPsqD/6+11HhqlJYwSkSU4unST+Z9JYRRL662qoxOnj54uuqIA/q1WuRFWliwJwHg333jeFi/Y4KPw/8XBHcwQpsLwX0EOknvl/dH72qFYKNBCv7BrKMFdTgplYmiQpWOmi8ogncuXMHa2sb1qEQICp43CCJECRZDADrSyJ5gDg4z3vAJAeB5SkB4i0Iph9+bmxcHJjnDOgIDyejEfn+UDJie3cbDQ6sqzT38hlBYPvwufQ+x4TwejIfwaoPvqdFENidq5mU9QFtScwEKqIPjM+hjoogeElQ4EFEhX/PYXLiwLnbYBtRJZ+IQMVzpL8x8ICa30D4YwTB/d7ccmCkf69/Tmym6gPdFy4mNJsYSqXw5LnzePrxs5LhYkK+n99DntXJ7Sa60YjroqiiTOmnfAGFYkXdFXxivdGel2k6cM3OH8p8LA4arvM511P3QPknxhKrBA+Ot3VW8O+sMo4vruO+qseexYAef8D83H++wFsdx7x+BHw7+areHNWmtR/7/TN8kIx0n8WrCBAVkharmWSkQO2Wfd3LUQLST11KeLjzoeaNpCn9PDjUUXFwvhpZw599vY4K76Nj64i1dXd6ps823zyBpLjAtMcvVY5g0HkzX2DnZDQqouIwifigdbBHVCiQ9e+JkQ5BoqKfw3kS0WKUzS2LKSbP1ScqDko/BeeQ5gsRPs0Pqyjl71XAQrkiJwWgn3mfE7Wq24Y/SAD6r3V811ERjOdGMjmqOyD9FIyj3wpR4cfRqh0bilkkX/31+eMG54I/78OEeC8ucmNI6QgB/s7o2QHxBv7bmq11XMQBiQr/jPjNsK2Xh6WfZKotHxqOrxFRXKu5FpOosPEkacQcwMmRunHk75hrUiYj2q1yi2zdUszx0hnMLBzD/NFFgQUkM0wLfBCsD3rjzTdw49ZrmJoZUf6mORIySQEZo2qTzqpYwsFQ7t0jgV3Rkyfu/frnO7Et1WopLlvXz8F40o+pjlx2xYwqxvDPmYu1vlOI30YQldTl9z35foTCCaytbGB/v6iin0IpjwtPPKFO4avXrqJcqYhgYDFNq96UyfPq8n1ksyOYmp7G6sYGrt28iampKXVvZTJpLCzMyCBzc3MTp0+dwauvXEIinsLs7DRWlpfR6TZxbHEOx84ew/7GGrKZYZQLFSOeS2VEWHASjWIvX9R9SVI6KBrH5u4u4qm0OjW4Z6FJNjusF+YXNEdt79KSJvmlS5SjmtTYUbKEwPXC/Dzye/tosmo1ToCnhDF2VFx6VSCicj/6+NSrOHfyGN79zvO4e/1NzE2OCwQCjXVnFvD5P/kyOpEEIFCRIE4dQ9xDtdpYWV0VgM5nkeAlfSkG4hHMTU1he2MVqcEU3vfBZxHudFEvlbG9saFz39/bw2B2CMeXljR3WbbTqNYF7q8ur6BaqWF6Oguw4/DYEXXivvDCy2h1gMfOnVf+mozFUWChVTIt81XuXSIxK1TIDg0LTGNvR6XRRCcSw41791HvdpHOUM/b8kzbQ1oBDPdCJkNsBXQsDuP3iVhEnciMnYOZIREb+4UCcrt7iDhTXQKrAoVIbLAbi4VZJGZrFQwPpKS9/tipJUmUEejl3o3FB2OTU+pcKdcaSKczWN9cR3Y4g7GJCdMpT6Rw7fpt1ZVXahXpsycH4sjt72jfxHyWEjI8Vz4fUi5Q3LZ9JkFEnq/PTwlkUk5VTzzBLwKrPdNemu1ax6SeRa1RBvb6IiFPMPP54h7e7595HL93tUID21NarmRtbV6G0QqJ/h/23vNJ0vS68rvpXVWWt22qq33PTI8fAAQBLo3EoCSuFCETG9JH/VeK2AhFyERIsSF9kMglCS6BJSAAA4zvae+rXXlfWemzFL9znyfzrZoGBK5WH0hNIQbdXVWZ+b7P+5h7zzn3XM8jdK4LBPTPS8ZL4QTxFc1eLOzBn0MyzuM+AOPYuyEMsWmlTyPPhDxVYG+vp/mA5RtiQPU7DKIO7c3qmReQBV2Gxxj9C/I0JXF94XqDHs7FKH5eyIZXAD0Vow7kShEfLXuUb4VKRfVzxGWCfU9l+Lazs6f9gIHj+wC53C9r3/tvRmvlQfW7zm8p5x1jkJq9H+Y6+OrWqgD1DoBLzX/UtUqxYB+8/YZNVQpWyqYsn8q45VA6b198dceylSErlEesFV7XUrWBK9I9NslbowVhh2MCsQ6Wg1nFhqxJnjvXxrNAdS9hCu8FltFsac4inBseGlIPJFeLHwqYTad7lib/bNTtw7evW7N2aGvLK7KLA9T99OtbtltvWrE6bFvgMGr+3BNRKTtynnF3UPWAuIH9S0JB+ndisyRRpNvl6Fg2eini7e+iVeY6c4P5zJx3sZ6PKfOG32FueTPjngvyAmEup44wb7h/z/85070akTnP/kUszHPl2j3n9fnhcS/r0O3Skz/T2ozNllXBQoUb5858v9raz1rAdb8x5mO9VhMxwD4V5yxrQtUXoTE40whwn7nMlxcBO4FBzs+1YoOOaJjcHzwMgF19WqNtlQj2lnrM5hg/+irRp4feFKmU8D++vIdGV2uGMSnSq5LKPcXyPRufGNc4jE1MWb5YFKFPtRyxzif/dj6GW/bG91+oEfVebV8YHWeBW1UhxHPHCARSJWGTWE87CR6xhNjs3MVe/vNYTBOtYcH0iA193AI9HMRf7A+xYhei4vKVC7a3u2P79FVptq0gTK2s15+am7Hx8RF78eqlHbSOZLVJDEhvMGy8mJJcIzE/FRX7u7taP1EoyvejdaoLszyWF44XnhlOEN5Pw+cQRJL2uf/fVFT0p8a3f/mnPgJzAg4DUBn8ANwr2b+PtyeLRrZCRUqs6MnQc9IhTVPBvEqOsGhi06BEnMOJzb1WO/CNvuCld2wKbCLeFMnZ2s2NdY8PQhMeVECUUXGAE6Bx4JBgwb7yeSh1aIYDcDY2PiabJjYqVT2kvTkxhwGN8GKjaQ8IABopl2srcKDUDCAVgID70cEOsJvJekAMPdwHtkFdPPBis1UCHZhZ+QhS9hfGkQMvMrcCA9KA/kUFWtyTyrwDe8+Y0AyKoKUtpZQ6N7onY1CWM94eCBIUHlmpkLV33r1u584tWKvVtdW1DZEsbPwvnj0XWHBIGTUKcJLifEHldeqBUCrrGXY7gDYccF5OTwCvc6rbtZUXLwQAXcP2pkwvEhplp20PoqlYtDRNyrsmz9VW+0hJEoEMbDhxWBMAjvtIHckfmL2+223Ja5xDDaKiMgw55CurTyDEGHIgHE0c5AFQEGDqgVpU6cb16STHIJg8DnwpTfegJjTHBKxzUIJGVqHRsCN1fcIhCc4dLzH2QN8bog4uWNcgNAzfcbf/qhSL1mug5j0SKFkoldRMjEZWKADGxqft9KkFO3XmjJIvyltzubKeF3PZyQoCYicR+uBtALLJAAiUW+2G/fqXf2tPHtyzcr5geSk4cwJGICrwF5ZqIKxx7j2qI9S0U8oRylQHIBv3A9nGtUSiIqopBPDI97qrZI8EXI3GQh+WaP0U1SLyM/XuuLJO+vLGXWs0PSDQHFDwHf05g2d1eLhJgEuGQIE8Ork3O6ARPJYDMUAC3f9KvC7ueUo2tLbdhzkq9tnzsLYAJCDh7Jfkds1u3bpl9boHgV408s2+D35fnqidJFT6pELSXiWh2HDCRXKofnIXiYoYeMYAMEmGaA8jcbQj2X9dvnDevvvd79jW9qb97Of/l71a27C2Gtu5DV0Mtn+XMw7iI34WARRf7CX6XihLjj+PSiFfDwNLsSQw7j/zstskWBivpT8G4RvxPV9HIug+Eu/zDeun+JyCnVTcG05aRkVwOZIRA4CV5Mz3nSSZ13+O/rA9iuUcQj/T69rC3CmpxIoE7VjrtZpSrHJWtegt06GS4lD9mCAxUd/u7tWkroyVX0nCIbkOBPUHz9xIBrgv/iC4PgYGJ4gs9j6dQYHRGIDRvk9GooL759z3poCeaGm30xxLAA8JQs0/n587gC+iNWEtGefvyTUhIDRhE6THnnK/e+3JKFlpaCjFmNsqekXFwMosgsxKyNTM2KtByQp4XbSypHdS8it5Vvi9D86RJMjeJ4sDSCzAJvQaUo+C0MAxbGrHPoPc/hhREaML+SPTDDgtIcXASjJsL/GgDO+WJKvUXDzcf5y7x0gMRi9UwsXk0p/FoALD93wHOPR3lFs0Iwy+/yIjgtpMdmH0KFDlyKDKgc+Q3Sc2V4m7jhU58dqSA5IcSwHd/R4Vvlh5f/WzIdaKANIJi7q4NnStYZt/nfVT/NwI3qjqFsvT1xAVPr2PV529bg/XVYYqFpJnlKWyoQi2R4od1Zsp9GrB/oGGpKF/W/IzRLwlelRIOdfFlikKEljqLiogHkgSFTojwhmq+R3AJoCLcjFrhaOGZSEcpCDvWQevacNDu6qzbWpqQsBuLjti6+uH9vGvf2kbWy/tw++9K1DWLVfdRpVknHine0RlrK8hiQgi6Bf3gRA3y2KDPgBhX2JpoUv3vD/Qu2F+D84x32djRSQ5BY1UAYwloApkaSTJtI/1vJHq9dNvWS5ftKWlF7KpAuiiCvu9995RHvP40UPlBAtnz8oPmniD5qt3bt+1U2dO2+johD178dKePluSwGp/d0fVFAsLZyTeobrhvXfes3t3HwgoGx0dsZtf37B6/cCuXrtg73z4lu1urMkXfHd731ZX15RnjNBzL4h8AGewmGI8N7dcKCW7EKy4jo5sd29P/efIo4g/6LNHXz1yLCo3UAxLFYuvO5Ym7a5eg3UVKmf6INy8fUfNvN0Co2OpTtsunp2zP/7+B/b0wR2bm5my9bV1WSQNT8zY3/7bn1uuNGSZQllnCmKkkbER7VBr2LDIfjStWBaLpHSvZecXTtvh/o51Uz374R/+QDFAt960+3fuWK5QsEvXrtnq8isBy8PyvW9LrOPsFp7cNMGt2c7Wpi0sntNYPHj4TJUub775pvYjQCOAR6wu7t29L+BNgpo0PfqGbW1t3Y5CFen47Jw9fv7S9g6bVh2fUD7C2pPCG7TVN2X3TM+yNop2WK/p7+RYVHfQbBfQn73oALub1Q01QYdsAkQij7l88bw9f/FM1ePkod1m04awyqkf2vTEuFUr3lCVfWtrd8/GpqZERr1aXtGUJ9Y+e3Ze1k8IlbK5kn11846sUMmjVtZWbGx8xDa31qzV8Uap5JyQWarOU2NzB/IV73YBu7zfBfsQcfbz5y+UiwNYE6MBartimFxnAHa74jklhTnnCHMSQBJyhy+IPgHs2udcYOie6jxHgEm3f/H9x5F+jyk9L+qf5yISQp/AQExHqjvmM76Xu4UlMZQsNvte/T3NI9YgDgC4MDTpD0L1eQ4xBGdUxnZ2921tfUvXzb0P5NCRdEhUn7rEzMnzRCzcz39Uod8/dGOg3xcfeM9OB7/VWLmQF/GrJvBULQcCR9ZH9ERqt61Wq0vgKKIig7++E/xeMeeArkB9Ka1d/KjYhPEP1pKc0Vywev2p6tYb6WoPDoSNCGz6KKlEtmvFfNauX71ghV7HRitlG6/imJC1ysi43fj6llm+qIqF8vCwxDQVBIyIj6jkwvq6Z9Zo9kS4kvN3uk5Qg+uo4jbYsUUSwONGV98T20rB3mrZ6NiYXDTi6yCcqBwsZHqWbjXs3auLtnhqTk4UVBY3OmbrezV7/HzVnq9siMjiBOHZykY45nbB+onoRPagbao9oOddrMSUlI8/ZBKVmpxhUINhDXG9anatQnYn3rTnBVGD3C9aLtpxpxHPWXmNz9dQZVWm3yQVJx2tReXAod8pVtz8J0shCJRoUcWjx/anWBQxEC3UlaMB8tN3okPsyhVj9V22+dOnREKTT/Acyb2Jb8GgCrm8qu3WVhDSOa7FXOHLMS2v/OR93WLQe3pofaot3JEd1uq+b1CZEHpgqicFsQXvE2yR8sKxcFHoyAqQey0VQo8QWYUiXmT+hngqYIpU+bGHgTthryirVAl2iIXpp9iTQ0omV7Tnt673w8bpK18pNlXTchqYc77pWTkBQ1VLzEtUJQKJxD1LWImln4+D7LI5c8Eg5RLj4jqdEOoFy7o7XhmqmEQuBS765H+Xr16WNePu7rbeh3OA/k3lYt7Onzujdf/w8RNrWN5a5DAQDKlU6PXixBFVveB09LXgjGGOcVwRZ/d7ioR79D7AvgcLUw3nATipz8ue5um3RMWx1Ovbf/xTGIHRGkFYwRPDoBhAlUFQAItMEDc7Pa0GOTEgYWNTqR+bWr1uO9u7YSPM+MEUS6d6VBZwOLiKjcOXgzsmOGyy7PKVUjkoFXwzjM1kIpjI70cbAQ4/qjYiaUBQBfAOoMGmyMFO+ZgY/RTNz9wHMNrRAJRHRYpv4pRSefNcGv5Edp5ABFUMt+IlW749uWLUgzA2RTZblfYFsoNNRKAKVRlFH1cnborBHxkfxaw3JiZRarpyCuCFpAKwAvCD9wEMlSogi5oEoqMh4G+Ksut8zra3UeWjZnbipJjL2rvX37SRobI9X/LGgVs7e2rWmVaD7ZKCWpQMNI+DtKEvR2VoWCDQPoqu3R0rpM3evHTBhoYKVjvcdUsd+SMWbWVtQwclzZBX1jdtc3tXFQAQGVmYeOtZrYEPozfS5j+SboBgklsFynlXA8VAsA9kxb7ZCeV/BJGU2wbVckxSo9I+Egp+lPhXVKMJJMmkxL47Qw5gzyHhiSFBXb7oAI1USn3ALDSP9/ymD8wMgNWEF75AFW9mPPjTyyFp2HiEv2bHPd8B/qkQ4ppotJgvVFRRMTs3r0bNeCyivGQOk7xKlSz/8ATgJwTDk30OaoBPrBgePfzcPv7Z31sFb0Y1McMTO2Xt1xAVrgzKepkkaoRQTRDHT/NcRKRXQaGU4SsCLAqQCUSOSLLxZkx7ghaYf1cfRBuVlHtxhnl99949e/583QG6oNT2RmXBj1oA/+BZfpOo8GTo5Nc/hKiIwEjcC5z8cBU0P2Mdnjlzxk6fPi11B6Qi47W5sR1snzzV8kA4VHGcUA0nSYQkMOsgHwCWZ0IngXrdmVCdAZgzAJMHJgCx+W4cH34902tZOZe1Ny5fse9/9zs2PIRPaNsePnlsP//sK3uxuhVA8IGlVhKMfd2ZFoPTCHaeJCqw0Ihq+wjqxesF+I6BvweCA5udfqvrBEkTPz/aqfT/faIaJXmdJ4mK/ljHioqwhvVHsKWJ15IEfuNekyTz4pyPz+TYOgzPjvNQQKmWJQBoz0bKJXvr8mU7PT1j7cOGAyaO+mo/pUycijoqKw4Oa7Z/cGj1ZlvJNqQFKky35HGfdk9Efdp7FVXqWI8K7WXB69wVk4OKpOQcA7zD8zuS5RHc97XHZzmIHcdQTQWRWgtgEIubyN+Pr8FI8Pi6+H9PVDB3ODN0L6Fy59+FqMCKS3tTIA69SfHxa4/zwJO544R3kmgZjKuvQxol9gnkqNjsT87BZ0h7EKGTYP0U1y25XFTLEd94zvTN/S3O2fj2kajw7zv2O9hn5HfWJxeTRJAvt7gO3f7gGFHBmAdySdcYSAPvmeJzOJIJMRaS2lBWAIP9jJgtNok8OR9/M1ExIH0FBiX2wdftk3zvdyUq+EyANZJBgNUkUZHcA/WeYb+JsURyT+nDngHISgswo1EuwxKtjYKFoZ6Lg1r5fDlYZfh5Hj/Hq1HcNgvvfK8YIm6OVXKe9BM3qspXJqGD94U40hl0gqioFLNWSbXkDZ3LuoqQZsk0OU5n89br9Kw6UrHy0Ijt7vVsZXXflldeWbO7b1ffumwL5865oOjIVezYDMmOK+WqUB8b4iuAULe5SvYBQ0BEFQIzH5AdQU86Vi6GM9C5KI+1fOL7fic1eBgj3iODGAhP8mDrwZyVjSoxUtqrR6ezk/KAvn/vvjVRKheoVjiw69ev2+T4hD24f0/x5+LCOZuanBQoRCX2559/aecXz1uxUrHV1XU1xxwdG7HdnU1bPHfGRsaqAu+oAoDwuP31XYGOf/zHf2Q/+tFfi6i4du2Svf/+G2qwXK2O2Obmtj188Ei/d/HSFcWXT54s2fnzF2x9c1M5EVZGKIdlK0v/MjWfN1VsLiycs6GhYbt//75yE342NjYiYEhK+nZbfeSw+AAkpbqZiryxqWm7e/+BasYAtWoHe5bqtuzquVP2Rz/4yO59+ZnNz0zby5VVG5uctnRx2P7mxz+1QmVI1iq1Zkf9S8gBAcf5oroBP3jsY7E2yqV79saVRctle3b7zl37sz//M7N2x9r1uj2+d18VBVhdvfnWm8qByEOGq6PWpcp9e8cmxqsSqBEPkycxXisrK9ZudUWQjGGVlc7IuknV7EcmcQvWuQjiUj0U0S3LIJpj3uUL1k3n7Mubd63e6okYoXqUeUQFTZZ4H+Dy6MiGUbx2AAzNhgFkAbvI67KuMgdE9K0vbc+evRLpwbgyTwGg/rN//mey91rb3LB7Dx5YHtKkVLZKPmdLj5/a7OSUC+myOds/rNvZ8+dsr3ZotUMIO4jEtr3xxlVV1Wzv7FnnKG1f3bhjqRwxf95u371rF3nNwa41moc2Oj5qtdq+KlRonr655UCvLH2kTMd73cHTXLEoy5Sbt7BUDWAgIjnAdFnJ5tQfRPYugayOzXpdne4e9QBfkCjYxhzWDgWQyiYmBfjLmNaUX7NvuVe6kwLsAVL9h6/kHqr9M/Z5DOdUrB4Q+MZ5pD/dSpXvcW3CDXtdKxcLquihOgDr47YaKgPMZqxcBPQ3W9vasWcvVkUMxf6U2q90DvqJyj34dfv99on98HvxPIuCpZifRJFDH+yVCt/3LhFHsuh16yRhFGMjVhmiH8qQ509YKO3u2YuXy6qaUaEJlrlBHS0rmlg9FypcWDtgJA44+33IHSKQ+hDILpLqCfB19T+WOFQSgN/UrZhNWaWYt/ffecvSrboqn4rZvB3uHVqmUJIdWapYsOLIkOXLZVXEK4fDugkrn+qwbWzuiPis19uqqJAjTspFqup1E1QCsYkx94TYk/NWdkLqTdix6ZkZW4awgyhQfxYXNxZSbSunmvbPPnrDrl1asG6zYbVW1zb3m7a+37SO5eyzL28JK2k2OcvyslAWroELxGFD81v2OQF0lyNIkCeidPeqxFC9GdxCBsIpj2nVB4q+qdg3ysLZyXHmN89PNqKhH1x0IAA3QXzLelT/ii7EDvETW2JLIl8snOX80fbeFj4Z+TfVUBAU7RBThVgy2A7xudEOlIoqrq9UKdvo2Lhif2IBsCWvnAFET2lvrIWG5D5v3MKIeet7hVdQxMrSGN9xz+x7OKVwttB/lIq6Wr3uNuSyWyrJ3o8xxt6Ia1Jvx4Av5Kj4KBZEoEu8IiCd+JKeePT48OoLVUiJQ+tYB1xQFpp5a7bEKNnO3oH66GFPuXrvvf5+MnXlc/2d++bsjmSsPyfvs5HLhfw4YDYiVFX16VUwIjBVJeTCDz4f7CTGeVy31j5OCewb4dMdO8LVhPs/snbvSD009hjrrU2jO2Qe+3pL2Xg1b+9cf0t79t37TyxTqdpBs2M0X9j5AAAgAElEQVR1+qtwlmYyOrvfeetdNwXvde3Rw4f28OFDq45WZZ2P3bpjNNwrWOHAFoxqwePOBcBLVMC4bdi3REV/ynz7l38qIzAXDj0WhTzymq4UpsGyN3s51PdVOXGwJ9ZXiZUAdJhMZ7cJnqSqowEZTDuMaLB5ojydg8ob47nFBGXV2gSCDQS/K7V/tydrJYB9PpugXE2uddgDeDsJQCADc15F1XKEqmjXD3WBBxAbKBNyCrZQ0CkgZUMFnKU0VE0zfdPii0NQAX/oueAgr5faetMiygHZzF2dEoMFLkisdN/j2lQlARgSBRnVkREdDJA4nrB6csXGDdGiAFl+3O4BzEZFQjM6Mmorr5Z1cFJi1mjUrFQp2P5+Xd6u+AkDuIPpVoer1jg4tOFy0b734XWFfDvbO2rotrm7Z8srmwK/hqvDCij396h8aeqgJwghv0bVV0BhYx1bPD1nczPjOlharYatr21IJUAZeLvds2aXhGDC1rd27emzF/K7xc+Spr2MY61OSWhHTfPa3ZYObRRJ/Dk6N9VvGhQT1agGdk/vYMGTsOhhvnmlRqyuGJQaa+xR4QQlD5s18++wfihCCD/H6ihNxd2KBL9CEloFzumsVSdGrEACJFLJfbU5yKQechQp+Es6m63Pk+0BykIPIqMKJgJ+GSibVt2ePHhoRwQnHVedErSOjo1adaQamkblbWKc5o5TNjw8arlSUcpLgjEOYFkmpbzsWkCgVLte0UFAiqpCNmRtyp6f2y9/9lPa+KrcW/MM5UbAvb2iYgBixmuOTTsjSM89SFGCipMyTVS/IjMGPv7xtYyBAAiV+6Je89JYJ228V4SPDxZTZrs7e3b37j3b2qkLbI3BooMYXr46aEzna3NQteJdKGKzzhhcxL04EhXJRClZUaEm3IkkyhVf3p/CG98PwBHW5NzcnFSNqCEJuljnjx89lZLPbVaCYifa4HgmdCxRi0lS8lodzAn3Fv5yDLjjSpw1DuDXoNG729E4Yh2tafy1Lugvp9p2/col+/73fs8mRoYVFIOT1ZtNu/30lf3i85tS93kfh0Eze5Fx3wBaB6ccTm68Jjb0Yo7EigpKXWPCN0j8Qr8EAVHHgfN4r85F+Xw+Ibr3fXwwlKFk+ZsAvMb1ZEVF7BkSgf7kDApERUxIk+f4QDnNdz2J1ZwkgdTe4+eXSL1AFjKG3geB2yCN71oxm7bLi4s2PzlhBO80VpVFjJRD3sOIc4a1sVXftY3tbVcR1Ru2ubUrcp3KKl1FDLgTF6qxcZljn9w7WXFyXP0/GDcRsplgKSdSbgAs+3Nyryyf2074oryS9SNJiR5Z6HES7Q5F5Hs1ku8hx9Xk/64VFZx7nKMkWYz3/1cVFREwDrd2jKiIZEL8c0DsOBET7X2IJSLxGGd1XOTatWJTeVd7+LoMJIC80Hs9JYnETkny7OSaTP5MVQhBQf86ogIVns8hX7cRWPKp5Go77iHa8nlFBSnXwK7NN2Cf72oK3rfACERNUMl5xYrbg/oZSEl+y22WZHVwnDj7bURFfy4H8l/lAL+B0I3PJS6P31ZREc80AcLtbl+YE/eCeN1xPmguh6qBWDUn8jlWuYT9ifNR5yHWEsmKCj4hsccRfzHGJNpeyecEgEA/4iPADEQ3UtlS4RfiDmxXwnlMwho3xmj95OCekxUKBoPqcbiUs7Fc13IprFN8fyJGyxZLnggf9awyXLKjdN6+vvnE1jYclLRUy6rjVfve939Pn0sFB/Ob/jqZVFb7DvFAEAK7+lmxRVz/TrASl8iGBqsOgFLUljSVD710kuIEfwah0idYqcYYY3UFssOV9ABB5CDE8G79QkLvquaFCn3wzO7de6iYv1Kp2uFhzd58400bGxm1Rw/u66zAMomeHZAY3Bf9phYWFi1bKAgQf/joiQ0PV+zwcN8uX7ogr2nWMHOrVKzY08dLqvCenpq2f/2Xf2FDw2W7fv2KvffhddvfWreSwKeerSyvCiTBjoKTAfvbHsRmNmPkBIB53COVKvSRe/Hihf4NcM/vYvGh+XF0JBtb7heQnZvkzJ2YGLfd7V3dMzE8dkXpTN5WNjdEhACiaJ23G/butQv2wZsX7evPPrHziwv25OkzO7Vw3lKFiv3oJz+1oZExNa7tHGU0R8i/AKwBGqtDAMMtkQRdAOKjlr395mWrVLJ2/9ED+8M/+WNr7x+oGuPu55/buUuXLBN837Gw5LmWhoZs5eWyjVVH1EAbEHbp6VPFVF5VzjzL2u7urp0+Q8VLSTnZ8Mio9v9PPv6VV7FUx2x7a8fOnjur98Cqq4JwLZ23X312wyxT0HOkMp9nRKVBSueWi4gQfFGx0qwf2vBQ2fZ390Q+YSdC42+arkPM3L33wPYODq1YHlalCkKnfIa4OmXTU2M2NzcvILpZb9qP//ZHUq9PT0wof+BZbWwcmuWz9tabl2R/BcHAmt5YW7WZqXGbn5tXfJ/K5uzGzXuWKVRU0QMxBXn1+MkDt/80VwpvbBBzeoUIqmfmC24CfBULBVV95EtFWe9+8fkNqXPjuhuuDGnvpzJH1Qrk31SV0S8wX5R4DcGhGuUemXJS9m16NwI04nWfQYyEXXGr63Y/oRogWpXEc6Z/xijn50wIjYM8aAl5Qeh7RE6PXQl7JqYF5CpqEMsuFOxwdMayf2QtmzpSf5VqpWCNw32pt+cXzlhrZ1Pr69Xalt1/9FyAu8D0kKcziqxzNYiXBRRNoNtBLJjxCgzOR5rdBhyD+9EZRawX4uTYZJnrjGeq9lrtkexN7FFOKvP+VIFgoTY2Nm6Tk1MiHnnekEXLy6v2dOmZKqcAhFnE4Bh+1rpYirUhgVeoqOAeHANxtwuAb3K38dFR7b08l07Xx41soFDIWor8zHo2Nzlq3WbNxiBPikM2Uh1TnHnr/kNrk/PT6Bpb5qERVd8PlyDbUpbJQ6i+sGJpWMKysbEp2w0WTB4ju1Uoa5RzFTwhnvnkfDEG8HPERXFuY8N51bVCMW9HjX07M1m2f/bRdZsYrVh9f9d66Zwtb9VsY78pW7rHSy9tdWVT7hC7+zX1ygT0VW4awHMqC1i7zB2J99Sjy8/GZOUt1x0r/ZlXIsxCrKTqGIkanbRTH4BAVEitLkeMQdzN86fKTXZUkOlBQMj7cZ+s3UrRCXP2s1yapwHGU9dzAo/h7KMKgudOlZdEraHCjvlEjr1f29daGp0cU0Ue6xUhrSzpsKzKOlFDJQyOGmurq7onXi/MKfTnUHULOE+hqLnjsZ9XyQLYY1WOiINYlBwDwh9HBu6Z9dum8gZxbrsl4hZ8RxiYHBvk66rxZk9ShglJTMUD65m+p7msLMARZsjxI1aEWloWywhgd2uHlisUlRO9uvV2P/OZe/MrrVnlE8qbU6qqYRxksw2WRZ+HmLuFmCTmreyZwg1bVKsGAZgsXj2vU3/cOkLrKAb0PCjGrhKOkY+AHR6Znb94UdWM29ublrOujZTz9salRZseq9rM5KStr63aF1/dsp1WyjLlijV7XStVhkRgv/HGm3bt8lVr1OhH4Wv+Rz/6G+9fESqcsaiHHOI5QWqxZmJ1u+LQUHElq7jQ30LX+q31UzKt//bv/xRGYIaeDC2YUfovlHRgQxSIQeWQDH0B2BghDtjYWCTuu+t2Rl6K6sCKDvgQgABkETCyYQNEuhcvShff6LVJJZTTAkYD6O/Jfkq+hsQ4lJDDHpP8sLA59Nks2YBJgFbX1nRIOZLtFjMcHix0gjIFF31/QM44T7rZmHK5Qp988MT3eFLNa2NyrwZHKiNrD/xCVVJLwullgAImxMz6ZzCOXAus//j4uIITDkDGm82PA+XgYE9JmBJZ3r/lPqAQLVwRTeBQBRmWF4b67ZUaBZKQ8B4oKkr5rAEozk4O29VLi3bUa1uxXCGSsgePlmzvsGF7B3WrHRwGW4y8vCYzWbf3SashXt16zZotnJq2s/OzdrC7K+WKW0ZhMdS2ZqtjmXzJ9ghM8iXbOajZHj7+bLIoX3sdO9jfs2Ipr3vyxpCehFNdce7aVW24/oz9/wT2heA2lgp68uolrt6LxBskcYhHIDEGinIxCb0RpDBpNuxgb0+EBcTJ+OSkgijmKcEOZIWmXjptYxPjUkHxxTwnGHQQ6sga2BkB5oTDkeA7JubMRZ65QAfZpfn9cJDm0h2r7Wzbi6dLdsRrOqGZuB3Z8OiIzczMhXmWtnJpSM0eSVBRA6VzJSUQVDNINd8L4Ga7ZQcHmwp6CHbxNHXmnx4rNas1Nm11dUU9SphrXoYMgx8C7qwDfhFUiE3BUDYolYsPI/hKQs5RJcMcVjPmoIaXMjWWJ9M0V3Zw3pdFwFloJOu2Ld74kCoRguhHD5/Y0tNnUgD68Pvaie93ck/9JqAcqym+WRGgwztaSwSArg8wSTETehYoSA6lnX3FsIMkbm1lSvQAAs4tnpNFD2oUcKB7tx/0ffuTvU0G2FUMcmLDareicpU5n5lA36NVma4tqnp8b4xuBUmAr69QO0JpzNJ1diKT6mntlvM5e/fSorxeZ6naobFYeP6M8W69Y3cfP7effvyxvVrfsKO0B+KArWp9krSu4ZIFHDlIqasjKWi1dP8qV5ZlQJjXSgiCAiUC1wGYj+rt+Gz7gZ8Cymg5RjXTwE+UBCSySnEOcP+RnEnOk2i3FkHLWBmhf0eVbqI8PrLTA/V52N1F2kdFdyhd0KPzvw8ANgebeZLyX5WlH6RGSqq/SxcW7eK5RSvlsnZ4cBCULk4sTk5P2dVrbwgcg0iemh+3v/7x39tRtmjt1pEd7u3b3t6mNbsAUl4BdhLk1Xi4PrAPNkfCwYN4t3Xyqe0kls7bIBwA2OP3IunlZIzP2zgH+oD4EWX/TVf16Fd8NvvYOdGvdRyspByApsLPQXCvHPL/kiRWEnD3oHtQlRSfrarweu3+3gtYFn2CJVZQw0Tvd+GC7IE9F5aHfTD8hPUTVYlRbebXFa0rvlnFEMc+/jmo9Ioka4gV+oB0uPpIXkawhF4AAWyPe1JyvgKgcq4B0LkVU7D2CGXmg2QpcY3HPP792fQrmnRT36yoiF7kfctFFGokeALOnaiQJduJfkaDcQjklpuO6/PUGFKij4HKlBiNMzsCFXpGgZRNjml8dlgGMgbu/3zC+qnf+Dv0aYpDHJ55YkftE9H+Kx7LRXFDnA/quyJQf+CF7jZwDpZp7EMjZ83voMjlHSWYCERTWAghmcXayc/awdwOFmlh2ZCAEhP6WHujTHZWWYCIpEBl6TEF10wlrYAEiABZjgb7x37MHHtUJar6ws/Y9yvFnI0XKWA9srzA/65ihuJQWdWxKAOL5bK1LWuffH7bdvcRD/GeHcvkUvb+Bx/Y1PS0pVKopulHhorZ9xYpln0jCE0hvXF9n5QMZ8X6BkQFRElWcQJxd/L5J8UPPud8DulZiFDN2drqmh31mmoM7cpBrD2yrhKXpziATcGms6OWPsraw8ePRQggPsE66f3337W56Vn74rNPRWiclc0mwhUUv3W7eeuWLZ67IICbioqHjx4p3t7Z2bKFs6dtZnbK8vmMFNE0rr5354ENlWmyPWf37t22Wm3P3n/vul24umA7qyvKWbBEvXnztjUbLTt9+qwsVGRnkcnrHGBMnr94rkbfjx49ltXUxsaW5sHExKRyq9HRMbvx1Q1V4GJhNTs7I/EP9iz83qn5edvbJZegcjmlyoXJ6Vm79+iR4gfiU64/3WvalXOnbX58yO7fumGXL11SFcnCxcuWLQ/bj/7u720YuyQFFTkB9FnsPIPqFFU9liJUvncaVCj07J3rV2z51VNrtev2wz/+I+up/0TTHt6+bViCVKvDUmMDupHfkNMAxlVQmAdVPnEguRHPkmuHCFHftoUFGxkelj2bor2M2ZP7DwR0jo1NWG3/0Gbm56yXTqkysTg0ZAeNjv34739h7SOEQBMi19lLt7a35BEPKA8oznVhLSM4KzTcRXHNflUs5CS0AaTb26/ZBtXihbIqIlDKYw9VyGEd40AnamfGd+nJE1U9XDp/QeuLZuTs5VTfcvh++J0PRMA0Wg31Inzj6hWrDg/ZxuaWDY2M28e/+tyypYo1Gm095/lT87aF6j7Vkwqdnn+4FgBKRhIXcoXP4QsL5I3NTYHKQ9Wq/eqXv/K4RMK8vEg6eitS9by1tSkAHVsS9hWsnhTjhZ4L/P7a6orel4qWCJgrB2h31cdga3s7WL6Fcz80oVXTXeX1ELaIYNzuOWIDOqujpV/YnWOltgsc830g3veWYDPZ61mpkLfRkYrNTI7Z+HDZ2s2aKimq7GVpgGmzR0vLduveU8titwtQnyf/9IbKxLmQszwft8BCYEX1osetbqOS1th4rE+/zOjf7/u47JZkUR324dA3AHGhizjcaUF5PKR1yCfUhzLL2V5Wvo7wErJ1e2dHlm7q16McwPEQiUCpAGrzXh3va4TlEeMJ4UKOQjCGwErVVYDFnF2IYZgjnntAOEBSD5cLNjFSsb3NTTV/R3XvxHre9rEjoqKiUrF2wCg6rSatwdTHh4qzcmVIorKjFBUDLkyNtkgeo7EWysq5exLmuE2RzvIodOkM1OmMgfJoxLHMQWvZVCVj7109awvz03r09c6R3bz3xLrZstVaR7a2sSUbPcDrOvhDoSDxFTn9EZX6PD+AWzk1uFeozvCAI8miKZBKzFGPfxgHFw1wDy5cS0nt75ZiLraI/QFkORr6QDjG43EKPWVYqx4b+jnIecm1QGTKtiz0gKOXEqQiRAvPC+xNoL4akAfBV+gnFW3CJYZERNxpC6dYPH9evSNkyQmR0WqLACEP4XPAgqhY81jFYyqvQmgFiyBIMNYa2EbQzYQ+B4qHVUwTevmxtlWVwXnfU89N0DDMxXpdmnAHoqPb0hnhWA02UL43oP7XuFCBU6DyySsyiG2oKmMOED9KIINlWOfI9ms4h6REmG88+CimAzYPUUHv11Dp4n2uyJVl4qb56gI+t31Vvsw8QHAqKyhEFo4Dan0gWJYw1nv1xArgSL4OKptjTx+zzFHH0sGObfH8Rdve2bb9nS3LWc+mRoft7WuL1jzYs1wmZRNj47a+vWf3XqzbYffI6rjQ5HJWHR2zy5evisBkzOjZAc73o3/zt/ZkaclmpmfUuwOR5KlT86pK/eSTz/TsZF+WzuhaB/b03F+opviWqOjPl2//8k9oBEZqhwL7HZx1ZRiJEgsn+vVFoAilCArr6I3JIcqGF70VpYxN+NERWFLyyjaiTSEorWMVQwT21fgobNQw0Pw82lFxwBBw40lKYOaCRGdtCYL5ZT6fDYPP09EE+N/tSjXPfcjfs+vMv6yHUMNL8VCQbyIKklhKJTBMpcIo1xwg5w3dU9AVDzDB0T9SJf+yffLSTCpF3DaBRml5seh8DuqUyICipsIHEEUM36fvBkopxGruo+fgLmp/khKeDxvt9NSETUyMiZHe2du2l8svxSg7MJ6ydK9t2aOUFdJd++M//Eh+wKVy0SpDVVte31BZd7Nrtra6bsvLa4atYa5QkYIfqyFK0LrtmqU6DTs9O2ETI0NqblUdGlaDJrocE7SgxDg4bGJiap10xp6trsqDjyAmBjA0yyKIaTTrSnq5PzxXGaOFK1f6FRVxKUUA0g/EaHngTbmieiVWt8hPMtGM0UFu7KRoQOmKHPphHKgKBfVW0cYmpzx4TKetWKooycATkekyNjEpZQNfKMgGTZdMRFsf5FMTLm+qzH/8PYLs0YbHgyEO845tLr+y9eUVM8p6sSXDDuvoyKpjo3bq9IIIL6kRsjlVMI2NjlpleMR6AANdrwrZ3trWn/uQLs2GFfIkSaFaJ7zWy3wP7cX6SzUrIzEjIScwjkElqjIdbKERG9cvW4cA9shrNvTsiAG2qo9IahR8Q1Q42BTBBdZ65sgbijqJ5eXHTH/Wqasz6dFSsmymZPt7h3bz5h3b3sJOzIPYuLfIPqpvAREZLP+844CyExUKwMLr4z14qeYAyIuAUf/1mSMvj1UnKwekCcKwD8jE5mg5Jyq4J6wWLlw8b+1e25rNjtVqDXtw55GDo0rCIF3ZcSKRGUmKoDbWHI2l8LEkNQK2TpxE4DeugwjqkhjwdZKo0L32MlLbUflN03r0KpVCVlZD7125ZBOVISuXsRJAdeokLJ/U7BzZQaNttx89sr//+GN7trJmduSWGhqHqLKOarKozmW+h32dNRjXB/NHwCj9Z0Kz9eR6dtDK7/F4KX0gqMKzcgtAVGgkuqGBYCA5TgLaSQXfbzqG42siMOrj6MR3Eop+HVGR/F7ys1VJ1S8fd2Lt/ffeVTK8tb5utb09NVKbnZ6ymakpqTRZ9+zx2DiQMEMav/n2OzY3f8q++OorNTQ9OmrbzcfPbGTmtF1cvGxff/qp3bn9hbV6DUthn6ReD0koNoxdKEvW/EDjEyqXRA5EYjJR5RfnlYsEHDAdNFLmOfkcVgJ84svB5qZRmxXXVyQI+vMWEiRUzrgdQqyUcWCTtR0JieT9SP2UaAh9/Hmzl3slF99n7kWiQlaSIbkMCyWQUp4gZQtFr3ph0yL5D6pFV1u5BWHcy07Og+Ttx/Xnc9mTnrguj//p4oj4Fe81XrtbWg8EEMfuM9ggMG7s2T5WQSJCBVCiJ8TJcR/sfX5dfcKH5DZUy0pEEQidkz0w/LzyxqAiaaUiRanod5IklzRe2H+E8vjkuRz3Yq+aHezZkajwnw9IsyRpIW/poA5LXqv2LZWK+X99EDwMcjwbftM+EMnF+Jzi3iHv30C0xecT75XfkRI3YQPY30+k4POeKCJlZPvn80sxAiSHVJU+eMln7M8GQCsSd25bRJzHuBCPEuN5VbKrfmPVRQTGvOLJif34FdpkB4UqdpP+uYiNAPLGisSDKStJiEJ1VF32koCa+XTKCuVh26237bMbt61OcKhr74msQNn+zrvvWqfr/YSwMWKfZl3FeDnOn8E1DogI7mVtbU3XE0VIGt9+vxx/L/1bTLlXfUQrkUwGi5ucra9vWq+DZY0rX0VUqDLaCQpiV/6cy09YLluwG1/fFDCCJQcWTB9+8L6NDFftxpdfyEZpempK/QioWkA0tPTsmZ2aPyOPdipAqKjg9w5r+3b69JyNjY9apVISSV8slGzp8TMbH58QCCbB0O6Ovffem3b56oId7u1IrQoQ+fTJkgCHoaERWWhgIcQ+C9gEKUU8Nz0zrX4RQ9VhESGQEhvrG8obzi0uyj6Cv/MFGEg+BcFN7HXp4kV7tvRMCuf5U6dVkUdlxdPnz+X1TQXMu+9et3SnaWdmx21mpGzPHj2wudkZu/vgoZ1euGDZctX++m//ziZm5iRcAIzc3N6x8clx5U2cX0Dz87NzyguZM71OQ0TFqxePrNlp2B/8yR9Zqt2xw509W3r0UD0Gp2anlSeifRARRyVPNicy4lC9JnpqkM0aIK+kIn5qckoinHML5xS3T0xOBPFC1z751a9sfGLKe+R0EcfkbWJq0pq9jpWro7ZXb9nPfvGJdY+yUq1GQAfFq2Kg4FE/NjqiPIFqIlmFSFTX1HVOTU16hEBFPs/v+SurVEdtZx+CpSKSodNqKK8i3p2bnbN6o6Zn2WphJ9exK1cv29mzZ+z50nNbXVmRf/zbb79tz148D2fukZ2am1V1A9U7IxPTduPmXauOTtrmzo4qjrEbfbb0xCrVqqpGGq2mHezuSdhGDkql+OK5RVtbX9O40iuFOTE0Omz5Yt5++rOfO/FS9J6EiLKwXmsKAHRveOxhyI3Zz8ltyZEQO7EfQZag8j91+rQIJAhdehIg8IKsWJN1EQ3cPX8QEJrF8cABxwgEan8WSBn6m4Xqv76AIADG6k1Bw95iUapmHkbcq0WAd3s2VClZMZe2hTOzdnpmyrbXXslCbKgECMxyz9rdR8/s5t0nli2WrdHynhiA5hL40ZdHbgCozAFhvcIQoSLkmVsv4/1etFaz4b1QgvgsBo3R/kVnojQakBbUrzspw7xkjYhYyKJcpxo04/a89HUQ0WHWoqKWHkmqbvXcVVZliuW8Mp0kSuK4cI4QEwBYK/dTDwoH5L0IGvsdYnx6fLhLgHJUcr1U1yr5jP3pH/7QDnbXbXN9w3a2dlRthe0YpjcNSJxKWaI0LpA5y9nGvHr58lUQouTU+J2qAvV/oWdNBVGFO1xgFc6+3JB41G2V5SAQ4r5oleTNgL3nEaB9IZu183NTlu3s2dnJqp07NSMi7NXatm3VWnbQpqdS1prtnkjp/cOGbexsizCjfwKAPymW+huGfnmKE9LmxI72IPYMPzMVB0fBRBCRRNGO5/kpJ/Ah9kIzcO9hQPNp782XVPQTT0JUpHKE+xBxUEr016FqgB6V9E2gcfSh1irXUyrmDJSDsRE5YWbVatXKlbJIUkhR9kyvzNoUuYYNUrFcEvl+9tyCxENRNBwibe0/gN70Z3314rn3yFBuZY7xBXsx9aKhrw72lyFm9zZhXtmD/bmqIIgbZb/qBCOC35FKQUB9uwnwn7a33rps8/NzquLw3rA1XTd9WHiNPkO4nCdhEgiJ5GD9MQeoaMrrrKZJOxUckFHY4vL3pS/e7Mc6p69/1Xdz4dogWVlTEP+cyy5M9sb0/DzeL7EAJAX3ze/y5YLXnM4Bd1MAe/M9wXPVKMiKlcfeTzFDBRHxbzqt8xniF5yJOzwzM27nz0za2vNnNjk+qnihl8nZ45Udy1SGrZtO2drWts2fOWtvXn9be8j66rrGenNry5ZXl9UT6eyZBZudmdN6qh8e6uy5dfuOYpKvv74hkTaYpdv0ufUfRIUTT99WVPzGfODbH/zjHYHJlgMBLCo1fc5lrEmwEDzfWCQ6cNNp293dUQAMII33opdqumcqC5zXA6y7eJjUhpBu0JWeUSK4QQHAhiWgNiTXBN6xrAn1h0ru9J6ucGBTKxbcrocNhY2nUOLzGjqoAbefcw0AACAASURBVJSdMMjo2qK/P59DUCj2vpALpWMpu3rtqm1uboitRFUl/75sVn9GsJo78PJLrtlVTEq4g4JUm1+rrWDSG2y7Klt9OhI2Kq6iy9nExITKkbkJvFMJxlHGr21u26n5Gau33c+xXB6SHy6bpXz02pTo0gujaePjI16qvL9nr1Zf9ccaFVPjoGZDhZSNlFL2p3/yQytkXRmAamVlbV0+eSQkvc6R3b37yF4ub1kuP6SyadQKhULGivmUZa1lM1NVK5PsUlK+sWGlQlHN9DbWN21kZNSKw1V7+GzJ9vG0rZRtdWtHjH/jsKWDqNmC8aevBcx9IzQ/omy1Z2cDUZEEbiJREb2PI4gUgYtIUvDz1xEVCkq7VG44UUEycpKoUCUEFmMKBiAqHEYdm5hQKT7vwQEQN3zmMPeUJCqcyXaiIoKzsRogAilKvntNW2F8dnath0Kli1IGj08nKhYWLvh9QMTQtL5aVZCBSmR9c9sOKAkmIafKCJ9C1mmGChvIjYjdUIqOPRS9WNr2cmPFltdo2pfVfCmVKt6Qm7JplA+hMihebwSauT+pDQIw7oFbOrw2NPMKih8HqxxsUYDU9aTCrb1cEUKcqBJ1qYoAywENC7a09NIePnhsjbo3XGcuxKAiaZ92EmiOZIbHl7HJVVLZHUA6KV8HIE4M8uOfvQxNjgk2vFrAAzGa4OL67e+h8l0B62mrjgzb5SuXRFSgEnn1as1ePVt28F2f5V6kobtPqHFXKOsHgubXwLOc33QA1/FTwEtX6w68ch1QVubVfx4R1NPvEWSJ//GKNKopRipF+/Dtt+3Ny5dsGJD6qCNAQM3FYkPh4H9bp1dKu22PXryyv/nJT+zVMs0y8bjuGfVQkWgOpV5+DaEaJI6jP2MH0gRaZr2cNqqW4nrx9eD3FxPPeC8CCKNXsZp7e3ApP/foU57w3I+vi4THbztxdfZEACwEyMm5EF97EqCO8y75PAa/643mvJICkCNvf/of/In24ubBgR3sbMv+gcSLOUR/mla9rubZrIMCe87QkI1OTknZ98VXX2r/YL3b8Kh99wd/YsPlEfs//tX/ajdvfGJHqZYAomh7lgRltWZOEBV+zQH0kzL+eFPgmIxp3fZtmhj3CJ5/k6iInymxQLNh6dDHRcr3WMlwDGiMtj8niIoEuXkSaP9tRAVrrHdEub3HE646Z4/3hp7YGvTfr189Q6VRRkm1XhcbNQfFf1hBfk6EeZx87nEPjM89SVT4PhRim0QfA5+b0r/1p2WcQ3F/894fxys1+58Rqib4N3sl+70+R54PTvgmz8PEhwThxqBEvU9UqGJg4GedXLMnAfS4R+hcEOHkDVKTX/1rR1mZWM+RPPI1577bybkaiYrk3tAHqiIRq3NksAfGGMDnqlucRaIieTb8PxEVnl8PKpIUSwEQQ3JpQxicP/E5xaqjWFGS3CN4L1lGxA08kGCRqFDlBrGByO6TBLsDtjodAlmIsMbjVNJcr1qMvUQieRTHKu5/J+9ZR1mwWPQ+FS7ioaICEG+inLYCMU8ArlD7cnZQrAWgnK8M2dKrdbt9/7FU+V6ScmRHac6Qsv3+D35o6azbONQO6vozEhXJsT1JVHDdjDXxdSS2vBn48Tijf386D9x2zokKxEGARXkRFd3Wgc5k4orYcJb3Yh/m+mjgfCo3boVCxT7/4gudwXiDo1imamF8dMyePH6o821qYsJmZmbdWrbrfRZmZ2YtXyypqfPzl69k34TYZXFxQTZQKECJ1U+fPmO//vgTAbrvvvO2/eKXP7diMSs7oPfeu2K1/T3Flpxj2KWSC2xsbtvCufP25OmSvXq5Yh989JG9fPVSXvXvvvu2iAhyDgApVVFXKiIZAK2IR/ElP9g7sPGJCdvf3xXwRhNPKS+p5tOay9ruwYH1jtK2vrmlCg5iV/odYEtxenrMFmYn7cXSY5ucGLc79x7Y+MycDY1O2V/+9Y9tem7WUiidqcSQcrjnoLGlrFKuSIAl9SeAf/PArlw6qyqXRuvQ3nn/XeV1++vr9vLpU5scG1NuRaP20vBQqFZOWY9m2lT/Njt2lM/b/Zs37cL5i7pHSCNIGvJHgDoImvnT8wJqqMJeX1+zoTJiIgBbU0+LUwtnrdFp2y7zMpO3T7+8ZUPVScVHkBASTWFH22yKrFBMSkVzpWyNQ6okilov+KqD8GJJRWXz8FBVvQTWNncslS1YqTJsewcHNgwwax3b29m2aqUiYDJfymt/fvL0se6T5/b29Ws2NTlh0+OTtrm+LmKM6wccJmZ8+803bHx8TE2vp+dO21/8678VYUH/GIDJq1cu6/d7CNDyeVmVQR6wFzYOaYDrQDQ9JKlQArCD4MnkyUna9utPPgkAOABdTvczJzDxIPTnaes5sFcDYPKMAfHIkzlb1deDnCGbE9EHgEquAliO7c6B+g44sc3z4n3Yc+pN7KNyAUx0qzaR06izQ2yOCNCFM664j8IH1jTz/aBec6Ii7VZg5BX0TRirDtv46JDNTIxaLtWxtZdLdv2ta3Z6dtr2tja0dm/cfWy37z+x0vCoVPeAl1jjIprDrlj5TujlRF7FemrUG4rBqcyJFWECOCWW80brsrrueCWFN2X2Rr5sleqByR6kfB91eLMvuGph00aczD2jYO90bH+fXo7s+4CsnEXkTCnhLuAqvA9AP5/pVR6eK6hBd783pvd4IO6OojXOOlWWFegx4EIq+niMV4o2VMhYKZeWLTRzq1CqiIh79Oy59n3swiDYqXiPsQCqfPrDsIYgtBBEYqeNQwXzgbMM4LrZqsvOR3evs9oFKd7417MH702Q1zofxv4qWGoT5ODpf/7UjDV3VkWqj1Ur2pN3ai0bmpy1Ww+eW63ZsvGpKZudnVMM/W9/9jNrMyb5nDXBA3JFWeERH6L4lyjWPJ9RBUCIzzx39ErkSAIhIFIVBQ4hIe/lvopF7Ln9vOG9Y67v568LQgCKwVZyJeJ7xL68V86yKSzU23bU6VkO4U+nZcNDBTs1Ny0ShDW+s12z2mHT3njzosSykLrPn7+0qZnZ4LRBY+muKlp0xmcywnwgcU6dOa31CnHDenUrcoRUhDQ9WePRN8FxCu8dqcboYR/kqTCPeS79/CaIjHUeH5mwCNYBlWm8cTpFVVPOaruHymsnqzkbKuft+7//fbtw6bILiI5M5Dy2gtzP9PSs5vdwdSTYaWdtbHxc4Rz4xquXL2zp6VI44yo2MTll8/OnJehaXVvXmvnf/yX4nn/9R/8167BjDx8/0nkRS+7Z78EeJQYrlXTdkdwvgs3RODxYOnmfL49BFPOFfmD82zFHJy1ivDrIA1x0h6CRPBC8ZOHsWdvcXLP63p66hi3MjNm1i/PWqR/Y9OSkPcNNI5Oz+883rDw2YblK2dZ3d+2w1bah4RHFKM+XXug2uP5CGQeatoguBlN29lQvae1n7E//9E/t1q1bbhfXbmvcONdiA/coPv3W+ulE8vLtP//xj8B4wz0Po78yC4BSNaoAANIBYrQ5w7w3AOCzYnOpOGCzJlBh8XuplZMILK6YcPkZ4b6++oxQ7RCTRj7HGy65MsFV0aiHKsEWyMspYyLENXGNHHzqg0Hio1zWFzNN33QQQiDQVDiTVuAflb2uxkrb2YWzdvf2bSWt3oTU1VoKDhQ4EMDFQy1jQ0MlWU1xvdGrks2Kz6W8HVsqfsa/OUDUk6LBIY5iDr/eppKfahU/SQLEvMaRLw6QnT0a0JHcueqCw5oAlA2XgI3DE+CRwEnESyZtL5ZferNyAj8O7IxZ3tL27htn7PrV89ZuHqiJIteNmguQMl/yHhN7+w3b2q5Zs4WaI2MH9YaC+Hz2yHrtA1s8O2PDpYId7h9YnrJ9AFTELSghcqh8OpapVGy32bAX6xu2x3ORh5+vCbBWAjX56+nPtqybSDpOX7wU1BYDtbADBKbnpvAm0ViZuRR9L528+mZFBfOMIB17A+bQbyMqAPBpNEjwxbzEFoqeEYxj9GcVQIiX628hKpiXkYGPCbcTdJGoeGrtesMahzW3fkLJe9SzoZERW1y8oHmJpyRzDkUUibDUqByIoRcKSam/p49JvkBFD0kCyg3+nlEwRuC402rY46dPrFFvKsHBUkqqTZK2PM3hHQSOasSoro3AUzy8o+pRwALeli3IRyck4nOJZEem5xYy8k4NjZMBGpiXJNBUBuBx3Wh07fate7a2tuWWNikHsJMAUXIM4xyIYEgfoFJj90Fj7wjMRUAJZdMguBiARYI+0qiMj4x2pFJZS8lsshAohERg0GSvZ+VKyS5fvmhEIWwLDx48tt1NfJ9/d6JCddY+o/UfREUE9VTqHUDfeB9OVLiqOTkG/D0SFS2UXJBLWOAVsvbGxfP2/Y8+sKnRUes2GuoNgiqL50eg5nZWJIsd66JyOTJZta1t79lf/NWPbHl1zbqpjLXVpTmAexK3OpmjBEn70nGwNZKL2ZyTzCeJCicVXEUUiQonL3y/ThIVkcBR0bEatiqt6AON8fnG9zkJtr7uJNZnBXInCRzH5xFJotfNlzje8WdROe2KIF/3JCHsxXPjYzY/OS4Vs/aNXtsqhYLsKwrlsnHCqI8MkyibVbLv/W3MGr20zSxesj/4D/8Te7n00v63/+l/tCePblk631EVVt8uKDz/uB5OEhWeQAWrGzXFHvQKiM8wEqzR797VbmDAXlEhX2j1QAkjlABbBVp1WeMDQFkFU7H/SACTfX/4zUTFN8ih31JRoclInyNhyq5idZsT7/dDxcqA+BAt4XOLxqglznxXe0IER2sin1OuTIwVYv6sveFmtMlKjkHc8yJREdflcbLGq1+SXzFu0e+FfeB1ZIWiq0DK5XNFVaDxpcSJXkeJ8zD5/icJtQhkaG0EoiLGYbwugt+qvjlBqsQzwXsaDerSkveu9w+edJGkZN1HYsF9xQfnhFRtKOMSe0Nc+3Ef0HjoZn2f5NqTYgVVeMhHIDSaDGX7cZ/8bftA5KzjPcTKX1VFhliU5518TnFf8ng1aePk+2KsqtVeyAKOZEVoOMkSpArRX6s76j+yQX8PSV2CxRdgArZIgGi+r6jZZAAjTxIeybNa7+4hdb/KWPMdtbOIipxNDectz1kBOBMsMQAe8J1GsEFFxdd379uLlQ1ZaPRrIdM0LTP78DvftYnJGcVKVBSKlg8VFUkSxUGeQbVEPNcBlBlf/h2JhTggMabXHAhVLKqoEOICUUEz2aKIik5rP/jA+x4Qq00Yt1TOiYpLQ96j4ubXt2VtRZxBjP3GtWuyYbh757ZAHSoREA09ffJUecS9e/ft3OJ5Ve+srKzZ2samzk6A3XPnzsjCFOAZ3+8zZ87YjS9vClQ9feqU3bx1w1rNur373pt29eo5q+3tWGW4KsuPp0+eBUvLnG3vYoVasnabZ5uTdUez3eyLjqis3tzYlGBlaemZzcxMy/6T8eNneNyT+6yuLuuMYQ4vLCzY/fsPBP5MTs3KNqJaHbMbX39tI2Pjej/il1IuZfNTozY/OWrPnjyy+blZu3v/kU3MnrKxmXn7y7/8GxufmlHMtlery3v7/gPed0RE01EH0GlGVh3N2oFVihk7vzBva2vPLZNP2e//wQ8F3myvrqmiYny4aqMTY5bNeuUNFkwox/e3dmR7AaAEwPvg/gP1pyBfBOCGqKBqnkqJ8TEaiB+qJ16zXref/fRnEnDp3ts9O33mtK2sr9nm7q6lC0U7dea8ffL5TYHUCAHIj3b394ONHH3pSgJeISLwlKeKYoRm0fRgzGRsqFTQ+a2m6fWGejGsbmxbNl+yQ4C+FIBfw07NzVi95iIiSDA2L6qs2r2O7R/sSR08VC7Zdz/8yNZXVuRVLtBph4bEWasd7NviwhmbGB9T5crI2KR8zAuV4WD9tGOzs9Oq7Mnk81YolfTcG4fuSc/OQS7J3KP/hgR4uZzt7e6qCgZ7qS+//Fr7B2ApleIIy5jnO1tbVi45OUMODPlEnw3ZrgQrYuYlY8LeWR3xJu6clVqrEOiWUo+2KNDTWqQqQDZqNZED7FFScyundntI7WuyW6FyOllx7GcNynJy/oPDmpTw6p2IqjvkdKPVYculurZ4et4Wz86JqKDiv1jIWLVUsnSuYJ/duGs37z230nDFWlKFuzBNRDK5SA8bSyrkzfYP6uo3UiqX+vsZFSuuxHbf/Si+lC2Q1EG+9/E7Lpgrhvjdf9ddF7yPIsIxrG7Up4FKOc15hAPkHcHqiWoWLLGjnWA/3nIlU4ytpO6OwQnnuM4W/xxuKsaI8djXGZtyKxo887dWX9ip6XF7/vSVGk9TjbB46YIaAj998UqWd5BxiGaY1456pKxeb2ndct8AzuypEqbK5aBrw9Uh4RLgRfXDmvqYIMxhLccz33NV1OzBeieV0pqX+LPVtGqpbFcWT1sp1bGJSs42VlfcAqiXsVo3bQc0WM64BZWqF0plVVTwOVy/uHXOLTWT9rHhH6xJOdkRiwa7nEG870SFznieacj9IvCNABZ8xvEqd8mgcTQYT6xIVoPqQPJBVOSLOWvWIQBD1akIrJz1GI+0N2C+dmXRfvCDj2x3Y9NadXpK7sl+bHObvnQ99aqjWTkVN802WE3ZnwT5NZaHnY4wuHMXLqj6TpZ6GcfhuE8II87/vR0qMdb7ldi+fr0pO7+nChiRYf59xxxwpHC7cjAJJxlZOm41nk1TFdK2d986Z9/74AN7eO+OCFuwE8hH8pzZ+dP24uWK3bl73yanZ+zswjntUVNT08Lp2Eti1Q7Wd5WRETVOZz5ABGMNmIUg6fa0x1A98q/+OwgJ//rP/9u8rPs2Nzbs7r37sk7TfYQUm3msr2h1q+bnNNP2+MMFlY4lEXOoskqOKY4vsqa9qj+sr0SwHeMwsiRGC7KY83d9dcWaB/uW7Zktzlft4sIpy6V6Nj5a1Rm/trFjN++/sJGpWSuPVu2TG3dtfGpUe8Hebs0mqFzcrwmjwS+LqkhwP8TJfKlHjWzG3H4LZxlIGsduYnVPcNkIZ8G3RMWxNOzbf/xTGIEpSrOkeqCErx33apXy8W+azomBDAclmyjlf17W5X6xsb9AbDTMok+CVoUSYH0gH/D0gz0s5BWI8EXpM8EAiy+CHwQY+HpCYgD6E9wSbHEIyncueA5GL06CAVfQuboj9s3g95Q846vbaUn9gDqU+1W1Ac3BVU5O821XCCuw4tDD37E6Iq96gg4CRoIZVBhuldPT6xw8Q2EAgTJQjUEQoJwAQFeAEso7Y2kZ4y4PzSzOkV0B+QTwKBi4BhRh0Uwili7GUksOGJrnESwDLghe6jTsyoWz9nsfvGWZTsNah/SXwJsTNUfbaq2mEk5qJvb3W1Zv9AwHp43tAx36qL9KhZR1mvt25eIZ3T/vC0jZbTZtqFhWWZ98TXMFO2i17FDe9w2rE6yjyOh5nwcAY9R7JGOAlfydSIJnAFERD4u+Kjt4nKvJ7AlAlKCAMeQ1CnZjfwSBkIEYCESFyviCjdjh/q5egw/zKKX6AvBIWoZEJqEgI/CiwgE/YA5piApZQwSiggAhCS55OWsE5/1apeo7Vqabtubhnq2+WLIm/UAAN+XR2VUQBpCBMm9ibEIlkMyh1eUVgc/yOlVTXgdwpOoI5I2AgKxZWeAzZesQhASl3tMAGIESwhcvXmlOujo3EBUFb/bJWhKxKLLMSzJjo9QkCSFSJJ/XzwmQZGuR8JkX6IV/NiXHNC9v8ekeELjPdNpS9MRIu73F6uqm3fz6rrVa3lwyNuyNz7oPooayzSQAFQFxR7J8HOOXkqIQ6EfrpySA2P89XkpFxZH1iQr2DF1vPiul4AD48ya+JLdYP+WKBAVpJYCdRrCcEnyI9VNAi/S0jls/ecQ/ICoEXGHn01dWu6Is3kOsHhIYJeu3AZHXfw3PWgrajo2WiiIp5ibGrFop2flz50QukvTx2Sg0AdIp/1fQiQs190nTtkbHaq2OLW9s2f/5V39tq1u71sX6QV4iYf+MGBu4Z9hvI5gYr0cAVCAq4vXzPSnwRGA5Get73kBRrD0zadQlkEwplveH8X7M/a8Itsc5mjx74/vGz+B3kvPj5H6SfG1ynr0O9OzPiWDxEokKPaOU2fnFRfvh975jo0MVq+3s2Nbmhr6PT3k2JJ4be3tSIdYOG/LWJRilySKe5Uf5Ybv+vR/a8MSs3fripv3kr/7CmvVNO0pRwRD3tsRAhItXVYMjobJ+8v1nQPLEYD0ChgrMUViFJr79uRXmI0SF3iNUAsYxjGcWyU23jSVCsDOIPRgc2e9bHPi8ON6jIo73SZA+Bv/x2ca51SczsFYL64eEIoLuUsFRil4/7M+p+BrtW8WCys19bML5FayffFxYww4Ia8aFpNWB/mDBEACJ+HMfP++BlQS2+Vwf40EfE33uCfufuGcl52Ycj9D+L1yL27XJxlI9dzwZf93XN0ifZK+PExUV8ZodHM4IePF+A04O6EwLc0Pb2Amrpf6zIxEPZ12slhisr0GSGO+Tz+X3FFsmvpJEhaLP4Gcd98I4hn0AO1xPf8zCHhrX7Mnx1keF6g/+KiImm5VaWPfrv9Dfi+MZEqtKXAE8qNpL7ifEDEF/0ycq9CyC3aGszoLiOD4j7jdWVPi9ubBGQAQq0NDz7XVr5OSz78caXvvgYGz4pWgvoR4VpZzNVAteTRH2Kwk6IP/SWKGM2mGzbZ9+ddPqoSeaS5J6ZmnWhzeMXLxwRdfJ/kX8JIV0omdVJE+SRIX24m5XveOSP9fvhOaRx55l3HsiUaEpmLN8rqS+EUcd+uMRL3vOwRio2hlCIpNXTHVxaF7x9o0bN92itoeKtGEXLlyw6YkpWT+pqnloSEAvtiaAVLdu3bG3r79t+VLJlpae28rqmo2MjNjuzq6dA1SeHFXMgZBkHMLj1l0RB1gF/eIX/5f6V3z3O+/ZmTMztr+3rfevHzZt6dkLjRUVi8SaxBs72/s2MgZQ0bHaIYpIX+fkQ27ngDLX4xLlNiE/gLwkd1ldWRbgw/yanp6SxRQWPYA1VIZQGbm2thGa2rbt3NmzUqCfnZ+yseGSPX/yyM6cPWO3bt+zXGXYxqfn7eNffWrlSlVWG4DRAHWo//H8RsVbyHrPM3o5sKs263t27fKiiIpytWS/98PvWxPL1P2aPbp3TwRAdbQqANP7uXlVMHkEuWINIDyVsgf3HmgP9gbxRzY5MSmwe+70KTVqVdNV9unukX3yyafqT8GcHK6Oas5vbG9avd22biptleExNVJOZYpSXx82yUGIS5krbhMmG9dARiMao2ku4CN1//jSjwwP6R5RRh82W7a6vm3ZQslqKMmLJcukqcYoWhsL1uDHDmBK7gaQ6hZ9YsdtenLKirmsiIpSPi9rYtZ57WDPLl88byPVYQd/SxX79adfijAEvELcNjczYw8fPrSR8XHNY9YJMR0qatmlZLI2NT2lvJmPA7zCPpiqcM7Gn//il7Izwh0AEotrx1qWnJVej/KWD/GYmlTngmCBWC6ft431da2joeEhEVX0c3EbV8iIhu3TBD4IGpirzMV4vkSS2YF2rIg85ov9CsgjlPdL0EDPM+/5x/2x92IdBDAKKK78mJyv17WRoZINl/J27vScLZyaVG61cGbOSoDBek3Gvr73yB4trVgXRXts8hbOf6oY1HRXhIMLjWIOGq3kGGdhEJwX9C0JMQBAKns1MS15NHMZwFg9/mKeGGx9dKbEeIJ9TnEutsgu3hJOobwg9NKUPZbv433w5fXH/Te/Gywd6UXBy9XLIPj/03/l0rkZ+6/+iz+3jRePbHN52axLpUHG1rZ27cXqGn5Jtry2a6lsykZGx4TLAPwCjCOSwIJna2ff45vQvxFyhpiB5+0YTlrg8draqojYw3ozYEU8cxcugMWQa5KHyD48EBcISOjjdnZuwkaKWTs7M27lQt7W1rfs4bNl20fwny9ZDwtsAH+qTto0lj5QJQWiK4BngfB8luQ22HBxfmFnG/IYS+s6B/3nnNiPcUHsCeb9kzJ2FKww3SXDK6OVPwWyjfcRjhJ6MsnpYLhi7ZZXsMpJBDwJ5oRqfCqNMmbXri7Y229dVK6ZaiCk9R6h7V7Klp6/skdLz1UdSBUXVSSqZFQuhGMI/aNMlXT0pAF8HxmpCv2QcDdX0JnMeQHgzxqWHXawW4vVIXESRaGw8jAReW53hDBS/WtU9RRdDxBl9axd79rvfeeqvf/WG/bpxx+r2m3+9Bn77PO7Om9OnT2tvRIciPsijuX6qJBTxX3oYRit4TTrQwzO2nBxiFcWcSZyRn754/n+vH/vj16KtMYCa2//wO3LVOHKugXn8MbzwspijzW5D4BHOgHB+6snBnMF4aaanvvPVJkQ9ivleSfySL8Qr6jntRcvXJTFVuugZsPFrF2/fNbKWbONNfbMYWFMIGh3Hzy3yflTlikW7d7jJyJ1KHra392XKEnCZPI5CDZZTzkOKmyJGED4hm8ZEMrsY7E6SPZxad+vokPFt0TF77qBfvt7/2hGYEbNbsLCDlfNYSAQv90KXp9pqXrkhd9oym819mWInrtszgQsXkrp4BubIQqkapVGxUE5QbljoymFCQeKVz4AvGJD4Qm+VH00ae12DI9RL1N1oCsmPbEppJT2wQLCy/cy8gYkqBcB0OlINXLI4daoS8WOz2u5iI9sS4EHpdqoOShx9ubXJW9UlDIxwgTPKFVQ+ajZcvDI5WDnkKCsjI2C4FdJqPoglMQUe9MlZ7K5p+iPSBAZmxmzq/L+jB/gHN6wGkMUA6EROZUiaoSoADun8i+UQwQGvP/w8JBZu2kzY8P2xsUzlku1bbSS1yELQcCmnsnh3V2wkeqoHakhb8mev9ywOw+e2vDouPyEhysFGy7nbHZqxCqlvNUPDnyzbDXtcO9AJfJsqutbO5Yrla1BwrB/YNsHB2o6l8vQIMrV9dx7n9sxOQAAIABJREFUoYwaYk//Bvzlv7nzF44RFfGZEhBFMiImsRH8jKRYnFcR5IpggpQAzAMpZV19i7qNAIfqid9GVIyMj8n/j/eEGEsSFbGiIoL0CsxDM7WoEopzUcdYUGkc7G3aJhUvhwCOA6IiFjvTmBDSi7ntIHBK9lqA/JT0OgHhinDuxalEwPa0Dn6CPSopBNyGnh4H6tHRU4JMKXghXwoHeN4yNAEMzRG5/ggka25KeRTeS5ZOvga9VPpIXqCRSEgCxirPlj8+KiRUCgE4dexSrwMwBBC7f/+Jra5seOk+Ys3gHxqfX1KReXLz/PdBVHhkQnEE6lJvqMW+oSbAqFf7wBTr1YMX+rvMzc9adWxY3q9ff33Hei0P0glW/n0SFRGgi39SURHHJI7HgKzoCRi/cn7RrpxbsF67bo1mTcHRudNnrURPm5arzWNDTHfGIcihWSwKnZTt11vWy+XtF59/bj/95a/UwM7JFJ+TaqHhsdk3iIoIbgpQyXtzryRRoZ4jr6moSIJTSSICAscBTwfvtAB+R6Kiv+5i4+LXBJjJoNNvyolAJTXxNgMwmZx/8SxzAscbBnt/EjzqezY3O2vXLl+y+ZlpWYWsraxIeQrwQdLE71ORREmvyG+pJMu2vrmpJGvm3FW7/O6HtnPQsl/+/c/t0ddfmvUO7Cjt9osOZH7TMkj7yDGiYgB6xsKKSOrENat9K+xdDioOemBgHaLS/YTlGA9eFgNBhdVq1LQ24nrsEwwniQoStXDtnHtx7H8TCBvP9eRz8HvzigrNq36S6GQoPt7379weVFRIxemAO0AbXsE+ejyugSUO55ArlLzSJ3lNLjhwQUGSVBvM2UAEhdfFuUGcoWlBfhxA/Dgn4+/ECrIkoB7fV71uvL2rQDWAJchdRiAmMK8LKPvvnZi/fdKW8QpxEffDdcX9xJuJ8u9QgSOyJlRCcP2aSoNeRBrHMAclVAykweuIiqgC5TUC50M1ZNJmIP4svu8/lKhIXk98hq8dn7C0nWRyu0bOdz+jA0GfIJQi2KYmkGFfiGssOTdPEhWxLwTPLxhDKQaUnaGAgADWHdtffC5F28DYP+u15PSJmzuWQIeKitcRFUPFnM1PDlkBwA37DZHxPesw97MZGxqdtKcvlu3ps1fWkPiIUDHQLWHzB/x8572PZMNARYUn+xAVx63TonChr2YM8boU+aGiLlZB/C5EhduoZmXlRE+1XudQYBNndrSy4P3Uyw6iIl+wc5UZy+fL9uUXXyo2ppE1oMQHH35gxVzBPv/0U1tcPCciAdsG7w3XtV/+8mN75533JGh5uvRM9k/E2ZACV65cEhE/OTHmfeeyebvx5deKg2m4/eWXn4v4PH/+tH304dt2sLcnkJjYn0qQBnZHAGX5goiRyckZEdSsB0QlZ8+dlco/9vMgR0CoNDIyZs+fPbOVlVWbmZmxZ8+e2dWrV6xR9x5qADunz5yRmOvCpUsag88/+1yAKE25yYWImS8sLtrqyyV74/J5Gx8p28tnT+Wt/eWNWzY6NaN+aPcePLaZ2XnZvwJUb+/u2ujYqGI68gz2/3y2YIVsTnZi9YMde+eda7b0+K4qKr7/B79v6Vze6hubdvvGDbdF6rR1fcRWxLrMF+IOLGUAGolLHj96YpXykARS+HIDVm+sr9qZBZqde84IOcTE3NjYDntkRkp/9qftvW1rtNsiFehNcefeY7NU3qpjY9YK+7tgpSNItkP1vJCtK30C6J2XTsmKpoAQhTywkFfMi/86pM3qxpZZtiDAli+uqVzMyiqKnnEooplf/FTe6PStazdl/0VsDnA6VC7aO9ev28uXL7XWc7mUXVxctMnJcXu6tGSZfNE+/vUXdvHqm3b33j3b2t61D99/154+fapnwRiSL/P6xfOLIlawYF5cXFT/Oip7OJNlh5wrqP/HJ59+arl8UUTI6Aj9VSqq1NnnujLeMBoFPEQQg0GuyqrHoaBcqtjL5VfKMehJsbK8bCOjow5MF7GGztvzFy+17sj1uW9ZP/dcSCjhYlAnM2YQ7iGE7PfeGVQAeHzBecSf6idZP5R6nG0IS2Wq1iCGRqtDlrWOXTx7yqYnhuzV0mN75/o1K2F3xd6VztuXt+/bgycvzXJFrQe+uG4AVQmyyEVCfy4qStiXyNtlH40ACDU1Z26oImafJXcEvFU1NMQXIjaJ4rxyn2unqsttxSCU3GaHWIQzhPiHtci/wQ70Oj8A+62ehYy41+DrjrHXfs9PbpUDqq+CYnSdM8T8KTWiv3huwv6bf/Gf2urTe3bnq69td6Ohyp2RyUk7df683X302O4/fGJl/PMZZ4k2ewKI6ddDv5rdvZoqR2KfKMaA+cL6BgeBaKUSSc8gk9Ye4uJQYk0qsV2Ix5+MEa4TkahQQ3MshTJHNj0yZONDBVW+QY48frFmrXTeLFcSqU6FRFbv544TEFp7YBuydvLm3OqjF6p51A9BhArNwzlLBip5/7vHz5y3cskQZtBVlUSuhNWfu4RAAjH/iO3BkGTLpQeIlTh9XeoitbHlZpyckOsqN6C/2vzMhESLpWLGKqWMzc1M2vhQ2aarVWs3W3KmqI5P2quVDbt176H6hvD5tXpbNrF7B4dqvo6tMuuejyZWwD4K0SNnELgV4DX7NFVoiFf3dna1f0Ju8uWEhON8EBLCxiA9RTIGFDxYYvVkYUU8C3nQUXVOLtNVVeZ33rtk7731hv2bv/qJZdI9u3LtDfv4ky+t1mhbcahq+UrVDhpgclpxssFkTKjsF5bQDvbpAd/wChW/vmj37r1vvHr1i7+b68//7/4ZVZ+QXnl7tbyssWc/4n2plGLOFUoF7ZesQchZNW7HRk3WVE62RhcM8EwnoNzeO1o/JfPYbyw+xUXeL2VxYdHWV5Ztd3PbFk9NyMJsf3vD9na3RdKQ3yEA2NzcU7XJQatpj1+8sKERztaubOAgmBgTz72ozuvJstst9EPP4H4Vsecn8ctdV/Ky//M9y3/yLVHxO2+j3/7iP5YRmGh1+gGEN7ajDLOjgM67yjvhoM2y3RZRwaJwxRR2Nl7iyQJi0SnIHh3RAc5GAjBQbxBcN/tNM9kgCHT4HS37bldBD1YrbEJsLKvra1IDsy7dk9ZVOYCtUjpwIIRAAPCbDYvDhN9H9USiQCICIw47TBmeBxaAsN54uTpctbGxcTHUBHyUhyoBwx4mX1CJGaXX3C8VFWogaKbEIgLaCs6a3lQZEiSq1NnIaEQXdw8RKpTzQcqwKaOUUsMiDgW8Dgl4fRPa2t6SRyAbF6y7SsNyeSsV8yqNZlPlcymNm5iY1KaNGks8a7ths2Nlu7h42ip5ynsprU67ryQNvwI7m8kWrTo2KUXF7kHDXrxaU0C6t71p2XRXByx1HsVCTmQF++jU+IQ9e/5C5bJstuvbO9ZEKaKgIKMSRkrt8Rrm2aAYo6oE4EPenVlPNGcXz2vMuD8HefzgZE4RCCbBhwgYnSQqIggSfzc2So9EBX/u72zr/UhAaZj9myoqRsfHdO989ZtpB6VMbKZ9kqiI6m0Hg91ah/8ECqVStrW+bLsba9bBnozDg2QHyxEx9QMSwhdAT6ol+gowRmmIitDAOPpOY/Qk/8RMVs+SOe2BlFc76aBN9bQ+ll+uaE5gueQ9KnKWLXiPimgp4c3qXVdKMJEkKiIZxFyVV6oIBwd6tOYCQcJr82lvpO0JR6QjvfmW21JkbG/vwO7cvq/m7ekUgQvJgAOF8eB18icG6seB2QFRESyXHMH1BOi3VFQkQUM9zgzN5VKWB5SVyqmnNS8xP0lbAK7ZM3hGKApRC40TbDbbdufWfUsf+XztExW65BOVFIkeFb+toiKCpnEMkvcSm2lHUmwAlprAgsvnztnC3JxNjVU1r+qNA2t3GjY5MmHzUzPuCRo8ShW8BExS5fCakRnbB8jB7/rw0P76xz+xR89fOlGhMlOIihAUnSAq4pqMQHi+4E29Ikga1aBOJnr1S7Kiwu/Fqyb6ZESiR4WAOF8k/eecJMiOPdcAosakI1YAvO78jeRm8mfJwO8kKBnnl74fCJw+USGyKiQ7BNqsLfkRp+3sqVN29fJlm5+dtf3dHeu2mwqkUYEBCG5sbctSDjD90lsf2n/8X/4Lu3n3kf0v/8P/bKtPHlr6qGZHafr6BDDzhDpf1xWsgvRs/wEVFXHstGdJjcN56h7nGp8Y7MYGmOGsJzFt1g+0ByXHPz4rWSwEFZMUZaG60ZXj/qavIyrinE8C+IN9gWSvo7Naz1cVOm0ppP/5n/+5/ff/8l+qxP04sZBSIt0La3BAVARPbAHQDjJEa7EIDpNMQZQBXEBwA2TFPXLwuz5OcQ1EEDYSFVFVnpw7mj+q4ji+byWJijgnXbmJGAEbyYxsMGJccHJO/0OIiriP6F5VeePVIf5oXN2qZ8Wai1xhqOjSOg/PUcMX4kQsSJRkhQuLjbTjs+bP2MOir7QNv5usqFD1YIjniL36REDSEug3VHjE8/+bRKQrOrU7B9shfoc4SfEGDU8DqRT3hZjAxiqOOL7HiAEAqERFhe497A2qEJOKcbDnIT7p7zt9ICqIDtQfJvShCURSnIu/ac0kxzbuA3oeYVyjRR9NKivFrJ2ZrlqGsW02rVJ2H+dOr225UslqnZQaBmODAsCkOR6s7XqqbPAKzDffed9Gx8YHREXs1ZEg7CIRFJ9r3O9PEhW+7wzmU/9cO1FRoaa0qZwVCxX1eoCoiBUV5CfEK3wGcXA251YdM7lRKxWH7Muvbtj4xKQsTre3ttQQnNj1s1//ysbHxyW6mpmeFhiMLc5nn31u16+/Y6VKRX0kdrE7xZq1XrMLFxat12vZ+MSora9BGszZo/uPbKRatcnJCfvxT/7OKpW8/bM/+L7Nz03JLsoV7ju2tgqwgtqxoFgD4FhqScav1xNwOTs7Y8vLK6EfxaFU7AifyAkkUJFyHdVsS8IWB0G84fHixQv21Vdf2+/94Pvypv/0k88EWC2/WpENIDnHpQvn7emDe/a9j977v9l772fJ0+u873TON+fJMzuzM5uwCYsgQCIoUyZpkZKqJKvssv2Dy1XyD/6TXJZl+xcFixRpipAAggSwADdgsdg0GybP3JxT9+1wu9v1ec77dn/v3VkEKhWkucDW3Nj9/b7fN5xznuc8j507M20rS49UIP34k1t26eoNQ1nlvQ9u6r6Yi5xRdKewton1pNHfcfmTPMUwulm7LXvtleft1q2PbP7Cgl179hlLH3dsa3XdNlZWBNSfWVhQ8VNSMdL0Jn8hbk3ZPqz+dMZu3bypIiOHDjkbBXX28+kpOgkyKqhTSD9udwUg0ZkCe5ocY2YOwKfhoI+kUvq2srotoII1yDYFi157b9qLcZB32INhIpN/0FEBeY2zAPNTVAQo/PDQtrZ3bXe/btlCWWAIxfP5mWkBD/1eW7kjZzoyHHRI8jyQj61VqrZ/sCfmL90AgBrPPfOMCruSFmm3bHJizBa4/lbTJmYX7PUf/qVNzc3b4eGRSGp0/aysLCtHpqMfUArpJ3Ipxa3HxzY3N2f3790LslppScfOL5xRnPqTn74bPDn68mFgrZBrkh+TQ1PY5nUYYyRYmF+wlCENSko4lbaDwwPvykAOqOPd7BTtDw4bAtjimUu+r/w3kA5jHsEc9d/xTgGdtyoYOyAfzwbyHl4bLXwM6jEIT+fJBR2ExPQbAGl0pGK1Ys7Oz0/Z7NSIdY8O5cE4gn8M9YdUzt5890O7dX/J+lk6Kr2ASQ2Bt+M8p1NGpz+5togPDgrGPRfQyX0qXC2CIj1zhIIn8S0eJFH2Ll4/98e98nw5N1QwJ68PhAdJ68D4N1NXrcht2sRD17DkYAeakwLR4r4OOVGd5/x6+Dz+cHA2xY74KMlJ17QknM2unJuyv/Pbf8Mau2vq9t1YObDN3UN7uLZjlcmK5F539g6tWATIIv91hYejdluyOhiS0/HD/R3W69qb+D4DCohULpZVVwGwkIlzgy4mlwNlTvBcycMFZlBQPvbP1cXEGu0dW6WQsZkxSJZNm6xV7OKF8/Zoad0+u79iVqhYOwVpQHRPgQaK5/DL6B7bzv6BxlZqFZ1jARWoEqjDEJAidH5IJDnEbK4eEIyR1WURJScDAU1SkwDfeSlKqFsF4Kx7LBDATcRrek+6Kng2AFF8ItALUG10RDJMrWZDPg6FXNqmp8bscH9H3dZ4GIxXKwJJ2UNyxZIdNtrqbmTM6bA4bLYUw1KHcv+H0AUcJMEgVkY5IKYGah6xI5Y9CY8fAYCDTgInF7A+Y0zk7HyvQfkUdG8YpLI0Xki99js2NlazbKpvzcOWfe2Vs/biM0/bD777utbn3Pw5+/Gb79tuo2dTc5PWy+atddy3UnXEPVhaeJ+6qghbsaTaw9rws99BPxHoAlmHvUqS7Om0/ezP5gZh75f/1qZeB5mk7a1t29rZ0WtK6g9AkK4p+R06aUm1k9AJRt7rHR2uxhLjFPZE9oNYT4r1nNPkqZioShWDeVupCqSlvoNqxuVzszY9WrXt9TWBwJVqTRJr7JeIfFy78bQ1ux27de+BamdHRy0ZjnNeROIz109MQDcZBOTo6RXHKJIPGC8BxVJ4KSoukIJJlK7Kzr02hDMelwk/+d6TEfg1G4FZ6Qq4BiJFZJdNIknwpJWDxlkBzowUezq4y7tGmgMHsT3JzWg9ASPoQ+8SZJ2DKhYlPAnxgYp+D3zp5kCu/6hOjRQmwW0ZUIsJRutrNMEMLXFiz5NcpVM6LFnMBFwKHDg8st6C7qauzsxcmJ+1SqVs46PjkonQBh4104WIewsabBKuX8FGNqtANxbE4oamQySwPRUUheIpmw0GXTLGDW2ZMBYiq5HNJpqQkYCBsHqNsCcWEbIzJCoAPE9ff1p6eG/85Y/dEwTz5HbbLl64IG3dt97+iQ6q3e0tBXMjpay98qVnrF1Hpsk7Y9j0CRIwPGM8VaSCJVUdtbWtA3v4cMl29w6kVF7KZWTQC/rfqqOD6qVYxgLASkxK9NOzOcsWK3bn7n35LnQ4OTFt6nRsYxv2vFm7C6utLfCCrhGe+8zFSwr84ljEwjhfJ4GKZEGIOaGxRn85yCTEjgYvmLqxWJR+orh1AqiQ9JMbyRJoEADwTAnMxibHBK7xAbgmabPAZI5ARSwcxI4KDsT4/rE4Fa+XubyztWoHO1vWAqwbFH2HYjcDM09CL64BM+1gZk/xXIl/MGjnutwwi6DKdfG9eARQ4Qezij0svTRJRsMeLT6yev1ILCKCSjfHC6baIcHXa9Dmms8FQ8ahrId3OWUl+yRmEOsx4S/gfjIm7xIZp8GaDKwAnrUbwcLsR4v4jm1t7sAXlpyD1j1sjeCBwAJxsMfZFaeLMZH568/Ag9b4Ie36sP6ijFJcgzEB8WKWCD9K2EiaMZSjxZeuD4KiXquuee5tr5iUw2xG8iBrI+hIHtbt3p37Rg+JV6aYIg46DfXeXSt1WIH3AmX4Zd3voKjMXirGeCKkYO8NcmYk+bE4H9eJF7x6Njc5Yk9dvGgzY6NKngsAku2GEtFuq2NnFs5qv2UtsQd7a7MzNiKzOpXOSe4N9sthu2kffnbHfvD2T9S+TJFD1xqKucmOChVkA9s4FpkKxayCJk+efM+N8mwEwf48kywm5nZG9++378CUAwUBpDoFVEQQIc778KKfmysOKjwmTDslFTOYP4nf9ffwa0j+fABU6JzU7PXuP3UchESHP6GA2evZ5Nio/a2/+V8JsHj04L7t7GwN2P5rG1tirDIZb9x41h5t7NirX/u6vf/RJ/azt9+x4yZScYC43mUVg3m/Lb8v7TNhDThoFrsWTspmDQvhQdonoSEfjSPV8RD2RS9AD71R4nkdAcrm0YF1YBQOCtihaM11sjeoIQNWG4MRruUxHSGxOO6HZehq0a35/flt+mnY7bpuMl9GIPO5556z//F/+J/s9dffsD/8w38pdqzvJxRZUkEOhoRo8AaSBuCcVgKScja4YFQYdUhK5iiMOJNLrDS6RiUdhFmxI2qSFggdKS4jEC42+HNpD1bBORaiw/tr2nih5sT8Ck1DSV8dMfVESvCuTu//GHpGnAbWBl8HMC1KWrEveteIAySDda89dghUOEAxXIO6dkkgJDt5/He09iiDiJUH6AY46Sw1uV4Q5xXyNlIbUwH49qef6tl0MUQNMVV8sjpLkp1CUb4vdJFqxENXh0LUsHfFdXkamEgW9uN7KJaVEakX3MWuBagIrEQn5njsQGJLLOpgixNoTgOX8esBUOsr1H8v7H3O4vR9PZ6vcexPMGbjNiWQwU1IGccBYBQOwniNwx1p+JlvBnEN+sgQy/KnJOawjc9NV2TmmTo+lmcObFm6KbKlst28+9AasB+Pgy9I2NPY1zDyjVIJ82fO2tlz5514JA3uoea8gK2glay1EQpwUdLzBFCBXnkwGk/OLx9zBzp5Ma7fz+y0FYtl29zYsk6bONxNZAHHvPiaUTKfyznBaaE8Zbls0d57/wN1ADAniRuvX79u5ULRbn32qRioMzMzdunCRXv//Q/USfvuuz/TXhyBCuJgzv5ms25nzszbyAiEqa6KyHRSCKgYHZWfwU/ffUdFgm9+4yv21LVLtre5KdIJbMkH9x8pvioVK9L2p0hzsN9QIZ37oyjB9VerNV3nvbv3xHxn7UCYqdZqMielsL6ysmJXrz4ljwNABMZvdm7OlldX7enr1wWG/PTdn6mLFpNm+Qkc92xydMQ21laUD0xN1Gx3Z0tgxoPFFZuanbfWcco+/PgzO7NwRvOes2l8ckLXxnjTicCaJ+8YqVQJkASAPfP0JVtevmeV0Yq98MpLehZrDx7a2tKy5ILVoYzZefAsIN7qtrwAdpzqi8RFR0Xj8EhFHYqM46N0evdkwo2cVqmcl0wURK2tjc0gowspo2nPPP+MlUeqcvARCHREYbkh772Dg4Zt7WzZNh0HFbrkvZjF1+yLdNhzpuATgYQPa+7gYFd5IV2QAMUbm5zThwI56IY5opA+VrNWA5+Lqp4nnfjkCns7u1auVLVnk3sC6lD8Ik+jkIREGMUrfrcgyZBLmjsQ6aqj4/adP/u+zZ87b+sbW+qaR07y4aOHKqIDrKmrhVg1dPLzOphxI/HiW7dLQ0HGQmrtw48+FqhA4Z2OFZ434Mn42Kj+jk4Mum8bR3Xb291X9xBeFnhzCPjL5pQrqlgLwCHp16xtbW2LqMiYAvgSS3My6eehG551DOgQ6wR00egkD3Egrxd3sLifRmCXswMwYAUZoWJRUmBLS4uWT7sR9Gglb1cvnZWE2dH+lk1PjFi1wpi3LZUr2dvvfmQPVzft2PCF8BqGS9x4PgfLmX2W3JDu79i9L/+EHN0WgeQQOyoDAMy4aF/2EE/Plf2B3NH9LR2c9piAnMD3TtUR6GLj+3gzNJHOdLBE+VHw/vS4IPiKBaZIlDSOJ3/suAwntUtCxu0/dAZo9wz+I/1Oy5556oz9/m//hu0s37PVR4vWaaacrY8ZeD5ni2sbtrG1KyleOmkA9ukoKGGejTRWp2sbG5vKD7luCsTERQ4WUEvh70rqcmBskT/j7+TLGWIlFh8FXTxhAALdX4caRkaSXZViWt0U45L2yll9v2GpbFFARbpcs2aPWJexgj3u3TPKa8oV26crCNkcvBWIu+S3FnwJJXUbZXp91JKkhijtMwAwQo1LHQgpr2lBkiECyyPtJO+ahtY862Nmdt52dves3jiSXwY5NutUcmZB7vbyxQtWq1Zsb2dHhFFySfLLfrdjtWpJ6xsgEElFJPswCm/SzdU+lqcJn08hY9doDGS9AHPd58TzKoEyIg7QrdDRdbB3U8inThLlgBzsZt77WMT6BfNe9Ss/dAUY9OmoUKeB5yH/8L/9fRsbydve+pJN1Epm7YZ9/N4tndkjY9P2sw8/sUbHrDI+bd1MwTqQzlQ/RFq7K/IuazSSFwZy3fLGQRYc0q4DhCKPBFl5rv/NP3UCKR9f/Z0d3R9qJJCJ2N8O6g3VzqIRPbm7x5Yeag9ymzBnibFiPCzSpbZPz7vJYaMM3MnYbxgja1b1u9qfeH2Ap26zZdevXLRMv6uak8BGybmn1ZlXhpSdTVur27Wdw7qeM/vD3vau5qxLbjlJjFiX7lX+jnyEZ0s+ILlH9k49a4/n3RwdonRT+wxnjWoGT4CKwZx58sl/JiMw0WJjjklOZ5BosGlJI1VF/KHpa9S2EworfVHvplDykIYF40xA193FvIZkOepBw3CoqLjDRqODgxbPgssciI0A4qqgwDdTN7U2tdrKFBjEV6wIL3QqgJCuvzPo2HRV5A0MQDRHYakTKBJ8oU17ZmFeTBptirAnOt51waFBgZaNwAEI9F7XZfRDYUlSN2Kl5xR8KEAiuEFGKhTelaSmXPNRJtu0R+Zoz0L7FIQ6Goq7kREfGlO173qLGtcr9k//WF0aKqD0zUZHa/biSy/ZD7//AzFeCJz/2je+ae/+7H0FkdubmzYxUrXJ0bI9ffmCpKAw1iUYx2yQA4KgQQecAp20VUbG7Dt//iOZuhGwwATKp1O2MDNtI+Wc9dtHCjCQv6rUKtKY5GApVapWP2rZ/kHDytUR29k7cNZI68jypaIOvNZxW2MgU6tM2vYP3QBq9vLlALhEbXXvrOCDcT8ZUPghwvcJiBlfzQu1LnrhyQsBDlQAskm657hjh3u77lFRKtvo+HgoSmRkdqhWSdrjux0bnRpVVw31BtomAX1cgsbEpEoW/Ly7x2V5kj4skfUfi+LoubdbDbW6AzwxP47VveTXh04IBQFY6+lu16bGRy2HKVUBD5akQfxJCQ6CQhLBWMBgnvthSyKclvQEgc761qatrm14K2G55F0VQTc7mlr637iRJ+BILNJw3+p4Ivlg/Ua9RxXWhoFALBp3AM9UEAoseIo10qkv2vLyqhJwFb4HBTIv+gzZAAAgAElEQVSXXvEWSy8axgJgDCiHIINrRfp7RRb+sBDNMxgCpycL1BFU1BqT6TgdJznLl6v21I1nbf78RWv3emJmbC0/sMbhvvXQhyb4RRM1gDPpYt4O9/dsc23D0k5l9+RLxTOX3vKPCFREBXTtauFnXvzHeEwa8QQcHoJ7YKOK6PD62Q+SwVIcD+Y4Cdsz156ymclxOzs7bbVyyTIYjPe6tr9fV8FlemJK3Vd65hSoB8XklDpoRDlKp6zebKs48Wh13b73xttWr+MpQVEvdkM4wOsgRMJIOcw59l2YeeqYCz9XYRDZkwG4Fg/LkLzJKB6gwl8vPt8TR+rPASoGRUkR04bGjHoCiXWZfL3HvsepYmRk0STX++l7jq+ZfDZi7wSdeGTe8qm0Xb140c6fPSvZgb2DHe1/FDOQ5cC0EFmH8xcv2mcPHtlvfOtb9r0/+zN79PDRoMlEvrcD7S1/1/ieGlfO1AiYnfb3CNMwec+xWBrnkToLJdeYUeFMUgQwzwUkxkJ7fD7uO4O8GMnaAJhVAul7T7w238eHkjYRbIkgp9/JkAEuMCTo6J7UhWWdHVurU/dzNrwq6wRG9Ne+/g1bOHvJ/viP/sge3L+tLglauHk99jMVyGLHS3gPAZoyYPTOSPZeaSxXKopbyqWC5vph49AODxvWOEIHmXVOEdXXuVh9AbhwX4rgT8F7JYDA00XugTzQY+Y753zygzFEesMBKXcNiDtDsisjzgklJ2HvkMyVusy8bT85ZwYFc8mhRGadt7/HuULxCbmWuKPpGtS5GqQBAW9gTB5jBgwBIqP2dv6jaDk1M2VTk/NWrYzYH/zTf2b1/S0yOTc0DSCY9s1o2j4AdXz/03ojETsNVCS+PjFYp76Ie0McM16PeyJZhslJfKPfCYbz8b6S6+v0XnEaoHjc+yf3ibge4p7AHpUkM5ze51SEUqHeYw4/2wPwx7wTgOBPJLnW4usM9sPQ6cDX6lrOp+zMVMEMJnW/r+I6Jp3FkTEr1Ebs0eae4nOKqxQFGKP4DPByZEoRozprr+wFkxBvKfZKdFd+bn8J+zIdyXzEjgudRYH1OATPhgQJrcsEcEZ3FJ3NR038GyJRitjZzbnFOswUVCg7V50VjfbO3bsiRRBmMUefeeaGlQslu3/ntuR/AC0p+q+urYkZT0fFlStXrVip2P37D2xza9uq1YodHdVtbm7aqtWiOqphDzfqDTvYO5R8FHvRhx++Z5VqyV599Ut2/vwZ29/ZsdEabNKeffbp7WCUXtS/27u7lk7TUeHFGIpcdGdj8kwXxsrqikAOvqYghQQtexlFCl/THRUlFOfig0RnQLtj07OzVqmO2k/feVfElLv37smfjFyihLFt48C++uWXbXZ6zO7euaX4cmt33yZm5i2VKdint++Kzd48ag081KJUK6at5GysIeJO5lKq37ZsqmONxq49/+JzdunaFctnsiqGPrx73y6cO697BKhgDlFY6qcywt4hcO3UD8TMbh21BUJwMxQbeewquqR6NjpWtdnZaVtBPlXdoRCuuioUUhC9cPmCvfK11xTzuCY5/jMdW1ndEkBDRz0F5jv370sCDK8Gin96j07bmgBB1YryK/IyFlm7fWSTY2OKM3k2u3v4TiCr4fnLSLVkM5Nj1mrWbX1zQxKOyjk7gNCcemk7f+6cra2uWb1+YGVev+aywvt7u1pjE+OjNjc96TnVUdPGJqfsz/78hzYxM2eHSLYc7MtIfWV5yeYXFpQHEkOMjIxqvhHrIuH03HPP20cffmgL8wsikJEb0VGxur5m7/7sPe0lnE8QsCisAoBwkiARDOubtQ4TV91KPaRZSsrLWVN4s8jDL8ZSKe/IB6wilyJn4DoAUSDCsGYBaVZXV1RY5XrpukAlQcV42OcyrfVx1F4b5GeS8d/ewZ7Nzy8oPiJnBbTj7EfvH43/kVLOnn36smWtY4VM1y6cmVO3Knr12ULF3v7ZTVvf2bd+tiSdfAEodAkJ2MM3rSiCHQVouqXjdTA2fGgfDFrvXDdSzvyNuvBCfs5JLMDDmNeoFUAAYyyLA5lszfeeEzBc+s8BiyMkygRUDOEHxSjiugw7T3/e+RZ/hv+Ce1d5/CQyJaAQuRRPun1kz1+/bH//937LNhfv2q2PPrS9rYZ1UhnbarTt+ddeUAf14vKaVUo1q5SqqvUgNXQAuRTpb5lQe2zn3k2Y/R6pwC41CMYYmXC6/CVX1FDBmNiUa6L2oi4EnUdp5cAQBhgrchOo5qg+XJibspx17ZUXnrftrR1bXt+2z+6vWmFkQh3fxKYU/1EHp2OZ9Y/U3AHFWxXBvavT4wY/I1QToibgBiAB/Pbzkw/3IvOuykhKkFJH+H0ZLKvD0A9CiJvsKRcunFNX9MjYuG2jKNE+tnrzSPtSs8We01AxnSL6aG3Unn/uWVt8+MiWFpetlMfnJhiokxemUgL9XFK9KSCcucXZxtlIl9nm1qbWqeS4KmWdBeyZDlhArPDrZ9+gu4xaE2cmslLca5QAVhwXJNW4R+bs0GTbB4gx4VqG0k8QhLp2/fp5qxZTVsp07caVczZWztvmypqVSlO2e9CyDz++Y+u7hzYyNW/9fNnadIJn89qveTA8cyY5hXXqMdSz6Bjc3t0WqUnycahFqHPf/TDdUydrP/pjOr7847Xf3hnUCxhfdRW0OYea2gM8bgveEupipobopumDGEnddS5nq72p674/3rXgHh9JEmqMuYb/ujS09oa8+xV1jo7s+pXLlkuZLT96qP0RiKsvoKZvly+e1drYPTwQORCIiXN+e3PbmvhbVCpSRimXi7a5vW17eFUF+SvyavZmJOhZN1wb9xs9R+jsQMre1W+8fvYEqPhldtAnv/NrNQLjR25QrAMvSCmxlasNFp3XFia5XkiMesMsejYbb+v04pC/RsqOgrkzif/xMXprRTEsZLwr6QZPjNR+KwNsZ6WCNjv6SyLjTAj8Izj0o9E2h5DMc/oYORUdFMEAudHQIcEmTVAdCHhC/Xe2Nm1sbNTOnTsrNkm5VLSD/QOV6mFFcE0wqjmIuTaZZPdMrY7c561bt8XyOIIFEFgjbJAy34ZR0u/bzPSMCnVR5oJAkkMDYAWzHJB2GZLLhNARZu6Zw5wuFnWbBHScN2fDbDYbKjDDoILtyUYE0HL58mW7e/euAyMps0tXLtve3oE9fPBQgUG1mLdL5+YV1I3Wyq6viHmajAcxuyLoHVEwOLtwxn74ozcU3OULtLXiMXJktWLJKoW8zU+P2nHz0PJ5fx77uzCH0EPMKplCOqp+1LRHi8tWhDGF9isdIc0jMZByhZx8MfDH2NnbUWEW3duFp64NtEwjyj4EKghoh8XLWAD4RUAFB40fdl5YhV3+RUAFmpwylAao6KEFOWYTkxOaixSoJGchBvjngYooqROLsDHQjoWIQeAN3wU2PcmFDmiYFJ6MsaYO1R7esF67ZfmU2RQJBWyuPPJmtC07UzspqcB8hFFSUudQ1NB09odAh0zK2phNHvszWF3flOE6gRMJbxKoiAwiAAxa/eXVkDAsdWkozMo6zrZIFCPjmvd7xsO9pWIKewaTUq33KcDBvn3wwYe+hmWs5lIzHig62zc+32RxSMF2YH/HwtywqHGC8K61kgQqYkCiED6ArRobwCxShHTaqhOT9trXv2lXn33O+tmcbW5t2fL9O7a1sS5JiCoJ3MqqjJEP9ves2W7Y4c6ONesNS3Vj18MXABV64ygFJb5ZOA9Cu3HamVvMhK5M0xNAhQpS/hE10vW7CckY9uB86tiuXL5gl86etTMzkzY+WrMC8bz1xc4hyaTldmF2TvtELJjJdI5gRm2iPc2JZtCQ/fTeffvB2+/aYQMzPALLaKbm+20cz/i8YuD2RUBFlEM7eRgGoCKFjJiz8aKkzucKcL8CUCGmW7LbIDFe8f3/SkBF6KBI3nN8veQz0eiE98frxDpdm6jV7Mb160ZNrt44sPVNCgJ96T5T3JWx6v6+ioa/+Zu/aX/4L//A9bgTcyD17wmoiPce15T2lQFQkbU+DHpJoKUtw7P/HFDhRIB250iAdbK4m1xvcb9S90GQFoqvFa9h8BxC5f0kUBHMSMMgU1A4ah2q4CYRyiC5w49hG3/jr39L6/973/2uiAexm4C9vVAp++xSZ1Dopgiyjr30sb7H+ZnPpG1ibFTdmMgc8kbEKyQ+O3sNlx3gXuIeG0Hb0FHWD07XAqvCuXUSlPGb+VWACp4T5AeB8SRviUV0GgDxAubngQr5QXVhkgZmfyiWx26BbtcLEPFZ+vnhRqdJoML3/QRYTFHRYFs2RUSokoy/+JKNjs1YOpdWrFTM1yyXK9q/+uf/wlYe3VGHkHdnhSLBKaDC97jQYhCSVRXnkx0VfwWgwp8JILUDFY1DdNnDfnwKqEjuP6f3iuQefHr8474Y/42F/Phc4r7gnTYOWCT3pDivBlagofMtxpIxlhXQHIosnwPBHuNhw3vks32bnygAO1sulRIjvpvO2NjsnBVHxu0I1feOA/2sLxVdVfilyOedilxz1LGmYBc9avhZ/Ll3XjjYMAC0EkAFTyHG/zGeiTFE8vfjfSWBF4o0W1ubYn/DliQuitJP3k3hQAX5wFS6ZqVyzT54/0MxnwGGDw4OVSyiMPDWG2/YtWtXlTdcvnzJHjx8IFNkZJAuXLwoCZQHDx/KvBsQoF7ftwvnz9roOMQQJ0tNT07Zxx99rNe4dOmCvfHGj+zCpTN25sysXTh71j338kW973s/e1/XdubMWRE+6Fy5e+++PX3juq2tb9jDh4t24/oNu//wgSSg6FiZGJ+0re0t3df42LgTtLIZ5SOwc3vHHckGIuOK79rtO7ft9/7O35UJ+Ec3b1q1UrPV1Q39S5EXXwW82l545rrM1d988w0rIznS6dnY5KztHtTt0aMlGXIf7B+K0JIvFUTQcVNvcrojyT7ByD9uHlkpl7KF+Un75Ob79sKrL9rZKxftw5++q26KF559TibPjL1ytRRdFYAmfSvkCopN3rv5oTo6ACeId/M5CpcN5ZSVUkEFdUCKq1evaA+jOEiMCqBBt3ZpdNR219dsb39XcTvgR7FSs431bXvvZx9auVy1UqGsAjOFH/YWOowp+DDfyH/IpQ4PDuT/QYEwnaGIX9Ec4whf39i0nd19dd6SyxRzLj+ELvv4SE3XA9gCuetw/0DgF2uU50+HDKAV3Q1Iyo6Nj6oQyfmOx8iNp6/J2woQb2Jqxv7FH/yRXbt+w9bWN21vf8+effYZu3v7tk3PzEhGhsLjwd6+OvTJWbkHwDAMjF0a+FB5cLU2ovtdXlnWmHKmc89u0MrnsSDo3mUAOHTvIIG2sbkrDwDWNDJgB+yVrP9AZJK5erFkzaYTxrwzyrvHImGQOUt+WcgXbGx83DY3Nj3Oi8XidMpZ3iE2FwM8AHGVSklnupQFJKWZU+xdLpZUTCzSrYec0fl5m5satbXFezY5WrMZyYTl7dgy9uev/8QerW5YGpKCgBpTvk9HhfIvdjn5/pF3dBUjU5+QPC7KC4HQIC+PwDSncCw1ibD/8lqMP6TCuBfKzJhYutkcdEcBMkr22DAFdh8OuhE4AuN5zozRWChejR1lJyPmL/qKsIM0Q1GH9umsZIDV5U6xuXVkE7Wi/ebXv2zVvInItLm2LS/J5c0ta3KuZ3K2Xz/S2sS3slodkYclRfHNnW07rB+oHsCeLeloqW040EcdA3CCzik+Z25HH1GRx4472jMAAVUrOu6qm219dU3m7ToHrGcT5Zydn52UBFS2h5dm3fqZgt16tGZWqNpBy/NPJIjYyzi/AXwgG27v7iiPIl/nvagPOUM/EFGCtFPSh07+XJIeGhJFOW8kGZtOSa2AOXqMZ2iqb7lMSkz5yfFxKxYpsGe0d7NX09VBMR7D6+roiPYj6hvsWYQZly+et3Nnz9lHH9y0dgv/TNPetLO/Z9kiRtqsBy+cA+SoS6DdEgjOuHGt5PR6DyOPOFJRn1wWwMLZ9B19j64OajNSpICMIyn2vPbXaLQM0YA9V13vuWzwCQ0eqip0O8FBklDMr14bwWm79tSCrT5at26ra3/zmxflE/PG6+/aufPnrVybtFx51Mpjs/adv/hL2zo8UkcFkmHkOKwdvDU4u/ga1QjWIoAFc4p/OeMYV+7V51HaapWaAMa7b10ZLIFLr3yq84N1xk0wT7lWSF+AaoCoACsiG+O1Ihly7+ZnjWoQqaHQHRTIruwDAqrDnhTjtighnIxFPOd1dREUF+Q7227bSKloz1y7alub67axvi4QTYBoJif586tXLlm3f2yf3b2vuQ+JinVDlyCAErkYxKSnr18TCHfrzj2RfakP8pxRQNnZ2xXwxdzmXINYAIgt/xuAl6wTqQGsngAVv9we+uS3fo1GYOKopckv8IEDn6AmaNd7koLJDa2daLw5QhqLNHzPJVW8yAmrIrJSKZ4SCLAZcWiREPmiG3WmtuR1hixRNmoh4LTxHuNn4Bqt7hdBB4O3VDqqCIJfsvWNDX0fBFaMbNqkkJAJhQla3UfHRsRaErIKG0xGxRFY8VbNeJDJDIsE7NgZhAAAy0tLYgXxNUkT9yBNOBgWIMaWknYjAWocF7Wnd9FNbStIF9qv4mvoAqDYmM0HoKanQ8MNyfyAZUzZhMrFgoLoV159WcHfzZsf2t/5e3/X/s23/41M9NCxf+nFl21/d8fu3PrMapWijdNRMVaxidEax7ZYC2jsalzQe4TpENgyUzNz9s57H9phExmHnoJQpIQoKpRzOTGw8tljGcMe7O2poEOHgF9k2g6PmkaK2+2nbRdEG6+NXkeM7cNGXRqy+WJegT4Gjkg/UQSavnRF7Mb43GLBhH+TXQqxeMD3f2mgIsjp0Gr6hUBFtaYNXkBF6KjAPJADvFF36SfXJk8pYYtFWf6NQEXyYIsFiHi9+jfI7IvB1fbAjnVFIORJQl0gUq2Yt72NNTvY2bFyHvAhLUBJQXPoHhFbJjBP0eKEvcYcJKiIHRVe8Oh7yy6HZAqvkz17uLQ4MHcXKIEXCOs6MN6VmJL8JIAK7icavQtMDNJTzo5ycEF7A+wjwKcBUEE3CAXPlPXSKfvk43u2trbuIKaK9xQzXDpJXVaJAngsDsWicBKoiD9TUWMgVeKbbJwXybGP229k9vtrBh4ThcmZOXv163/NLj/9TAAqtm1zdcWWFpfs/LmzNjs1advbWwqaFh8+sO21RdteW1WLZ0ZyMF/cUTG8V82QIOGjGRQkmEL7Jl0bCaBiAFiEi4/dBhEEjgGUZPl6HRsfrdi1y1fEKpueGBWwSFDNXsUexn5UKZasSsGAIE2AssstAVLSwi8mHLILmYx9fPuefefHbw46Kvoyt+YZscd5VTk+m2RB6YuAiliQO1m0PQlUDPR3o1FvEmD4VYCKU2DO44qJfxWgIgmAnH7NuE+Fpzw48emoMLHMUnb54mWbmZ5UUXdjY0MmrXR2kawQcMPeTeeL9syNG/bjH/9YzK2gWO8JrFOpBx/xGgSS/godFXG9ngQqXM9XjD8YXGzyJAtyOjrdURG0ZLtNBclJYkJy3cYuTHFLgym6GNIJLwAnPJz0ahCAmyiIxxvudtvWONpXl6QK/ZKM9PWHTAQmrq+8/Jr983/2L+zenXu+N0mKyKw8guTHsPjN30Zd6r46GFwuACmOibExK7IP4tUjY7pjAX5b23syahVQESRuKC148hJY78EE3osOQ0AvCeZo9QfpLoGGpwrLpzsq+DlFH+YIYxmwkBPxUhyjLwQqSJYfA1TEa4d3GefFif2ScxHSiL+bCjQyCg0sf0xi292O5nSnd2wzc/P2jb/+G5YrVKXBXyiVLJ+BJViw733n39rtm+/TAK+kfyBX8BigwvdNB/zQsma8/mpAhfuq8VIqrKCnnWNvdOlO/TSASuqqSJiGn9zXhgvPSQt+7j3uI+6L/CzK9ek3o05yBFFVyHeJg8EcCNJPrHyt/oTklj5PdB+dWGunLiQ5pzwG71km1bMz0xUrIftoJrnTUm3UxmEtd/vWzVY0j8Uk7FBIR4vbjefbQaYkkhu827Suol+UdeL34/hJSi4wQQfPrecdyR77hhg94RdyGtgYSGoFQIbXIYEHqKAjWuasAaggDiBG8TiFboeCLRQnrN/P2v37jwSUcX7zUkinQmB6/fUf2vPPPae1/8wz1+29998XgHHzo0/s2eee1+vAfF1dWbfqSFUg6cVL58V0RGecol2pULT79+7bxPiYvfjic+oyK5UwMT20MSSf9utWKVWs0zq2O3fuSpYPEg/MW4y1662m2P3EmHQ/wpSnOE23MkWKTD6r8YecNAagAGsbmYidXXV4UuienJ5SoXy/XreHi0v29/7B31dhfX151a5cecrqB4e2vLSicZenUKpnlVLequWycqSNzR27+3DJxiam7bifsgcPHsq0ub6/b/2Mdz2wlnnm2zs7ygsrpZKKV8SoraMDe+VLz9lP337TXnj1JXvq2esqsBErIXvE/KBgVi4jNXVg7XbPyqUaCqcqKO0cbInAhCzRysqazL3HRsf1LCis0fXEfz95+23b3T2wZ595SvdMwaY2MuKgOsU4o7C5r6Ix18y/77//vgAnUlWY1h9/8olNTU15N3mhYHv7+8o7iMkhsBEfEVOZwcw9spnZWYHU6O3v7cNwzmseIQ84OzslvwTOCvI/vBf5e49Bu7a9taXzVFJKwfsAjzNIXUftpk3OTHveI7Z+ScAQ3gDEyKVKTd3cKfkb+HmIeXm9fqjODwhKxbIXzXmm5LTrayvqLoSdznWi108s74VXJx4qt4Rxz1mnMXIyF/PLjZMp1pcFRq3jMbK+KdkrnWcQKiiCo72vGDJjqZ4XxMRCVk7tRVR/GjrtA1jpHefucxYUFwIQ7vmUS5e4VHRfBV5yIwEVMLKRNoGpXiqK0FUrF6xWytuV8wti4fePG3ZmbsaK8gI4Uhz/1k9v2sPVDUsVylpvXA5xAvGvG0B31eUDqBQJTvKLxDsBxQEIkxpHByL0fQEQjYG0H/sJ4EWsjTC2FE45r/G2qSBz1OkEWbC2QBB5X5DztToqqtPlLs8nAI8Q+4jgFaSmYn4xdPNwuT0/Iv2c5PlAYpDUjYILN0qOnaepbsfGaiWbHx+xXK+j8SMeGpuYska7LU+UT27ds0cr65o3dIDR6cYZVA1rrN1p2c7ujt7PC6Jcg7P0AZ5ZQ+xfgGd00FDIp5sGENAVDlzkiqKwCAOQQSF0Er/SedE5sslixr719S9bpteRfwvx1uLajq3tNaxlecuVqyLd0V0sIcwUJB+K0fjXIKfVUm4dJXvo4qHjg2cAsKZumqC44FRaNyjm90XMEOlyX8RZ7lFpB/5O5aKVkD9LQzQ8UmcFxWluZH1zSx07jNP6+rbAPDo7qG10unQyUHbp2KsvvaTusvfefV/ensjztbpOEJN5ecjLXMobGR9kyH3fHRAcFGrSHeIEh1g4pwivOROktbhv6jreRezdkJynMo2nphXl3BEvJgdXh6wT6XrAfBBUWHeK3ZFEwF/i0HKpnn3puUtWzPWs3zq0G09dsdFaxX78/bdtYrxmnX7BPr67bNNnL9mDlS2rt/ouC85hIfEQaC3+/v2uKzgILAqdmdHbhitRl30wheYe2D92Pn15EOnMXP+pJNFZp5AV2HFcJp5Y1lsxWTsaX+KY0FEtcDJ0c3HvTsxgHnhXBd1v7Nl8P8pIx5wlxnZx3PU6khjrW6VYtHTv2J6+etkWZmd09uwf1mGXqnOCjgrW/tkzc7oWgGsIIIw1APHmxkZYy5Cm0nbp8iXldbdv3ZWvKteIvCq1Hs4m9iI+eE3mCnN4IN0VyORPOioeG6I/+eav+wiM1htutKWA1rVidaAEHwq1QoaWUH5Hm09oq4KlBkLqi7qvtmhQWwJAJE5gX3JQUxxjEwLxRP7GTeXCpqTdNySoETTQBuxtk9K6DB0PLE6+BsBgU46JIYU5gokcevwwkcbH7Py585JyEC+41w0tixW1fBIQ+qEUJK2Chr1r77oPAMEHsjXr6xuuF83GG4suqmAFk28FrVwTDDTkFjwpIxihWEwg5GwOjJm8SMPntNcROMokr1hSVwgHfGRpkKBI5zhtMk57+eUX7fatW3b9xg176623lADm8yUlTwAzZVrTsykxTMZGSlYqoIfI4UVh2gEAtdlxL0Hyp1Cq2gcff2abu3U7ajHeOTHG6EIZqZRseqJm1msaxbcciK3TPwSyUMih0RIt4+19N8eDhZMJPhgEOTw/jqmD+oHMwmGCYdI4ce6ixpcgIVnQjCBX8kDW2GIAGdry+Dwmz0npp9hRQWE1tpADVChgKZXEPlMyD+BUrnqrs3z20lYZLZsDFX07arhBaGzFlelt+IhASpS1IZjlmUcpqBN7QTBBZB6rfZlW53RGQZRL5RzJwHl+asKW7t2xnbVVy+GhQFCVdSM6xkaBc9L0k8AWZnappHWq3xej0QvLABVMYVoHYWDQ+g7LiTFQV03wnohFAuYgGqS0JgvsC3I9vH4cX0VeiY9YeCDJoGjVx8is79cBKxsA6BGST/ceaHHrsJciGgGFt5hK6zHIG8XXi28Ri3yxMBSDmtjB4WDF0C/ncXtwDCy0FtXCnLZMLm2pXN6m5hYEVJy7ctXwOIfJhmza4qNFm5udtbML89L0RUpmeXFRrdMbiw/VpglQoedBMMp1JIJK5owKscde0PJA0CWcxGJhz5FTLXc/7KiQTF3srBgMwnDMY7Ck9UHASZfGcdcunF2QxNvCzJRVywUr0cGEb4xM3VrWODiUMaNawUOrPfOZ4Gdrc1tSFxUVBwp2b2nF/uQvfiid5xQcXHU8Px6oILhUwVXFWkzHSea8fT4J2sW5NHw+3qUUfTqkb35yasXDwFlUoVya3A/ic00WfGPxOr5f/Jq/ix4NSiwAACAASURBVGOnxDIYqn3RmX26EPm4r73m6CBi8mMg/wS7hbnZoRAyZteeumKZDPJ7LRUkSAqnZ+fstde+Yn/67W/bwWFTBXSAZ+3LjA6SCzzrLwAqwhWckH7yAN/XcFAXHBQR4/gNCoOK6V0yTh2MmFfCKGR/7LnfhWssu8av79F96/bbYinFBCuObyxMevLt3RRydAgF/dgt97ig34u53qUU508svmMO32weusdU8C7wGAWAJW0vfvlF+1/+539k/+oP/8S++2++q041Je0AgHRwwoQMBXARGmQuSGEF40sXnEZ7uFZGZiVvJSQomdtpL3LDqN2AkZtC61ejqDXtH578RH8QJd8BeE3Ou8EcCUaij597AeDwP/QCkyQSiDuy3tGW+Ijj6P8GRmsEQoL0E2dBt+dSWBGgGhTBdVYMZReTc1nSBEXXxj0NqHAJyBM2Oy0BFYzT1WtP22tf+2uSySJBBWQv5JCGKNp7b79tb73+Pctk2EeG3R1xbUs/OEqBxHmgPa7HA/C5zBiH30lezxcV7Qf7Q+iy4u8BbBkHmMfMB42b/FS8iySeJUnQ4vRcjGsoAhHxcXwReMHPk/GMvqZImOhsifGIS05Ajz3tDXJytsR7ToLXcR+M3xsWP5j7xzY9XrJxSXWkJHNUwbR4YsqakD96LkMUE3/JbgZAr4v/yImOip5ie2IeFTmj30vwkpDGdIgfkh2xALRxP45ghcZcXJfE/QaD7dN7PfkFZ/Hhwb6AiuhRQXEndlTgS0Gecb46Y9bL2U9++p7NzMyqmIF80/Nfel6M23feecfOnT1jk1MTYux//PHHKnx/8vFn9uKLL8s/6+6dB+qoEPmo27Rz5xdktIzsEvriABXLi0uK1b/2tVctm4OQdSBpEvlCHbX1O+1W1z75+FPJnWGIfNzFl2FfPm54QFAca9SbMv3e2Ny0QqlgjdaRDJkBI/gXQgo7L6NFsXyCToKdbf391Jl5++Tmx7a1u2Pf+q3fsvt376ur+uKFi7a5ui62PGOEFJBirU5bc6BcItadtNrYlC2vIg1q9uDBAzH8FZcBBoU6GfEx3eDyhEubisJ4VPDfSy8+b5/d/NCeun7Nrj77tK/RdErXXt/bt3v37tnW1q7lcyWbmpzVeHQ6aOBnLZNPWTqXkTQQxBWKNkhfEJOz7l0fHsJNW0X+Xrttd+/ekawK0l2as30TAQomsTqh64fKsza29gQ4cysqVLbQMm8rjp5fmNfcdR86WLR0tHdtYW7OuscALO4Ts7t/IF8KCvYAXBh8T46PSSKwVMwJtCDuZo8lN+O15AEoH0aK3fgXHGvcILZJGvi4pW5nznbmfrPRVGc/fml4Z2BmT9xWqdUEpkTQEDNu1g/XXamWQ0cI6zljtZGqe2ykKKyTs7hXJPuOF9O9i3cg7Rd06rkACvMQCAEIAHK7HVjdEJmQGmurU35xecU2d3YUFwBaIPtTyNJVgb+gk7EYW+V5oRAa82diStaffKaOGWuK0+5lQKFOf6d4wTRnANXJTTzn8XwYsBSQBnmnSjFnU6MjNjs5YmfnJq3V2JcMV7VUUIEYPfg3f/qRLa5tWSrPuekxMOsUIMf9Iry7x1UNHJBg7vhcYOqRc2V1n4AmPKtImGQM2R/JWx0c9a+5n2T8GQudvB57pYyWZeyOIXVDeVDE5JXHBAka5os8J3TWE196jDkEz2P8EQylVdkgFvJOalYtYJH+XvyoY5ubnrDzM5NWzPTt/MK8LS4+UqfE3l7bRiZRtOhLAq7V69v5CxftSN6eXeXxSEtLDjiDNHVBoB+5W6lYDnO9oC4hSfChSgHohB+mCu7UMVxyWt2wjGPQ1AdgiDkZYMpI+thevHHF5qcn5TeChPRb7900K9Rsr9U1yxa0DzBH8jnyXEgU3uHhgBzdJE66YA3sbO9JkswBdYh01FC8k0eeIgKa8if8STY3t5Qn0V3Fa0jyvNOSFDDdiAUM1Yt5EYo+++yWrRLH67XTAiwkj4z3xjF+nMGfJpWyV1580c7Mz9sHP/vQHi0uWSZfsBbnJyALskDBm4G9w7upEz5ZIQbX8wwgVfR5ibLXmlfIDB3jZ3GkOpL7PXhXNCRLjw9dKSSTdrCJnwkoQqAIOS22dcZRJ40DkQBgnVZdBJNrV2Zsf2vHMr2Ufeubz9v01JS98cMfa8zSuYq988FtK4/P2NLGvjWPia2I23w+8h//U90reL7F7kqu1etdbj6vuR7j30xWShAP3746CILOfukj1Tzk1xDI0Yp/0l685z2y+KMg566uLydOxk4pkTcgfUpWHkKAd4WyF0nBRZ0VXhM8Hd8NgIog8Qv4VshAdDK7coFaY1G+Qnv7hyBymhdk6igjzM/P6rX3dvaUnzMXiVd2drw+xXoB8INUzf6yurrmxFHJdfUk8wXJDZK2nmuof7IPA4TTvcn180Gt50lHxeOzrCff/TUegRqTHL06FcD8oORriiwsLrExaCutVh2pDYchC4zNVRuCdNCd9c3vEYDs7+3pQKDNloAA8zQYQ0gl1Ko1FVEJvthkVVyW8ZUXZgmA+L5raeYVwHBwwhTi9WCJwOwHdfSNzdu9zi6csanJSbFy+D6ySUSsI6OjasejfZWFTLsczA0vpsQCiSfmAmjECnH0nL9RK2PX26C538i0YGzYSBg7gmJ1VQTzSoJ2NikCIYIdyT3xuzrUTHqvdJxIb7ZPS2BZoAPBo2KNwMbjXmEsaEPa31OyqHHJF/S5/C+sb1OTY9LIu3j+jAEPVCsFoeLZrJtCCRw59iBWjLi+2fTcnG1sH9ib77xvpeq45aRrC6vu2DpHDZmVTY0RnOdtdWnJZqamJKlE++ZTV68p+frs7l3LVyrWaHasg7cH+n3lolgQAFXMF4rZfF8dFe2mTV28rMBmyNYL0mJBbzYeCjEQSQIVsaMhsvpiEXsAVChgRuuWQu2eQAJYnrXRMWf6YKZdHRkAFRSvyyMOVPBx1KD9Eqbg0KMieWg5MOEgV5Q/iAX+AQqvJNwLrZG9I7AvkxEDK1vIWwvmRKdts+OjtnTvlh1srhkhGAkQRYsIyFCsip0MGhc6jNAFL3kbO+Uy1qsHLB0VjyiCw46BefJwcdE2tjYHHhWsEw61WDQAqBBIkcsGIz0Hj9yrxT1AkuzxWNTRs8tRtGp6UalPYcRNQdc3tu3TO3dU7IsSQO795YmT1o2KaMNAPAJWsUCUHPMkUCHDLRJKMUG9Df3zH17M5CMGxQMvjmzWpucW7KWvfNUWLlwSwwUTw/2dfXt4/4GAvrPnzlqj6XvbytKibS3dts1HDyX9FDsqnAHl7zyoXQY2mSxIAviZSoeifjDYi7JQFOu6KRdD+UVAhYpc0WyWMVOx4Fiayc9ee8oWpqdsrFaRyaPYPUSevZ4XGQCeg0RdBL1omX74YNGmZ2dsZGJS+/F+q2N/8eZP7ObHt6zXI4Ej/flioELJkILovphUPAsScoLIJFP2ZEE/AhXOLI5ARdIoMIyos/SGAxsSuGhq5uObNFn3r2On3LBTLxa9I4Dy8wqLvxio4HU9iD1xX4G9JEabvGfAc70oMTM1aWfmZ1UYAPTG/JQEBy1nDFJTWSQSj9UaL2Baskk+scIW9LmgWe8fLBn1Q+0XLpsYi7vRLyG5l3oh1ouELoXmwBJSPzJ95POery3tX2r1Z292HVxYpyT1sNSS958EUh1kjEVXD7bjz+ONnPj6C4EKkgjW99GQ8a2z2ecdicqZS2ftf/1H/5ttru/Y//G//2Pb29u2TBrtfK4PWSfvIJNWbSpl83PzKv5v7mzazva2NMxhh9XKZXUvUoCKTDDOx73DupJSyJkCcfRfvIvQVRGMzH8RUME54PMz7gfx77mhoWp1nIMq2FC4ISFOABWxKHICvGTuBwaaAJ0gbeEdUb4Haz4NugeIe7yzS9MndO9pv4QZT2dfQsZnuL86kAY7uAUJolSwL3/lq/bCl16yTZjTkC/UUVGVqTGFzL/4t//a0qmO9Y5hNob3E9DkxYUT8zSAvscU/oIJtubZXxmo8HMY2RaKU8QcAq4kredM4CH4MTTWjuOSBATi934VoCI+ozh+p8/RCJJozajn4fFARYTGhtfqrxjnSnx+Yi0GQEx7fapvpZzZeK2qc415RCo+d/GK9SABcWZrrfY1Pow7+5DOfLpAJY8x9AMjiZYmuQxq3f8kMjjj78U1Eq81AhUx7oxxB9cfCQlJACbO0zhmnCmcY5gdu940xA+ARu+ocOmnoj7/3v85O5yq/xE+SzjtPPbdHt9/88teWCxIDl/ltKGu5kDoekqC+r/sO/z7+r1YHB28ntdaTxANftn38nuMH86BDrP9l32J/wJ+LwzwfwF3+uQWn4zAkxF4MgKMwNT1d0VE5uyXNLsAh7T76eCDQjde9IqlkweSdFDjQBpShKfQoapaHsCcwCuPzYlvvOPbjcqTMdYgjwIcolaZzViaumM2bU9duiDCE0AFcr59OpSQSJN3kon4SDfv+saOOqiQN6Q7EHAd3x92c7pAFhYWFFfJ1zV0nRGD4V+1trFpI7WaYjOARPzGACggNOCd4l26Lgn2BKh4sl7+sxuBqSBZREIvEx7aFAetWV7YkJklci4qumfEQpeGbiwaBNklJbcUSANbHsBiTYyevlq2aPWlVc9bv6KhkZtR06IJ3YCFiGcEBQXACv6Wa0DHLnYn4N0g+W7aWSkupPtWrpRUkKPIQ5Ea9hrgAO25kZvLIgbl9xbG0OIW4mDX2KUAQkusa7jnc651R0LWta4M9eSnAVu93vAOFBkDwjrge/VBC6nGodPWRonxjjZMDI6QvWq1xEzw9mjG3E18AC4AWdCbU3taYBXLTA+ztnTPXn7lFbUpvvXmmypW0zVy6fx5297asN3NDbWh0SIJA6Xbo82YZNw1SUmE2dRkoIpEDIXkYtU+u8cGS4eEd9OglTgxMmLVYtZ6x00bRTIAz5F22yqB4bO1tWWZQtHGJyft3sNFsTFSakvuylxKSXOqL1SfjopWp2UYgFEgGD93MbT9eoGdD+ZOBCRi4qpxD1rIv6ijwlkoblLN55jyNdQWfqzOFTQtY6EOXW3mulpnHwNUyAQqMGYxNU4eWrHTIRbs49exsDNM1rxgRMFFxfTAEAXIY9yaMHvbLRuvlm3p7i1r7W9ZBmBJ7cDeLUASzoHER+wKEBsgtK8qSYcZPShAwZJEazOrwhqgwcrami0tL+k1JPMUvCqGQEVBoEYSqJCsVOiq8gPzJLvfiw4w9zGIq+Nja9lU1jKprO0dHtmnn9227b19t2tPA0Dmta7E5JCxHkVI12+Nr58EKpLP/3Sh2U3dhiDRaWa7j/8QqIgseq5Xe1cmZ7Nnz9mXvvyazcyftXr7WCaXjd19u3/nno1PjNrZ82dVeGcNLi09tK3le7a19MjaBATat1iMw1bt4egEb4ooB8PzT0eNeC/MJYGKXvAG/2WBihg4wVCjywkhp4tn5uzqpQvSyZycGFVHE3sPc+OojryYF58o0En6C5Aql7Vbn922yelpBypqI9ZN5+yDO/fsRz9+S/JPP6+jIlnQj9JP/CvTyP39EwXRyALy5/J4oOLzh2oA+RJEcp+DXiiOxdo4T+LXyQ6O5DWeZh1/0SH+7wRUxK484B3We8rPslI+b2fmZ+zMwhmZZ96+e9fqdfbHnhXKZckKqfAnvyZvaXagg3lzsmsjeX0/F6gILKxYCIz3H/c/vpb8WwAkBkAF53gCqGB5uv60F9hTadezJ6AXAyu+jxjhQy8EQF6knyT/dKrIHvf6xKZ6oqMi7ge8n4CKblOyNAL4g8eP1kHKZGZ64/rz9tqrX7W//PFf2oMHt61SA6zp2ERtwva296QjPj05bSO1qo0DVmcytnt4aCtrq7a+tmbFfM7GR0etXChYng4MAb2cUzB222rzP2wg/+Rafr8KUJGcZ1qDQUIo7lGD/e+UF0n8O/cPKriudvg4zaaPACYvMZDuGchZumRTsqNiACSl3F8rebYJ7OO96J4UO967LpL3TDdfvdmQxEGpWrIvv/ZVe/6FF217r64kDMJGPl+1XKZg92/ftm//8R+Y9Y4khUAxVWs0rGH3iQodPIAYNFKE9vuefKIcMBNt9ASoMAQYTq/ZAfgSTheeN8x0WLKRrc1rEYdoH4+gYACi4pqJ8zQCoHHvPQ1UnN5LfvEeEpiy4b3jOQyb/5cFKmLskQSrTrNvxVzmUaZ6kjKcHBu17f0962VzdumGSx7SPeGwpRuRsgcBWEjWtI1kqJ/fkcFJHBoZpxGo8HFxZqfPmWEnDtdJ52+8XogNkU0Zxze5hycBzziOxCLIn+7t7QTAFAa0k3kkj0Y8E4CKP/8nc1+0tf8H+36AlAexzGA9/Tu+o2CKwKSN+8TplxwAJb/g9/4dL+WX+vMhaHPq12MH/i/1Kk9+6ckIPBmBJyPwZASejMDnR2DhSzddHjcqGkCooINMvq5d76CQeXdG3nLqmBIJx2H8GN/yL7VC5VnqsvDucTrtXIbLjchjXhljz3hFxMDlUt7S1EFSZteeumgLs7P29jvviIAN4cvwZ+FaMxmbnp5U96A6elMQPzwP39vdkzw8MoHUPGemp3SN6xvETHRzZZQP0j1Ezoh0IfdKHgnhtdlqSQKNzgr56IgMmXoCVDxZPP/5jcBk0820CfgraGFSZAkLm4K1e0AgQ4CxdlstmiwukhLaiNk0pIEe9BW9Dc+THlBCWsgwyWEjoPhPSygbB2hgfN/I0EIbGtAiekiQANHVwWu5Bm5G16bWLlqmKJ5TxOjR7eDAB6aYXBtABUV3mK1cW2yJZ/OSYEPatbidEeYFIQovsMBlVtRsialOa6aQyg6FfJcjACBgk6AAS4BOYQPZKXQGGavIKo5jwjhIMqPtJmRiy6cyg1ZE7oHEEgO6nZ0tq2KK1Ob9vUuFMYbhvre7I7Y3nQz1gz2ZHdUqFbv21GV7cO+OteoNu/70U1YqZqWR3mxiQBgkaABK2p1B94wYjfhLpHK2f9S2Dz++beNTbujXRyqn37dauWhjlaKK/8etpo3RzZJJeTdLCbOwYztADoC2S8yNMPlD6qiLoZW3I8Lwrh8dSgLqqHWkn42fvzjQ10sCFT5HnKkXCw4RoPDvU+D2jhDXaoU968WV2FERgQp0SwEqJBNWLFk5ABU8T4AKSRsJqMhYqVbyjop+Sixbl37ywijeGoOPAJxIzzEkYNxvlH46WaTwecWrcA2SfqIzqVK1dL5gTWl0tmy0VLCVB3esubdlaUyeZBjpBydrcmx0TPN9IOnAvYbCACCdPCqixj/GUD3amh18ANBf29q0h48e6aAWUEGhmqJ9kL1QuzXgWM6L2xyOtJDGTgTdu99s6OzwQgst4vi9tI6bKjChbt866tijpRVJpgCC0c7Moe/eMS5hRQFWz3Tgx+LFKACFyJ7zZ+9ySbENmnXLNWlNS/P2pCTXIIhI6L/HIp1fr8vR0H5LJ8ULr37ZxqZm7LDZtN2DfescNuzOZ3dsZLRmZ84uOHOz07HlpUcCKjaWF+240ZQUgxe4gvST92WFD39uUd7JPX1cH9i9OUKFVf/QTu/8DldACjJSseRBwUdjH1rFo845vPbjtqWYd9a3Sj5nN566bHPT4/Ko4TkChmLo2WP8W20BzXRf0c4OmIB0xOKjJe1T0zNzAiqsULYHm9v2/R/8SLqrrIXh3hjaeIP026C+SQ0RLeViPhQhkX5oeWE0SJINu2Yie9v1iQnYHi/9FJQAh0MVuidiwXRoKjtguQTfgpNF3Dhth7JCpxnJp09zZwgnOJyJQq4eXWxPflxHReyggeGqAj/sZu/uYs9kT0d2AN1rgdB0LbEvjY3aM88+b/liWZIPqyurdkD34c6OddtNnVDJgDles7dVhw/k1CjiBw18H9fgiaL9JIAIodgegQrJUPAs6KgCyObrvneL6b8g2+bvDziHf9Oxzj7mFHMzgqQMlb8tf+ugeAQqoq9MfM2k3JeDd4EdrvEO74Vpcx/wBhM8Oju8e1E+FJL1cVNKTGO/9Ru/afW9ut28+Z6Nj9Ex1rGxypitrGxq3p+Zm5dMhEB4gMl63Xb39gRUoAk8MzEp6ScHXmLDOvqwDmLu7tVlmKjOtsGoszB9jP2eoQd4HPG450UBfjizw8KOr0VnVVjsJ4A4QF6kJZBgSLDt1SY/kIYYakkMgQpGiL3HzZAjCDyQ5lI3E3JWYQZJjs9NFrXzZl1K0OV8/KzzD7Qxe5KoOe51rDpata99/Rt29dp1W9/a05lPUpXPlnUGLT96ZH/yr/5fSVD2kVAMZwjgBGcRXaTjE+PqeM0Vi7onzm26cXe2tq1+WP+c/FtyzT8uGk8CFVyvOvpoiW80QpIbZAMH3QBDsDxZNHdQzxPdWECPoHnyrInPO34vCZzHa0lep+8hniD7+PvgysScPTGSDgI442eGPxifV87F4GyRfEMYU15FMV1I3AUIZJEmSEu2BgIMZq6jU5O2cPGSZAkU2xNfhs8FTgRiCDGQgAolzO6bAMnFJRU8ho2mnZKRw3Q0SD9FMIx5g9ydAxVIRjkxZTAfEwDU6e6KOI7Eaej0E/vKRwcSSigkJKWfSP6//38vPG5K/Ef5XpL3/6vy3T/fURh5nz+/KyEJDvyn7KjwnSHedYJdkBj5/9TX9x9lEjx5kycj8GQEnozAkxH4DzICCy/cDDGJS9x5UOT1CepKxANE6MQi8qMJJBfVA6Xi4PGMxz3urwuRT95X1K1k/j30L0nme8mciIofpCYUTPB+mZuZVg1gaWnJmp22AxTIpXXpGE7ZhQvnbW9nx3b3DlR/kcQe3keNI5Ew6JTAEB3VFGIbOi2ivB4DSSxGzcZ9VYi1UM9w/5zopYM6DTUm1FeedFT8B5l+T170P+UIAFSQeLAQZbJMsT60d+NYT3sUSQRJJcVzNgYBFemMm0r3cSpIqSPCJZOcNQ3A4GxqWFT+Pdqf+B2MvngvCpkkPyxatDjFqMcHg7apkIxIdiIwuySHADs7Q8cBnhrO9Mzm+botxFHhcmB7svGQeKGdSHEZBrjLn3C/noTSWuW6ks7E77SRLnJNY7Qy2eAaGM+mzXLFaN6XUnEPsGV1dUUbjlDSkIRxnzIrDjr6boppdoRZGsnZQLPfC7Qb2zv22quv2Llz5+3b//Y7ls+6tAXXGxNtNibuR74AGLLBKu80ZAZKEor5U/Pw0J595rpM9yoVCpW0yMPwDZJU8t9IyRSKDodsvujSI6msrW7uiTkqHWKM/nZ2pGtZSKeskMtarVq27Y0tq9XKMuWDVUuxqFAt2eLSirwR6Jjg9Y8wN0uZ5LpyBRLkht4PFiOF9LGz5wXcSI4naOtJskTFYQcqkom/d1qgQYiElXtU8OzV7cLBFApratnTAdZVSx1gDgxBCoKV2qgXAZBfqo2aWgEpKWezVqg4UMHPuS8HKrx4luyocJ101x3lPZmrCEhEeaN43cOCqBclJO0StN4pFkvzU8/k2Gqlgu2srdjm8iPLAZwEtr6KF9mspM5cP9FlV1zqwA9etGVphYxJfhfDMencOxMWIGplY91u3bsnWS70GzkoAcWYA7wWnTLpAnIfkUXrMm98eAtksmDpIJ8OxIKvfYzvtUYaTRUlDg9g1rKevEDabuLPgf4lMkyezgI2aVzD84jX70wJL6CcLu5EmbD4XJJzJLZqJotysdMl/p5AjnTOsqWKnbn8lD374stWGR21vTpycHXrtTt2+9Nb6nDCUJH1S1F2dWXZ1h/etY2lh9ajIyoYlUpKLRSPkkCFF169eOlFJIqQXviLH48rmJ8uajmDe1j0jExe7c90mgGIHPctm+rbwvSkXbt83mpVwE50LPELOrLxsXEFY7BmNzc2LZVNWWWkZtVqTfvwZx99bPNzC9KITpUq9smjZXvjrbfs4KDueJ8+JOZvXQPQHkp1xSIb+32hVPQiGoXGFueFSxB5wTpowoc1HUFIjUdgxsR3Sq6f+Jz5PZ5l3CeSY/i4z+PffdGZ+rlxPrXXJIEKxcBhKxJUkwAqTs/PaNwM20Zrb+AV4F01wy4fL+QIIGQNVor22l//ll28+oxVxiasvn8gv5rv/H9/bDsrDwV2xLmTnEPJ+Z8soGpuBXA9yQ7nPXXvPKewT8f1Ev/V2SRm95AVrTM2QPrHRrcHZ2Rb+6Qz1H2uB6+/ADBzxgFcOGCFnFKiseJEh5afuj5HNDLMoaOmgxcpl53yZ+b7ggq0wTSbbaJYytjv/u7vWDFXsTd/+LqN1fJWzhMT5Gxxbde6x2mbrFXt7PS4FYs5a3S6tn2wb8ifHey6lOL4yOhASo8zCslGbgiDSYCK7Z0DnRWR2e+HQ1zPfm36f/hWEjAbnGN4+XzB/EFDOBaoTz8zf13XDXaPH4BiB0u1D5wC1uJ7pFIkahGoCADqoLuCtecxkMCkUPyOa77LNAhAdtL8Wedhq2OtYzpMejY2MWa/+Td/y2bnz9jq+pZYYQChxFjFXEF6+n/yR39sh7TDd4kZ0YfOWaVas4nJSRnBostbLNNlSIzk3bBoiq+urNijBw8VWyGn5r4Hye6Okys87qnJdRFjWjpXOTvj3nMCSArgZHJt8fnptRafj8sW+rjH33kcIPHY/SdqBZ4CPX3aO6lBzz90MQz3RcAo59W73GjcpQIgGaS03B/GnzUfnLewC4nN3eDUJefOnDkjSK3dc88uCBTsV8TQkgeVbrPPV65JXR8p19FmzgE0xZgmSjrFMYtgRdxvopk2X8czPJJT4u8MwJlT3Ve8vxtJNmx3dyt0AntBgb/hdRz8KCovmMtPWC5bsps3P5NJMXHJweGevfraq7rHt99+0y5fvqT5ee3aNXv99R/ZzMyMffrpZ/alF16St9SDh49E5qGDA9+CGzeuWa/bsvm5abt367Z97StftTu37tjdO+6ZkCum/EYFlgAAIABJREFUrVTK2Te++XWrlEsC16q1EWmlExfn82UnhmSztru7p32i3WnZs88+qy5TyF+YbGJmzX1JGz6VlncGxCIMms9dumyldNq2drZsZ2/Ldna2Rah69ZVXZCJNVMX36vsNnfXkbzw3ZGvz1aotnDtraw/uWl4mwQCmdO32rdmCGFYWAYjx0U5Gx3cbqdaezczO2eLyku3tHdiFSxdtdn7OlpeX7Lvf/TPp4iP5CLC4MD9jX/nqqzY6N2u9o4bH74Pcp6S8Z3/Xiy942zWb5FhVa2LKS+cu+1iaPKagIg0EHEhyKspAcskX7KCO3yFd4tEfKmUHB/s667QnBrKdv55rsyM3zJhPTU3Y+fPndWahr85cfeONN/T3EJ6uXr0qMsny8oqYq9XqiIhq/C3zD4Ng1tG5swsypEcxAO+/nZ0dFYpqNaTunCWrPJi5idxmUAOAiNY6OrTecVsxZQTflJugJKA1JjdFFa0gkLBeeU0eijzxMhnFdDrb005yqx+1bGdvTxLI+EMqr8SvsFTWmkHjnfkYgUEV8sjPJXficZ1yHohnhaLOGOXdZPThPTgL6dCGKLS2vqHnhzk8ZAUOPFQDKI4hvwwY32k2FTGWisEwGX+VNqS3gpXKZfvSl17U2mCp+xjv2NbmpgiQkBTxKSCfZV/Z39/Tmnjl5Zc1dg/u3rOvvPqC9fEsqLtHxfTkpIp9vVTW/uL1d22Tv0EMOcV8yjsBo+9xqVQNgqwLsSrfp0AYfSRYz2JfQ2ySibYb2Hr8jvKD1yg4T6Q8EWRiWNvUHhg78kruDflg5qLMnsN76i3Jn4KvT4zb6PgXwTGcU9rDgxw2c1VnvZ6Zg8HD2Fitt3qOql/wTFkPxErdnj1345q9eONpu/vpTTvY2bTRasWmp6ZF1qKz/P2P8LjZd5JhtycDcDxf+JdnhZcdEs4um+h+HJAzqXv4PmLulYgUNz4hkvHuyZw9Es0AwuMZwfjxrETOItY8btl0KWVff/UFGykXbbRWs+2dPXv7g09sv2WWrYzZ0bH7oBwft+VRwdrOZJwYxZ5Pp+Tenq9jjQtnGiQy+Z45sRR2vQgHsXsyja8Q89zPXeZdNP5GIhQ8HPnrSxfO2v7ulo1UylYt+bxcWl6Rjx/enM88/4ItLi7b3n7d8viMHtVleI8583Gnb9/8+pdttDZi7737ni0urVoOgit7s87PkP8iEQ4pMRailbcHckLMvoN3KvcY52fs7qWuxdxgniK1zTrm9ZhDnB9Ij8hQm90F6fGuWT4L6fjIsup+7FulUrAvv/SilXM5yaJTN5iYmrLx8VErlQu2tr5o25trtru1YefOnLGxkTGrVvBQKqjreHF11Zp4oizMq5YIibit189bvlCWdCoePAf1Q7v/4K49WlwUqZcxT5KrmMItrSvvvNRaDUQ9nh33SGeyDOrbHT1XD4BdZp0aIuQ89iqAC9XfVBD0uo+ACnYnapYYd6umRD3H45m4xtyY3f1i48eJ+BI5+WpFJuujlZKdP7MgxYL7Dx7oOo7ax5bDLwRJ3l7XFubnpLayu8O+5zE30vqc+07Q9Hge6XuIPuxJSGZy89Qi8bbiXJCsFd5ceffZldRyoyE/LcZDSi3l8hOg4rHB95Nv/lqPwKSK3s7kkuarpH+cFYs2LExQCu8kldKmNgLcpjZ+2vzZ2OMBysHsxf+u2LsyoVZgTmBXtNGRESuVqlpwGEvt7uwoeCSgYj9hsyAQjAETgRoFXXZuBdJa5ATZML+cye4bGQbdDV1rpVRWoIGhN2x0AggWt67NnM2NjjIBNoEzgdI+ASumu92O0E4V8iiEH/eUMBSKZWf8pWDmHelvGBNM0DB784OCjoddGTkhfxJb+rk/mamFtvoB8+3Yi+wy76JYMj6uDZND/vd+//fs9R/+wJYWF0NQ4gxdmVYF469iIWcvf+lZOzo6kGETZlM/efMN6eGNj47I3A8DbKHG6vRAkxgjno5M4XiGxTIHZ0/yT1u7h7a+tWtNGNhNN68qZjM2SyC4t2djozWbmpyytZVlBYBTM1MKcPcah4POhoNG3Z8/QVYmYzu7255otpCKONa/FKgn6KgIQEUs8jtQ4Uz500XoKAnl5qAOVKhgGwJAL845q9jdyjyYbMhfhGSsZNURirZexCtXakooOJCRwSlVKzY65h4V0mEOvgePBSpkkObvT7cFh2Usop4GKvxrlzric3XjlGGb5l3uq9d2M7iDPVu8e9tyAGwUoENxjt+PQAXX5Ii6g23qqgiyFvEQBaiQpAsyTByAqYytbm3ax7du2QEFn5SvA3wLeC5lJLEqFcsAVOTQegTIILgouAxNMOjjUPfiZTAzQ0Yowz10jGfOPkFSeHTUCpI1vlYloSZmJhr86Ms7c5hDORb+4t4zLOR+fjtl7GKRw4PLIUs+BvtxD4qF7ShREYN6/r6QLQiouPD0Dbv23PNWQKoI35rmoSSdbn36md4HUzUOfJLKlZUlJfmbiw+tK6DC5ei+CKggkIzsZyUkCSmM00FP8k4/V0APeu6xqBaLbH4/UGoRpTdL97pWzmft6pULdmZ+yuZnp6xQyNntW7dknjo2MioPCoLY5ZVVdc+MjY5rD6TgQkI1Oztnrb7Zh3fu24OHDw3ps88DFa0ThdZ4PTw/gAo+CJYoonlxM+if/xWBinjf8d+YoCXH8HGfx+f9RYfyLwIqCGyjEs+vAlQM9iyACsCAAVDBHPCAOhahBZrl3OivPFqzv/sP/3sbmTlrxymC565Zq2n/9J/8Y9t4dDd0ZTi4cbp4ehqsiF+7/4eDlXFf9Xj+80BFssDoxo5ewE7+vo9lMKmWf9Sx/JSQ5xGbmoQAjrZq+S5O57UqvwaXihw+kRPPgCQsVmH7fWvC2kbaJch88beSIwofce3z+uz3+ULK/vbf/l0bq07aG99/3cqFvlWw9clm7cNP7lsqVbS58VG7vDBtlXLBmj2z7YNd29zetsZhXcXXkWrN4wTJ7h1bR12YaRnN7h0c2Nb2vjuCBFDGg44AUPiTcUDyFwAVcW4mnxvfQ+IqPofTQIX8JuKzD14kEUjSI0lM9Pi6Xij0jgp1c4XW9lgg0PPN0DkTgIpwP1rTdLFishiK9cQnFNEEFAFM03EoecG+zczN2n/9279j1ZEx29jeU4GN843CBUAFc+Tbf/qntra6ZplUT+3ytZGaOiiI1ficvalcrVmuUPGCUpNzu24rK8t2+/Yd29/fNes7kBPn5OOAgQhiJMeWe2CdEQvEwnocruQ4e2I/HMnHARX8HWPpIPxwPfsz9VeN3TBftPcMTI2+AKhIvtDJtT70NfGzJXYf+jUDagukiGB4uBWBDFni+px3KqfTik/PnTuni23TERRBGYCK4FFBXCUjzlDw0D6SACqYE3i2eUeFF4NOAxXxGa2vrw1uKwlUnH6enwPowiASp1Aw3N7aHOwjFGDYO11CIStwgpgIoCKTLthHH31qtdqoOphbrYa99MpLKiy/+cYb9tzzz2k/uXDxgt29c1fr/MH9B/b00zdEYMKUmmJ4u02Brm1XrpwTyDY5NmaffHTTvvraa1Yulmx5ZVmdHs1W3drHTXv2uRs2OlINxY6M7e3VbXFxRYVDroUOLnIEujXX1lZtemZKUrgqJqng674b5BcQxMhDor8dZziFm/HZaTvuOAsTfyOeE2b2xLc7G5sC+AB66YzBz+/hw4f2/Csv2+zsjK0vPZRcJIUccKz2MQbUR1bCM01Gt0159FAsh5jFMwYcuHLtqtbQhx/d1D5y8dJF+fy99eY71mjseTdpry151aefvmrnL19SLiPCWR8wKacuS4r6GI3X603L5koqfpNrEC1BoOH+YYpSLCb/85i654VzdR+WladBohGQIgNUCjZ1FcdcYrccyFw5dXm+9dZbtryyZi+88KzNTE+re+j+/ft6jVdeecXazZZ9dPMju3XrtnKmc+fPK1anI7jZbNvhYd3yWYAEiFLHNjc7bfkc/m0wWT0e/+zTWwFI5jzqWhmPxnQ6yAymVUTifsiZIJCJnKD8gX0fv0MH3dhbAUD4nByNvJr5RzwJgAO5j2Ibr8W5VMLke3tHHcGc9+SFjBnjMTY27uMo6ROPt4ntkR5R3iMZYbq0naErHz9puDsg6nsZ53ZWOR6xogr07ba1W3110sssHE14GMSdpohxRwc79tRTF2xmatRGq0g9l+zBoxXbPwSg6dnzz7+gPf39929aPu+eeHhKch6g2DA+NmatNhIp+ypaMyemZ2Zs4cwZ21xbsR98/3s2PT5mo7WSjVerNjU5KtNjXpui4JvvfGCb+0fWy+RULJRCAvk+Y5/HwBhCo5NeyFl41rxvBIb0nAoF3afnFW7UzGtQQJUHZ8VVJKIsnhMqHQBkH2S+i/iI7rxIlRl16fM1RXbACi+EYuZNTu5jzljzvrGz0oF538h5LswJ9o/okchck7RuUITQr+r1JJat7tZ5pGTaRzY5UrVixmxtacOs37JStWZXrl6TZPP27r4VyhXLFYqaO6x9zkvCm0wwI6buw37EHKQ2orNQBVavX1DslsExQGjb1RSIA/hg72YSkqtS3+A9GH8R96xrMyWzF5+5ahvLKzY1MWpzZ87Z62+9aztHPUuVRqzeJMcmW4QFL9kLgSwUuXlWvB7rVHNZ+waAkftfct3UoBh3FbODmbbAzI4DSTrjol8WYCcSOv1jy2XMzp9dsK2Ndbty8bwVgifjBx98pGfX7HTt6vVn7IE609uWyeWt2T6ySq1iR0d1qx8e2de/8qrNz87aD77/Q/mdpTJ4OnYUR3JPHnMEEk+I5ZQ3y7fU6wqAP8NcSCvTz/yQA8eYw+cK+4gDNCKg6AkxT1yJgjg1m3bSI8ojnRZgsNnC3HRQz6hYIV+yQ5j+RyiI9G12bkpAfKmYk2E0REeZbvdSVj9sqG4CAFMbHXFfRwiwaVNnuEy5M8SByIG3BeJMTI5pPSwtL9vK8rLqJ9TQdvYPBXBAEGTP0vwK8ZbLyPq9Md/4UC2EsyU8a92d4vM4kJ6ycPfRt0uAWVA2EDki/MylpDlr3HsvxlHJWPJEzNk7lpIJXpEQTZ9/5oY16of20Ucf67wHON7aO7R8uaxz4uJFpNm3RDBmYQE0cB/UTJijgBCRjM25Rf0FoIK9gT2SOJr9XrGCmc4YwDmPjZqKgRizKCX/pKPiCyPwJz/4dR0BOirEFBBLkYVRcPY2Pg+gzUFeicCExcX3KETD5mbxEgCogN5qaRPjQMhYWoGi69ETgMKk88WJBAwHSyDdOEM7sMnUQRC042TmG9qbIntBB3YIGHg9Dj5pz2f6NjJSHbStgxSzSfEanrSbCvNcG4sbhJ7iAEEY7fG6LwoUGNTWRlRcJRgr5osKstPZnFgHjWZTDJW9/T0hmgR3vJGQ3m5fYyjWuwAbD0SlF59xaR0CRQ5OgshysawNiQOeA4kDnX8xx5mdnbeV5UdC/WPXCEFVDCq5Xjobvv61V21jbVkad8gyfftf/2uhtxi4NhqHIoBGAGYYRPFMcwJqQG/7sMyLZfvs7kNbWl5X9wHjDFBRQKqoVFYAeVQ/VFIyOTlh7aOWNVsNsblAf4+aTflQBL9kscK4Vg4RkpvDxoEdMf7plLWPWzZ+7sIJoIK1o8IdzI4QJMb1NPSoQK98CFTEYDH+HnPR5VaI1Lpupn24r+DkJFDhZtrJjopSzYEK3v8XARXMSRnHk1D0nH0rplJgkHmQP5Sn4WtJVIWOighUEIQfH7cEVOBNcefmh5aR5JYHTnwQSGGkxL8RrNFzDAlLVkbJMSDB8NWLBnQOECQQEO0cHAio2Nzd84KBjGWdIQSLQ11IOQCbjPYBdVsEHwsd5ip+OPBATB09JngtEmoYLbCGFG+rOBl/l7ZHngfM37Z1CH77BP6x08AZ9RGoiIXvxxWhkkCFAneAjsAajcFEBAYj+4jxih1i+vtMVklnvlKzK88+bxevPm3ZYsH26wdWh32WSdutT29pnOfm5pQ8kQwsLy3a6v3btrH4yLowGgK794uACl2/2NYeWKmGmazSPmZ+xDmTPEP6CaAiBqbD3+tZqusdDFBkUr1jm5+dFAPo4tk5O7Mwb4uPHtnG+roSwcmJSe179x88lBHXyOiYEpO9w0N756fvWrFUVmK3tXcQ2IgkR/FqYkfFEKhIPqsIVDBndncwPIW5G0EK0VkeC3BoXv2cjorkeoprITk+yTH9eeDD6XP53y9Q4R1C4i9Hk+Qon/NzgIooWcJeVxmr2e//g//ORufOWQ85wl7fGttb9s//n//L9jeWdC4lQZvkfndiviQMkVVkUIE5mGsHCbUvAir4vtahnhtnuAMLJ8eKdAeDcJ93nFtdui0DUNHtU9zmdUgkvOPL5wFdazA0h4Xg5OuSEPv5D8utJaACsMb3r2RHxRDoCcOtvSiV7tjXv/41m5mYs5vvfWC5dMcmRnIGX+7mZ4+s18va+ZlJuzQ3ZdVywdq9vm3s79nm9pYKVZznFEUoZjAn6fyj+MIYUAY4bDRsc3tfxUsKwtGMnDU+7Pv7xUAFEpRJICGZBAHk8t6nO/N0nwmNd9iCvq8E0Eo4+PAqkmuGp8XMFCtZQHNS4sg7Kvw5D9dqfKnOMcUvnxNDoEK7jzXrSD121cU6f2bBfud3/xvLFUq2sbWvfZSOtAhU0Mn559/7C7t7+7aYeWPjI/IS4+xFPhNWGUAFBUZY8SmIFO22HdWPbHV11e7cviWyQ6frBbwIRsSkfDj/vagT10n8fhxP5lU8N2KCz9exuJ6Ua0p+f/j6Tuvj9VWADR/8/WnQKQkwnN57fh5QkQSik/u97/nDthkl7VFGUKm2z5HH7Yect/xtsVTQWci1MeYXLlzQemzh0xa6dehCVsxPrEKcHYolgh2DjB+sbdj6kF6Q+UzuRREUjWMan8faGh51/hEB2njmx9+JccaJfSFMRnVyt5q2vrGmecX9iPxAJ3XoqMC4nbhlvjBlxULF3vvZh5bNFRWH41H3/7P3pk+Sntd15819q33fesXSjcYOkDBAUiRFi5YtW6GxFIrwTMR8mT/N4U+OmBjHjBfK1i6RIgWQ2BsN9N61dm1ZlZWVWblP/M59nqy3Ct0AJc0HcwKFQHR3VVbm+z7vs9x7zrnnvnDjuubdz376t/YG6ux+355//pp9+OFHivfv3btvzz13TQA4AMHu7r6qBSAFnnsGUc2xXb64LGtVxB3N+onESsS+65urVijl7fXXX7Gx8YregzPw4LBuDx6sSdlNnzFEUWMTE/bstedsa/Wh3bl728bHJmxl5YLOXAeovGfK3NJS6CsF0JK2evXAhRqFnBVHSsMzp7q3q0bxbgPXEzlxdHgkYANwu1o9sPGpCXv2mau2sfrAum2U8wB5XWu2utrf8nmsdl1lL/UzhDPgbL9nW9uPrUpFwvS0XbpyRRXeW48fa65NTU5as92yO5/dterump2guC46EXn12WdVjTE9MyO7w2a9IVFXr+PK7F4/bdmcV0kgGiKvUkWiSAssLNxmDCUw+UO701OVCuCyV5l6fKUm8AjmVIlxLNBZIHwgxj/44AM9zxdeeMHm5+bsqF6zRw8eSVDG2rh8+bJdu3ZNFRFr6+v26OFDVZhcvnzV7t97YPt7VeWbiOcAQukHWBkpOViXSgkk5Ys/WTvcKzmbnmewDmWdxRzPz460qszZ/1Tdn0lbuZhXfJbPeV5BXgtphA2smqMKcPc1xL1jScga2js4tOOTlgPwoUpCr0XwJFAeq2bOYa/CJa9wgoRcMiOBnOfQbqPLnHEhlOfNqtwO+57IoXbHWs3wDAd9K5QA9ZsicrLZgQ16J/ajH75lVy4u2KDrz29nt24P7m9KFcy+LzV0q2N37twTUcCaZnyp9FpZXtJav//goeZz4xiSpGxjY2V74YVrdnJctwyNbwddO2nUrVIs2tTkmM4NBHc//fkHtlc/sRSAvg5Ot46W3SzKaTCLYPniOTqVFi0RBFJwdzsC2KPdNT9X01166iG2CvbVkCyME9+HBObvEtjJds/FdggOGTPG3M+ElJwFAPu9gsNV4JyvEoSFs8UJAI+bk+dZtDyOCvChDYyWQQCz9Z4EoIjR0jY/O2Xj5YLlBj27enHZ+p227e5W7ahet0arbfVmW5X2kNX9tIviwDCIdRgLYh/2AVUxUFWT9vtmLxOWE+2Cg3WOzlhZ7nhVlu479B3l/GGeoQD3cU1bqtexpbGcvfXqC5ZHI+Pm2vbuB5/Z/nHPylPzVm91RZjUDva1/lRdGogO1gL7sI+pu09AWkUBo9sU5kR4xYqL6BKQtF7kuRK3sHZx/6BKHVcLyMtCLmMTI2WdJawXzgbmVr1xYpefedb2qgg0qDCG3Bmob9fJSUNn1OuvvCzb0b/9259Z9bBmaUBnzk/2uLDXa1FH4V0QM3plCv1gHZc6PReD1VGSqBjmk97wUPGNxFLuNuJEBWOC2IFKLyc/sB5PY3Paa9uzVy9Z56Rhtf19kdhU2+WKZeE1XezFxyrCjEqlgjAxbD1zmbyEx+SOzOPK6IgV8hkrFXKqeIIEwZb18eMda5x0bXxyxrZ3tmyvuqu1QXw3NTVtzz73nCrrAN63d3Zlf0vFDmNNdY/3iHWRSD7r+xPPM7oxsL8pLkPIi3V16KfnElH/EkkYnDp873ZxlY8VZ64LmJNVt+djt9Nn4OXHOJhYt2MjpaLduP6c1aoHtra+4WQjRFZ3YBks3zsdWbNDyjBHOP8qoWJpd29Pe6yqkrJZVRdTqcZZzM+E0eQLcigplyHo6etJ420qk+rCa0QkF9mvXUD2jfXTl6Lub77x/4cRWOh5kEvQxMKF7VQAKAU/h7n7uXH4quG1DaxUqXh5cVBHc+iMj45LaaP+DCo/92abbMoc8iRIBCgtsYIpVTtQeUDwo3ImSsbkae+EB4cHh5vsdtTc2g9jAm0UzysrK1LuOPFwYqUizbgd2GBBt5pNAdQEPt5Mx218CMyx3HFA0RMyNgbY3PJISUw0wS5+voVcwfb2qra3vy9/OcogCUqlspD/OwywkxKMVWzYWz860mdDBACAsFGi3FyYXwiBZ1rgIeXjMKoqdQv+u7wXgQSBLMHv5OSElymGAFTkDUlnyuxHP/qeHdWqOvxnp2fs53/3UxEhBHx99QjxXg4EY95oKCOlbz7PPXYUONL4p9Ud2L1H63bc4GBQ4ahKHwGXAbVRkXB/UWbtjYi8B4F6deDvTQUOZAXPnUS209JmSvKCpz4KPHpUtLttmz5XURGB6EhUsK4iERGJCrfoonzXg2yBBMIHnQH38fGGqwTOzKt6rapno2cxkrR+mnBiJPgvR+sn5kkkKmKQyPyICTVWJyIcgs8J8ylJVJyqHE7VjXwvEhVcJ2ouL12knLVlJZRF1rd7t25ahgTiXEUFa8DtyvweBR4FlY+ICuzGAmDSS7nyEusnEX6ZrBRXX9y7Z5u7ewpChoAOiU2weHHPCfe4dgVuUGNLmQ1U4SDRUM0hwAznFwJLTzCjytNLb92mpZ9C1cQz6ooY63aCYkgK0KwCoeHYJgD8U+DIm2JHECQ+kyQ4FMfcS7RJKhwQ5D1QkSaJjEImb6XxSXvu5Vdt+fJVG2TSsn6COCxlc/bg/gPN2aWlJZtAFUgz7bVV21m7b7trq9aB2PRZ99SKCo+M/FkpUIrq1nPkVRLkSZ4jcTzCEA9/lCQHlJhAHvEi9kfKorNpW16as2cvr9hzz1yR3conH3+iBB0LqJmZGZXuP1rbFGCCKuPh6pp9cvOm9gCWDWs/pMOnTb+lHAe++DJRwWuZn1RmkSQARpDQRLKKP12V5oBecn1o/w1ExfCez1l+JcclaRfypLGLgeR5sPI8kHj+zD7/cyzsaFAfE4ivsn4aAs8h2dDjfgpREe+R+zjdr3pWGi3b7//xv7OppcvWT+dl6bW7sWb/z3/8j3a0vxlsb0IPh1874PDKsbhPJsdLhKNIA08WY6WKAEb2jLT3XUpK9f3apSvVemTOcTahro97SHBtC+A3wBeJ9tdXVDC9lByjWmy5OlL16dpTvCJJ43peUR8qNvrWsumpCSvnxyzTG9jEaM5Gyilr9sxeePUd+/jjm9bYeWxXF6dtfKRs3VTa9uo1297dVUUFnzk1jod/Xslcq3PiIC0WlcQBJy3bPzjS9xzYDwtaIK+TxCTwrMmv6lEBef40osIJXAeNk/uhplX8OA6yYDflikl62vhzjF9x3/PPIV7yCjvvF+OJmffoYjxdVKIyEOaEfh6t+VA6exVbJCriexP3yQ84n7GLVy7Zv/q9f6PEnYoK1OCAhcRyJWwl+wN797137aMPPhDIOTXnhCnAYqlYtNEKAotxJ8ZFrlPF2rPm8bES2UcPHtre/q6d9Fp+yjxhD02C22fnuVsDxZL+82dGQinzpfnlRNApsaa9NywIVbgEEP382fW1yzM8zHjNZ/ee+HlRMXlqfzhUCUo1GC31XDnrFx/ZDN8nkkl1Oj1QIiv7mDSWoBV79tlnBYKcyHEnVF1h7wFgHPrAKC4m1glVzHwESXEPkDSHqjs0I4+VT2EvSc5j/r63txfERT63Y5+K5HNL/k5yrXMvsojtdkRUeIwM6OAkCc/Xq8DdvmU2M2GZVME+/+KO7Ht4HeDA62++KjXoz3/xd/bSiy+p4eXLL71sn9363CqVEfv0k09EXLBnYe3BF8ukXj+0V1++YYVcygbdlvXabXv11ddt/eGqPXxA5QVg/qaNjFXsne9828bGKsoPsDKjouLW53cFjlJRwWvJB5555qp1s2aHj7cEGnnVuY+Ngy6+D8vSpFqT0vrOF7d9L89kbGllSeuL/GTQ7UlEhGjs1q1binnZxwB5IAUQZ1H5/ML156xRO5DYiDHjmD+qn9gglZUNm6z0hkQFtpxuM0sVJmta4F7KXN2+tCiBEkII8pRzzqTnAAAgAElEQVTlhTmBk7e/+MLu3t+wbIGqIyrRRwU+Ly4tW6VYEfkopTbaikFGDUEBdbG7EU2dzkr4gvCN6yFvo3KBPRkQfnp6xs+C0J+Na0JMFucr77W4sKDPJt9kjO4Gey4uHhJAytQipBZgOTkjJFjTLlxYUR7D7+7tYm87LivTVtOV2Zpvg57NzE7bxMSYi9o6bYOEA5DliziHuUTeNjU9ZeVSxfb294b7rqw5up6XAGaRC7HeeG8IXfJW4nmezUgxr2oEgNvxsVHZlZCrMQYA/pw7ldExO6gd2T7V+9iUKB53yy3yQc5UAC7fGvxsofcPlntedTEukBfCEbCdfIHcempySoQQYjPGBDDSbbgyqsTttgcikdqAYuWCVQ+I+YhHuY+2/e7vvGWXV2as1TwUuJnLjdju7rGq6lh3PD9y8NrhkVUqo8IFtP/niFfczhd8obpftd29qnLfSFBC3oyPVmx7a8MqpbyA5LGRsg16zKOe/dXPPrADgHDA2CAWEtkV8At2cap4tHNKQJFVBTl5LPfPehEQKosVJ3XYV/iT6hHmJeuB8Yp/Z06KBI4WmMH6mvXM3hOrU9n6mV+csbweABMCgHuPFlqcVV6h4PkT783859l5XuOgLNZMLiTlfHeRjLAY5cAD5X15iIT0wEYLGcsOeqq+RtQ2Nlayyakpm1tctvc/+lRKdlU6hKqPkdFRfSbrkLz+0dpaEJO5dQ7PjHxJtlasJ8i7SkXiTXfjaIvwgNQGL5JKPgjtmOvYJw1z+3bTlkbS9uK1KzQLsAr2SqURe++jW7bf6Fl+bNoO6t4PE8U6QDj7IfEM+wjPQZVauIKwJqhmClalYDCqbCHvCPZBnCOyXA0kXVTncyZxncxFrg+Bow06trK0YJlB38oAwbL8OrGd3ap1+iarp/IIa7AuMStzOpOjCrcjISzoxEs3btjC3Lz99Kc/E6FB5UETIWuwMBqWGYd8FfwhEmhcNzgL+4qwDVl7ncbC5/OpSIYxt3lOxIbez82JCo9bVFOrHI2KfPaXXNrswvKCNY5r1jo+tlQKW3BI7Izlitizd0BTVHkhciqIjRHfkl9DwjPu0zPT6ovabh7b0vyMFXOOG3Q6faseHlmpMmrdnguEWQdffHFbc39+YUnPlzOFShnGgOdJ9RykxebWlgh31p0Kr7XFIXYMsY6asAarJ8XhTlrJ2inY9fJatyBzVwv14A023px1ggLP9R9MVlacjeucqIBcNnDNkYpdf/45Vd5gAyZVNnZcllavCvbllcV529/f096Pqwn7GWSPxM6c182GxkL29bh/jI7IUj7mZ2BF46qSa/qzDRZ9IjFCFbMTb2Bd2LkvvHWaFXxtVPrNC74Zgf/5R2D0qC7wlAVAgMLiYDNSQKsGlj39HA9/yvIBg6Vskb+jA1SADBykspMpEXin5JPJ4js8qnmJKL7WTWx13CaJzYgvHYqBmWdTJsgkmGST4s+YeLk3f1YlvBwoChQoVWw0VN5OUsFGxO/E6xa7n0krGBHLH8rV/X490eLwIuCSOjl4JKtMUMy8+/rB9qq0LNHUmA2Bw4lNzhvVjmjTgLhABQ/Y+Sf/43/YKy+/LHsZSrXn5+al5uF3Z6Zm7O69+wqSUf1wDwSsXAPMqsiFcFB1sWIJVlt4lvN3CI5UikAna/Xakb+217W56Rm7cvmSPKRROOPDysGopNqCb2i/I3UFSk5PFDLWwy4o589lZKQiT0bso1CYENTpegSQ9+SdyqZbLONr6hY/VErwu4MM1SsAC57scJ0803rjWJ4qEBWTyxdC+avPMwEoAcyMQDMHSlIdz7yThVCSqAgHvB/SXsGiAM+wMehY/bCqw109KkbGHVQKPSoUEKrhZNZypYKCN66DZ8g1xGBKXocBQBJREQJHV3NRcnxaUSFg6ZwtBN+L95QkKrg+rJ/KhZyN5HP28PYtax4eGnpklWeHe/NKGIIzL6NXGTNEHgop7NqyoWcFzaAGvg4JSlV2mctbq9dVj4rN3arbLaEKVjk4MIcDkFF9EAHJCBY4mOBkQlTJu/VEBNXSquLw3wtVBIqnHJjuB097WXE1m5pPw1JVSNDYtDdRcaAgJADWcdyjMtYTwlMbjDjeDqi5Kiz6TEZQRAd78LPG+mlkcsquvfqGzS2jYE9ZvdmwY9RZ+YKtra7Z7u6uiFCSbNS9a6uPbG/9oe1trImo+LqKCge1XEkeKY0IaD0JVNOcTChz42uTRIUL4qNq2BVUqnKBEJEkHQKta8VCxpbmp+3SyrKtra3bzuPHduXyZVtE3Tg9bQ/X1u3m519YrlDQ88cPllJk5ooHQAmwDMW45jJ/9myQPvXYTwJs7GXlkYrm3VGNSiq3lBlW1sgPNMyHxLPTWAybPocGt/9QooLZmSBBngRkJgPQJAgWT+YzAKaSSRrauw2dZn+I+J7Wo2KYMES88ClERQTjzsxlSnuLBfuDP/5fbfbSs6qoICFau3vHfvKf/i+rVx9rL3vitSaU9F++Lwegk0TF6RyEkTztf5IkKtwuisT5bEWYvz84uSfEsgfiPG80/dzEJiBzqgJk/vu686SbHhWRcBzO7/CsGVeAAgHKJONgYsnqkFPXp2EsoLkTfGd7vaYqNnKpoi3NzNv8dMWK+b41LWs//td/bD//6d/bZ7/8hV2dn7D5uWmzbF5ExV5137axJMIOZ2LSfdHbbaluOc/YO+FMWB/Vg7qAmfNERdznmPNKFFJne+skoz/I2uRzPAtSu3IznmPJfSLR1kBExWnVGkTFuRQqjJvP3Z6VChn1Ioqe7U5UMLeDnVYgKvBbFlERLKA4Y3l+TqoxJwIxjdq+C3CIaCVr1168br/9o99R08CdPapMUTVTMZG3cqEkS5nqwYHdvX3H1jZWKbSRIh0QBXC1UqrY5Pi4xp7YBSvQ2sGhALWjWk2kMYBtDwuTBOGbvOvze2okGfzMcp/mSC7E8Y3nxvB3Q/Lrx2OohJOFRqJaJVouhAqxeA3JPWf4u08J+zk7k2frWfLklBg5v56136vXkcdw3jdIJ8cTKypOP8PzZhJ3YnFXS+flyQ95cdJzyyhVLwHEnJxI6KG4mFgcFXKoilLvGOL/qAgl9gkWmVxX3GvOExXYGyD+iFUUsQoijlUcv+Tcj88lnuHEdTs7j70yC8uqUHWrngCq6IYcy9nl0WURcB988LGNjU4IeOTzXrhxTTZNd+7csddff105x+TktIh7+ifs7OzZiy+9pPv++KNPNG/q9ZoVS1l7841X7Przz2htr966ZRur63bl0lUrVyr2ePux7R/sW6vbtLfeflO2QCj7J6dmrHpwZL/61Udm6ZzNzs4J9J9bnLdLF5ZlZZavoFjNWB+7nzyCLLOTo7pELO+//6HduvWF9psbL75km/JFP9R1QzwszM3Z+++/LwX8izdu2KvvvGPv/uVf2YcfvG/PPfesqkTW1tYkaLp85ZItzs/azuaGtVsNzxMsZUf1lq1tbNnYxJTW28WLF7Rub33+mSpmEIFdfeaK/eLvfm6lsje6pzIH+wpiCSylus2m3b19W/vQS2++abc/u2nrm4+tRqVBGutg+iaklE/yGlntFEqWzuW910G5POyx4K+vuzIW+xViiLSJUAC8BoyXlWgbEhkQzslsxfGKsb3iHMsm0gHFpZYSaUDDVM23PjZARbe4QqTWassDXNbGUxOqAJ+ZmbNOyytc9nb3df0A8A5ap5UrMk4A+Oxt+7t7WifkPFTnYbNFDxhEeFJzh7wXK1HvYVFQ/yTAKsgHNUSlgWqtpnuFTGGN4XPf73dsampCQHx1/0DPe2py2mZm52x7d09EBYQV9qvkMqiGuY6rl68oryG3ZUzJw2bnZg3wlnXIvgOhvAMpMzainJV/a71nsiJgtBsNTLko18d41CBJUqHiIogQwf2OagdWLDC+J/a7v/OOrSxMmvUalk0PrH7UtsmpRc3dtdV1gbr0d+R5qjJdHvve+4p9mufXanftoFZTL0FU1dG+D6AdMPTwYN8mRis624jH6ZfX6gzsb37+gR3TD6SbUs8Fzy29f4NAPOxcZU2KxVrDbaGC1RN/xkpXxil6+isPpSqAChJ6GZB3oTTH7hmAu+v9ExtNyH2zUiHruIjuy6sVyIvJFd1epqtKLM3hoYOA2/fFngoMvecx3p8N1TWEsp8XEB15gZwsEOduPS4T9Nw3t8/p9ezG88/K+um5yyt2XDsQ+b+zvavzGlKD36c6Z3p2xsYnp2VPx/8AyXLJ6HasMjoa7tHFFIwfGA8ThHXq5BJEFZ+btV7bba9E+DCvj+i542cx48XHkmPzlRl0bGEkY7/93W9bPm0i5dY2tu1Xn3xuJ4OCpUtjVmt0FIOxt/Y6blcN+ctYgOvsY+EJiB2+qO6nT4PbUmW0HjjryNv1zMLaZz8jLlKfVapGOl1bXFy0o9qh9dsnlk71bX52RhUVL71wXc/m1mefqXKs3gQzSavHJ4D0SQPSs2TNFs8E0swrKt5+69sSY/z857/QWs0WeA2iUd9/nER0FsXzfciJWPXEM0Dk66Xt6i4ahH0xfom5x5nYPtgZCdQnH5a4yH9fRIVYG2WobqdFX5xKya5cvmDrj1atdtRQ1THimyJnVCZlrQ7jS2LP7Ynq8Jhh4PZZ5A0j5Yp6eVAZ02nU7e233rRSgYoCRC1FERGQkfSMajRb9ujRqkTAV595xq2QJE427f/Ys3nfkaxdvXpVGNLGxoZ6PBwe1ATsY88H6RMrK1xohXCTOB5sxfvUsf5EXoceFNpzqNwLdveKDVMuJnViy0nniEl9OZRjdvetyHv3uzYzMW7Xn3/WHm9u2vr6phyZO+qvl1NNM2t9anJUxCL5MVV3zEUs1NhzdnZ3RPwSS4G7gR2ShxCT8G/OCeInCEJwRGE/Ic7nPKCKWT1WwKwy7orxDVHxlAD8m2//5o7A1WLJDjmcgqWN++J5Yxk2dZJINgz5ATYaCqYgC/g5Fk4EGST7bPgERFLeB6U7wRIqGZJ8Dg3KxCCGCcZh5QkaOdxgqt1T3ntOwLry2fGQJkEqVcryhoV1JJhjmyVwUJnwCb6HaalB1JxGqhtAdW++iaoLBQ9MJaA998IiJxCgxBGlN4A+myPXwIbJNToo7R7NXGe74707uC42lLHRcR04BJxUohBAMH737t9XECvAlUNayn1vSMjhTd+LC8sXbH19TQck30OZkMu7cgIigEOVsefAI1FoNk5EGpB483p89fDfVQAVSpEVyGVzKsteW1+z4+OWvHkJsF194SWH6QHPltem1dgJDX5H/gEoRNNWIZDi+RfdR5371TVJPQR5YwIh1CxZ5XmeSKMoxd+bP6mM4TlyYGBrhdJAiUavYxPLK0Mv2UhUxMQ1Jr9PIiq8/NYTmfjzJPMtQkBBU1/j9jSiolIZ8+oBPEQBuQt5m5zyHhaRqIjXc56oUFk1SRTBZCAqYhKeBJyTf4/3NCQqsl5RAZnD4f785Qt259NP7Pann1gBYiJPabArB6MCkX9HiynmLgQiRAWl/9Hzs9XDL7Zjg46DwwRS7UFfRMXOwZFsCCKIAVkh9bczB09UrA4BAzXXO/Uzj0pplJ5UTfjrHDwhGPJmcMx994MChAIEiQmfgFBZu5xWVJwF7vy6IlERA7Ek6HwanLlKMypn4+/o/rPZ074eubwV8yUbm561F15/wyZm562HJVybBo91K+Xztr21rWCeJB2ygrFcffTQiYrNdes2TywrXkDOl09spq3xBZELqnTZ2jyBkEmeGP84ooKAk71O7cE01iS22AUI6A0gEmWm7NcEMKubm7ZfO/R9QCS0+3q6hyeP8LSiwm1m/HkKKMt4b45IFMV5JIV02RueoiAjUHQ7mVMrliQJOQT2wryL4ODXgXwRUE+OmwL9JzQpP63IOSW24u8lwcoY8MefSX9EgKv5O/D+S08hKpLXG/smRGJDkH3C+gmwMKpjkp/Pe2TzGfvDf/e/2+LVa05U9Af28Xvv2p/9l/9sreM9JfDx6/waeVrUwTPjgSbBw7iW9Sw09qdrLIKLIr+wn0o8u1MgFlmSzxMHnbrWOoZ8pAw79E0hfQtWcd7jxIlOzirOUO2TQQ3n1gbeNBKyVyXYygGo5nNggRNF/VjCVyQdPbnzxDyTAVTvWrkwZguTMzYzWbKJsYJlx2bsR//yf7FfvfeB/c2f/BdbnijaxeUFS+VytlOr2c7enq09WpVt4mToZcW9ADzKD7pUsnQ6Z8cnJ7Z/UFfyE/crXxin9m6RqDhdP+efDCDOqVUO16798fTOhkBuXFfDH4VnFT8zEhUikH0CnxmfOPfLhYwtzIwpiYnNkdWDgASd/kiwMFLq0ZPCba2wg4KY6Pb9zPd5cUpUaPzxt+91pB58+ztv2xvf+rb87nd2D7wStFySbU4pX9K+xDwhETs4PLDH21sCRam0oOKiQjzXatv+3rY1Tw41r4glGZt26JNFb6VBruDXl6isiTcd57X/O1SNSFjgooHYePlJvxt/hz/j3PK9Kjav9rF1giDsh+eIiuHPE2T709bleaIi+TrIo2QZ0+l9AWK4z3QkKrx6kS+3ewjsv/4e+7n4ug1+1RkawRaHRMUzzzwj8KbVd0u22FOHZHpIVEAeJogKns2QqCC2/jqiIjT2/iqiIjl28YwYnhuhJ4hX0g3UsySbc4HE04iKucyEFQoj9uFHN2Uphoqd3nbXb1wTGXr/3j2NsfooUbVwTLWA293yWu3HWSwuqMTGFzpnK8vz9tL151T5uvd4y25/9rnV60014SbGz5dyNkgP7LXXX7bJiYrsjLAWbbX7WhNYaNDAlt5PiJEmx7GZ8wbnaQCaVNp2tx7L2ojYHrB7fX3Ldvf21cQaf37yLHITRFcjlRF5Wj98+NAWFxaVq3Et/Lm9s20T4whyUlJkImJaubCs+3/vb38qOxNAYkiCTj9la5s73qNCwrSMFM31Rs3aPSo0swK3Z6em7JNPP7aD/arAFoAXNbjO5W1xccEuX7rs5MdgYPuQkvcfymYUJe31Gy/a1sZjAdwIajyfo5I5ZWkq6GnczlrHaharXXr5ySo4VmB63sF9A/B6/OtxsKIsKWgF4QXgzM8fNbTGZpbcJIiO+HwAZXIkEZidtkg4VVZb3/NU+oTQaLzjDetlMRZ87ckLqdzHpihfcFU4ANL42LgEcwBtbiPiinmWJX8y//Fj59zrBSumaJum/iq5nCrMqKCAxGHcy4Wicr5+yq9flkzpjO3v7MvPHWCPa6VvAhV/osA576kcaHVsYWFeaxXAOlr4MRZcD/kN48xcozcfVocCxaU4piG25+qqiMaBIKjNY0WVjhzurVSy/b195Y9UTqStLbunH//oHVucHbWMoSqnopo8mlg+a9uPt0OPiLwqG1BlA2Qy96JNM9Uz/UHGNh5va41iUTpsXN3tav006YvYbtnUxLia2nbbfWt1+/Y3f/e+tbCB6gJ4eswFtkAuyywBLBWQL2GTzzHwC1fke6Nmxx0AsMsOIHOGhV4ijDljjFUY+b7EBcIb/Lxkv+R5sRaivZPi1hCLUVFCHMHaEfkWgHSIFglhQk8Mvy4/f6MFlCqHwq4PzkA/QMWUsuJ0iz+d5xIDQQ5m1Og31WvbpYUZW5ybUSUkRAPkz9Z21Q5qB+q1wPt2un3ZH4OpKJ/q9SQSOD5pKJ6HEPR1Q+VQWRjMyGglWEE1VEFFlQxrEiEr60KCRUieYMHEtUa7NBF0rWObLWbsR997w5pHNZudnrKD2rF9cPOOHdKrvTRm/XRB5EmxCP4AaTnQ3FNFKe9XPw5WyS6mjP0IWG/eWNpFFwKxWcNt+uRQUURPSvYIH0dyPp4p+36F/cNcNU/FAddNj6LHj7dVFYS1TzqHvRjnb0YCXNkMUpGTT4tkZKJ968039LPPb93WWoUcYrwF7hO9PkH2zrMn72D8uS7Pt/gYj+mT8U4UM8ZcOcYTAtl1zrGWuhonwHhpg5QvqsuEKgLomzNSytvVKxcllD08Qvzb1npqkUNmTPZuKbk1eNSZUQ9Mj9O0BmCU+wMbLZVsZmLMpkYrVqGSJ206Iz1zTNnYxJisw1XZEAgOqjG0bWov4Az2fjvrG+sioHh/eu4szM8rFt1Y29D8ZW/DlhAhNLZaEEgSE2FvFXrDQHpwxaxFrWP1yeRaPSdX3BeICvaYGCvGXDOZ657Gat6rr4STSq9r0xNj9sLzz9vWxpptbW3LSg07deZIW9VNKbt8cVE9Ow4PqCKj34+LoCW4HvRVPcbcBJ+E8CJm3nq8rXXG9YOfUVFBDAAGyDixHxDDQVhSWURMz3VDOH9DVDwtAv/m+7+xIzDPiR4AKK+KKJ8Gg15J6g28xNh5aT6LAX9n2cKoWbM3klJjMwDI0LQaMB/1Zu2orvGhIYynk95UjN1DFlNZT7wovyNohBSQni02mkLhdFR3wxWBaq4EV+NRbTiUixak9mPzl1KhRUDgdlICs0SA8N7erIdANDZSUhNtJUSmoJBDR8oHmEoyeUpFqZYLZAqs/Qy9GmRb5b6iCnYyaQF2BCoCTAFnBAq6byPBw9AHWkmUM+YcqBwGlOnDFkPIyA4qNF/2cnAOxKbeX2NFuSr0dR9lQU7lvvTmgMEXAYPNjhh4FPqUz6NaCUphqhLky0dDoqyACQ4KNRCl4gXyqNm0UYLC1okqYgAOSBoU+BOGcv16Tl7JgEc5G3u7TwDtzdYZdthwGqRBMmABxWsjURF7IUgBGpT00V/ySUQF18t48VyjMugsUeEbOGoIJyoOXIGiMk0apHtgWS6P6r7pPaJgPp9RSTQ/53DUWAVlpaysgv0RAS8BhKyfCCaBD4JiXAc4pE9QYgv8j77WATQWUUFimPUGn6lUT4H3MxdXbOPBPfvgF7+wvBTIDurFsYhAIgm0FN9S6/AMCcYg3UK5fK+l+x7gj0j5LwqOTtvuPHxg1aMTG8gj14MdgiFfix4AhVxnCMjEoIifqz201pwTWREwYb7208EvMrzO79nnuXzSQzJAo0D323SVPpMjemsPg4agsk6SFDFYU1ARAoxIDPE99YeRVYCTiBHw4O9R1SOSlH4quaJNLy7b9ddet/L4lLVVCdRRv5VcKm2H1UOpyai4mgtExdrDh7a78dD2ISpOTlTxEokK76cb4ScHjhxEPbV++iqiwvVRp1UBQ4UNc+eswDahJo8VFbEXhs8596N3Wx6ICuaBSECA91Cd1MYnXz0zvGmzKA6CRtm/UIjjIaUAP4iKkKjp/dNeeh7JIs1Jev6gcMqj8Dp2VaOI3eh/7+/Ba2XvQ3VSbNQc9uSnWbrEA9V1+mcbScd5y3mg5x0AgrOgpb/D+WDzK4mKMwkiYqKnExVxng0rKkIj4vjYzjfTZg5GUjbuC1wv1njf//Hv2cT8BSXZ6cHAPv/gffv0/fes3Tx8KlFx/l7PqrPDvJT9U7R38rNAz15/OlHgBApJqKvxKL+W0U0CeI3nbZKoIAnC+olETOeyCLloO+P9bJy8dJs0gaihMi3ev0QFPD+2gwAEgzDEZ8Z7RkVZcv0PSSIUYhn64PQMA71nL16xa89etFb7yCaXr9pb3/mhvf+r9+3P//P/rYqK5YVpnXHbhzV5rdMQF1u0ydExnaEAaMfNYymxox0J/ul71aMnEBW+Hyqx/CdWVIgjEClwbtHrMQYwOpA+Hj+ECjZtsqfZbmzCyKjPTo7YlZXZUDXnMDtnB88NQEbVogJ1OvKIbwOyqPkgMZmr0Pyz/bqG5zNiAJRilaL9zr/4Hbt85Rlrd/q2vVsV2CevdZo35/Azxo7TJIQhrkH9iPKMykRsBna3t62L4hFv47IDCV4i4IQoMeZB/djaKa++i+RvJA0C2za0v4rfV5PKYEvqdhpOnCYJzPPrh9gzNpbWWkqACF9aa8kfho3qlNB7eipwnqg4fV9ihUTpUKIyk3dDuXhaUeGgn3+FigpWbCBs4xqL57lXoKaHRAXnoKyf8FX3Bkq+8qjIhMgKFRUS8OBlzZkaiBqJDTrudc+6jGszntfx/HXyw/cWrDkAdGMlGa+Jgos4ZvH34x4WxyWe4cy/1dWHikOTVc1eUYEy28G1peK8pSxnX3xxV01VubNG89hee/2VYNE6sK3Nx/LNBizEpgThEqRdHD9V5Kbo3ZC1XD6lxr1vvvayTYxV7PbNz1QB9Hhr2x5v7VihVLRsPqvY941vvSqffol68OIvlC1bGguCjIy1UHD32rIVgTxph34RY2Pjdu/OXVX0jk/N2Pbmlm1tbguUWV1bV38GJ2SDACycp9ijvfjiiyIBGRPyIgBxnhsAB6QC+/G155+zxYVZq+7tSH0uxXFpxB48XLc791dFVAByLMzPSaxF7K6q9lJBAq7FhTnZVXFfVEbt7+7q75z7xBjMnYsrF2WFMjI+bkfHTVvb3BJQPDo64c/g+EREhQAymgu3Y3Nh5pB8c7W/Sn1OD0JZezhJLXtR9gIawKJ+D3kWz0zAqYRmPk9VCYcSHCFXojqKn3VksYsquyN7DQR3yjHUr8GrDAFpyWWbNPwGjLSU1PE0d4aAZQ1CUiD6IGeDhGA9kZNFZTb5I7EoBBM9wgBGOVtkqaNKtSBykX0i1QOAq249TI8RqidQkPAZmQJDExpAp7OqQOOey5URB0g7bTsktyZvC37rIisg1ROV3qfNx8k78OFnjFoSmDB+jG95pKzqIvZgCQNLTnBDirEv8L+aUyNGUx5M4+6W+kd0yF3ZZ2xgv/dvfmBLc+OW6jTMelRiEGuSP+ft8camGvDSB4S9MNr0uMWRj02+WFYDZRToAvPzuCo40Kpzodu1x1sbduXiigR1KLk5uOonbfvzv/lA+WdngCCCankA924Q1aGo92tXLCIBhRMk8WyI+xS5dLTCjv0C6XsSiW9+RhUOYx33W4+zsh7r0DBboCvPDisgr6KQQEAAI71MXBnxYpwAACAASURBVOBBPyz6VUIieFWQxxQuyAM78Ngq9qjgZ+Alyr8h8WTTDVXlhB3YA2IhsADGKI8Yjj6IA6rSdiybJ14v2PKlC/b+Bx+L6IIkbXVQsoO/eNNv5jUWzpCP6kMQro21E8l8CTgldHQyHXyBeJCcmn2JigfhEEFP4fGJW3qr+faga5dmxuydN66rXwWivZ39mn342V1rDArW7GUslS96zptjrTKWHa1J9h7eWGQkWA45D+4YhZLGZmjRyHgFuynZl8tiJ+RGQ1tmyBdfW+wTAOzkqpViQbZP7IPMPX6XPgrsyVRHzMxh5d1SXMNz4yxKZRE7NrSGr165othnd2fPGz8DhgeQ3r2LgjtAyMOZh6wz9aYIeZvOf2I3iUG9MjkKGiKhlcyXY+zC81eVAHODViHC2tzCUva8clRAlGUisThPiN+0ZgD7qfJLZyRWlf1Tn/lJfCA0IFTh08sVXAgbpIFlBwMr5/M2WszZxGhJ/TfZL0fGRjXPqa4BQ1xeWrb96oFVq4ciL8YmpjUHdc6BMdH/EiKsUhGmAhG8sb4hyzMqEajgz6Rzei9mPeIASG9IJM4eqs8gtyAuHD/wYE69Z0IFnjcy9/M6hZBX/WV93/T4I2ae5213A1GRz9qg21FFxY1rz6sHxerqujAWKgap8OqDz5SKtrw4a1tb61pD6hMiOzm38+Nre3tb+z1rYnxiXN/f2NhSRYX2iJOW4gMssNiPsWkjrmXOEpOBw+ksTrsg5Rui4ukx+Dc/+Q0dgWn56+UVsKuoPJMWWM/SpsSPjU8+gCFQ4TYVfKECqZS1OAgUCWpYVBy2TjKgpKa8rm3FcsUrHdIpkQC+cYRGpAKZTN9nIyawiGSEEiGXEGoj5H3jZ3tjGYAqDsqgCAm++1QYUP0RiQBtDATBIVh1cMxVoHHjcmQ1ADSh54TUKGn3KE3nfTPjEOEgUrDbbmlzA9hUlYNKIz3AIMDh9d6k3MsUdairssFBVP/yw4ODYHgEBaCRZMPZU1c9COAB8AKoz6IcytkJpV/5fFAtZW1idMzGRkcECnrj877AWCyxCN54P088uY6UB27hk9n4UEW7YopGhN7gm2fC9RNYcp+ykFKA1LdCHjIIoLjpc8EoP/YGcCSJ7o/YU1PD2MR85uIlr+ChQSDMelAKeLB61uokfo/7IRDhWcffiYoCgY+ybXHPWlkb9Xp2VIWoQNlUVEUO84/njbeknpGIioxUEHgsMgWOjyNRgaoo+D1G9j0kTTE4TYJokUxwgCCoLwNRIbVNUOtwHcwN1km637PpyTFbvrBgzfqh/dV//Ynlen31dWHc5V8rRZdXF2A3INU3a42ElYQ6KLLUNH3g/RmiGj6XKwokoDldlXLVYOOQBFVUYh/sJNyu5wz25XDIOe/0+PsCnUU8RGCTdR83QtXi+NxlPtOTQ4mtq5RCBerw2cffOgu0PNkSyIN196eOJEUcI7/eoKJIWIMxB4qFEZu7eMluvPGmDQhYAe16bYFmzBkSNYJOkk5ZP3U6trW5rmbau+uPPIlE8RfWre4jiS8N/xFf4Xer8ZK/sgNKESz3BpL+dR4M80DqyV9nXhuIWXE/wXKLAVZSGfYNB6hTIifUxC2s+CQRFi2Ukp8Yg/1hxYWbhymxZskB5HMGoBrdVhLk1RQCnyWzZ976Z8e1GsGo5JyK4xGvR/d3GieeGZ/h3NV27Wvgq76SAP6Txlk78DkbpeEMTj6f0KTuaa+N5dvC5GOjNv2+am+GazgSbxGsr4yU7Ye/+wc2MXfZjk569ujebbt78z2rbj+EGX/qrT31OsJvxPeP5wznJEE/z6dLH5nwXOK+5c+A/bEwTISSc1NHMNZPYT5zHqvxMT2tOOOCPOwsYOsP0U8bjwmSX74unNBH4KAEGEVSOAdUaaEeN6f7cFqJu78PZwLvzznGC/Eo/+7b78i+afm5G6pcfPfnP7OP3/97e+HqBVucmVQPoP29um1V9+3R1rrNTUzZdGXEvaoZgnxGcxqQEDkZCdN+9UjnojeqjCX4ZH/cX+wr4aTMk+aO9iRx26d9WuI55/uWN1mNc/F0DAFoHIBIgrrD5xKqVlR5wl7L3tTvWSmXs4vLszY5WrA8CXTwFvYlmVICRzilakeav6LeQ6U88Obh+8cN6/RM/3f7wXYp48+A/Z5Ef2Z23v7w3/6R5UtlJYkk8I2To0BUkOAXLZdGRd0XOEUSSexw794d2dDsb29ZakAlTM7yah6LrSENn1ECOghJzLl7ULVjNTIPdnKaR7Gxtqv6NIZxLoV9FqIMsCG5kZzfY8/sdcHmVMC9VI3+eW4J6s9NwKbI2ydIIeObDXuAPHn/9ud4Wp0YY6/zCz0ZB8V5dToHTi2k4g5zXm0Z388txdzyKTYchajgPGTs4v5AfOIAp8cXnH1RsBH7W7DWBVgO1chuSxH3kEgIDeODdFpATZKoiDaNcc9Pvja538S9OhK80bOZ+yGOlO0ERAUNNOWbnbPFPBYzafv88ztSB/OYiEtfe/1VXXOpgN3Nvjd2lpgJm9NRVftgVSsQ/aShPQjVcqfVtFyqb//id75vuWzKPv7gQxsdGbf9as3W1jZt5cKK7e1vq5LitddeFphG3jE9N+9KccAXiaPywQIlbeXRUdtafeSVQ722qhiwtaCxKMBXda8q2yfWJeTV1tZjgRTkMpAMjBc2VoCE169fk8UjKvvlpRVbXFyS+pJ7aPF/68TGymW7evmSPXh43y5fumQbm5tWKJZt6/G+egBgKeH7GnFjT8KkxaVFOzjYVdX1/ft3BRjdeOGG3bhxQ30b/uQnP7F6/UigMWBKH68LbGgKJfm3Hxwda72SCgqYLSBsO1E+CejIHIOYYB9R5SKCCpSj7RMRO5Ky0aA3isRyGesgUIIQDj3p2CO8l6HHnFHwwJ4xPjZiXSoFAFezae+1KGsPn9+sbfUGAOYamEhUlLCoqtmjXKzlzX9Zq61G0ytJEJvlsrp3YkS8+Dk2uT9ICeWHqK+nZwX0QwpAZvB82aoRCCBCY4saGxlxW91Mysqj9DLMqRcgfUcgLFB0HxxWdZ1U15CHIvjj2lAPQzCRs2OBonsPYiqBtUXP2znHuE7FIwCTEj+Rd3nFNj+nGjEC3Pwb4J/+KxxHVNCzJqhOIudVFW6aCqS8NY9rNjk2Zr/3L/653btzS/kLFmnFUkbOAJAUIosl5uNsMdvZ3Faz93F6XdDrSFbH5P45NUBH0FYqj1ir3ZP9kwO7KSuUy7Z3cCBgrtk4tnt37tgPfuu7Sj2ODg5UVYHS/29+9kv1NBik89YGx85iMdbQHCXeoVGyKm1QX4ccSnFvsDmMfe4A25XLht4VXKPjDtjnBfJe1ffktJ6PUhEju6/gPqEqihT7CcRfT+cueb/6FwgbGHh/R1UHQQ44EO2hb8ySYswQBKOhabdcL1QFwzkiWZETzCIxsXYzK+aytjA7Zdley248d8WW52asurcrz/9HG1s2MTNr2/uHdtxEcJqzpaUVYRmq0mk2dZ3EX8rzseemD4oarGMTVhKoSkNhroVxYB5z8TwHTr5YtamemrJ2HKhnJvsTObcj521bGivaj7/3bTvcXrcSJN8ga+9/9tAaaVg6JynARqiSqtWPvYppfEzCKAgP1hDAtOy5tP4YGxdTaI8oOHkEeciXV8z4niQRJ3MZdw9Zf2W19lwwMbBiIS/glzkXCUD2Sp6VKqFK9O7MCUOBuNKepdzUcRLeWyLWk5b2buJvzgVezxr0cfHm356jeQzJ9YkYKRRE9PgT9qiDfBrsDSKLL+6La2Q9+f7klWNcu2y3Mi5y7SNM1bPxPq/k4+y0BaqLUgP7wQ9+YHfv3lP+C/nJ3FfOEFxOKlit0dtHYoZQqSohQN0rErG0ApjH0o51BuZBD9e0WTGfscWFGRsbH9GzkwABC9bdfV1fo921hcVlW7pwSfMRlACLLPZlzmasWTnjaTDtvZOobKtof/VqJ/Z2x+ZO2D+bJ7oPphgEsFdCeQ6qeawqylh1B4FN02q3R9ceFyqKifkl8hMJ5ngVmB9OJMSt7WbTLizO2dzMtGKK7Z09/M90D/T3EBlRzKvyix5bwwbzlrLJSe9jdHh44JWZwb2G3pj0B+J7Ek3n8iJiaEwOIc5ezNwHU2NNsL4gflkXXDdY5DdExVPT5m9+8Js6AldyBGwx2Qje0p4lKCCLG67OldDkUvYYAYjX4lfQ54xlTDCSwFfcVEks3CvQAZgI6EQwln+79ZF7EPJ/VBrKsqDbkf8qC1bJE8okFCI5yAonBBQMQEioCsE9nRUIKEDLOvsoVYV7ApIwDK+deyRI5fNj4spmXixZo+0+iJRbSQ0Q1NtsMGoyyAGCJ1+7LcafA4RrlLVQUODr0MHegCoGlO+hUbk2SJq4QmQEGxau368tNEUSV+MBSXfA4Y1HsDcao8kfVkzYAJ02BvVKFTUrTblfJ8ED/1NeBmkjiFoNkx0mIYDjsAXgwQsWkokxVOAWqmlyWYAuxppDoC3Qg0oRVAsEZM02jbYy6keAcgplGqWQfB6ba6/fsemVi96cPYxPnH9SAGiO+VcEN/37TlSQXPAMGTMOJ8YwEhUq8wxEBRt4vXqoYJnAvVhBEeUN1LB+0nOBPMpD+phNTnuPCsrimQNSyz6BqFAlQ1BonicqIhCSBET8Os8TFT4H0/2uzU5P2uLKgqUHHfvL//rfrHfkDQVlNdZuD20OFAyPjOh5Dkva1Vy+aJXQDwbQnbXBtROIpVOuzLhPVUCtYb0E4XAW+AIoc9VpXJfxGTzte0lCIfk7p2DkKVERm9VrXAOcB7B5vqIizgP/7KgAD57h4YIc2Dv13xfAQiCSqKaIP+dXFLxKOVW0SmXcli4/Y5dv3LAupCL2Fb2ONfDuHZDAtFS2zLqdnZ3VJ25tbtij25/Z3uaa9bA+o/FhUGN8HVERQbIngYya3wkF9XkQ7fwcGi6KJ/xFYx5sP+L4x3mXJAZIgr3ZfFhfJPmhKkEVQOcAuFNlu1dpCHAPYXM6NOrFVzaVK4io8HJemqQHoiKkXHGfT4Jv54GquN69wucMvnhmTsaxTN7z145N4gXnxzmOz5OA/+T3hMMnGq596TMTAHq8F//Twd04b2Mw7GcbVhyj9sf/2/9h3/vR79vdB2v2F3/6E/vovb+2o721M9UE5z/v1yEq+J1TosKt0OgbQfNjF1P7WhqSrKpQyA1B8+QewJTvQVREgT9kcGiALXWbSNnzhFsgKhLE7en8DDUUqPWlwHaLIX2Xs5fEk8rM0NdEgDFjFog5xQeq2AokHL20KhX77R/8UMqrN7/zA/vle+/an/+P/2btZs0uLc7ZhYVZgeJ7+0dWbTTszoP7tjgzaxOFkuwTB7m0LV5c0Zn38Sefyr6ExB2iQo2+Q98Cr1QMVj2heiommcO1dZ6USZ+SFDG2ifsm+/T59R7/7dUopxUu/v0AgocxcQ/trqVQtQ76Njc5aYtzE1YupKycy1uBpBhwiscOWOUjFxI9fpf8Kq/qUCnfWl2rHzdt/+DYasctr8ChhxaKYJ3hA3v+2gv24x//rpR37XbPdnZ37biJr3/B8rmilUj8BRr0rH7UFFHB/FtdfWB3b31m1d1tQ9ZACT3+0yjxotI+xn3s7QdHR3bYarteNI55rCiRJjB4J0d7PVUZhEqTcz1vzj+js2vKrU+0xokhEuRQ3Lckignk2dP2HPb0J52ZZ9fSP5SoCCfil+aBx+nxHH3SNcX90qsP8lrrV65csQpqPTUNj/29nJzgXhn3aKXI73uvEre6idXTqqgIsVpyD4l/j3vLeaIiVknI4zqQnk8SQsS1ESswAHv9vQHBsM2kN5gLOvw9s7ZUWAH2tNu37wpMA6QcHSnbd773HasfHiryqNXq9uDRqirHBaCrmbFXXbsdTF/x7DGKaRrKp/r2z3/0XRstF+2jDz+0eh3gMWNbj3flaX54uGMT4yV7441XFX/TiDSTz6pxcmkCi1GvhKAJbOgKZof7VVnOHe7v2dTMlN2/fUfAFUQDwPPPfvYL9SIgZ6F5Mv0NeMgS0jQaagyOXeWFiyu2u7Mr0uQH3/+hXX/pZcUyWOGub6zaL9/90MZLOfv+974rQQbAt9Z5Omerq1v24IFXVCj/yphNjI8KSMMS5sKFJXvppWt2++4XdufzB2b9js3NLdhLL71kM7Mzdv/eHbt7544d7O3bWGVMBMzG5mNL5Up2eNSQgp69gfkSFcyAYyIiFa9gpxu82uWV39K54wCxk48SSuhJe+U9ZLJbnjq4HKtMUFSrCqRcUW4J8JSKTe8FXsZqtYEDq1Sls2cG0B57DtmZqs9f6H2BvZlU226jI6977OoqZQGDVJ8g5CL+4WzieUIM0VA7xrjsN+SiWHZQgXLcOpHVHWrzHOcp1SD9no1O0gQ4Y13A3FTKLizNCkx848037d69e9qfJTDDVocKM3JHS6vHBMQOwCkAseefJyJcALjYR1krUVGsfgJhbLkuKfZlD+Ngqary6dmniu8Tz1tDni6hFeBn81g9VmgX++L15+y3f/RbtvbFTYGR0/PT1j9pWKfbst3dHbchnplRL8dOq2Unda/AJGefm51XrgLAS58uXU+eswBxVdsera3rvF24cNG29w9sfGpKoD/g682PP7U333jNxkdHbWF21vZ2t3WW/d0vPlCD+E6f/gosupx+hzwW0s1d5MArCuoxoHsHlGQvk9qZn+UkmiQHkxWePOtd+c6DdeAdoPjUZox9E/Awistk9RyaYrM38ex55vWAG/AsASG9Ks3zfq+cclHHMIYI8Xiseue9yIHZK4Ql4HYhEYQ3ClaoQG+ITk+9FQBRxwpZ654c2VgpZ2OlonpOlGgW3+3b3//yQ2t1qDKhNwLCrb6VsceGpO11bf+Avjg+Ll5lVgj9SL0KSb1L0gDqvo5ZK55v5dRMm2b13CfPXH1BESw2G17ZpD6ZLbsyN2lvv/y8pdt1m5+eto39Y/urdz+1huVVGTMYuJrfK2/dSQDwGQU6JAVgMs/eRWv8rK9zDGJReSc2laDlYVGyhlgDbvPjRGq5TFNo7PpaIufUaB0LuTz9aArezySMg5P4XvHEGcK6EKnT7Vq54tbcEd9yiyePb6O9uioa8rh6+Fgl8zPii/jlFc5uTcZeyJxRo216gagfjdtwc2OyK1de5/sb6wtgnubVVBYS08UeZDF/Uw4LlmEp9eLw/dbdN1D4s88R+0axpPZkSFmcCahC4vqoRBRxfixbRvZkBCcnxw0bKeSMqy2BQVGR0e7b9MyoqtPYZycnIS7GtPapQNx8vGuPtnZsgLVjnz4PYF1e/Ys4gvsk7gQzcqGCP1LFL4ylzoqU9UJTe2FrWEAhgAqVKJw70YJQcQUW28GNQGd0wBV4rvwddw3GUqIN9dHhObSUnxRyacunzEax7n7msmzB1rZ2zGgIrrEMFT6loi0tLqpnFCLYUonzN6NYam52TuQFpArPDXHC0tKC5sTm9pbiEwhqKrynp2YlSIAAZ7xZf6w7WfkVPAZn/pP7fENUfBUi8M3PfiNHYMXcliOqrQBB3auPzd83dSlXQvmhVGXBfkmltulMKLt1AMzBZW9KE0vw2eRo1saGH8vJd/d2deCqBL3bFvCtAyyw1VJ2Uf4YAn02dTWhnpmxR6uP9H1t4ByWUkqYNiESlP29PYHxbGgcZmy+NBXjoNS+pIQ95aAdm4qaJDvoQXAFS446YnZ6xirlspKDTMH7bbAx8BoayhFkUapF02qV8IoUGcg2BtWTiAVUzAlCIgySxoGNFvKGX1QvhIx7TLp9i0JEb5QVku/oUhnZde/lUVQ589L8nIAjkiWUS/VjmG7vMSGFBWXNKj0lyPAG6FRZOOHh5bHyUUVtSRlcq22w6GyoUn1onHpetkkDwHDyczgQOHAYEnygGuCA5LoJdlHJ0J8Ckokr4ZqnVy4MKwySQFpMkpPgoTPcIXkO7xsrKuJBr2ScUscEUaFS6oOa5gjEUZKoKFdGfe7R3yFPU+2BTUxNal4z9z2Y/zJR4d6CCSuJhM94TPjjgZcEJr5EVASiKtPv2fzclM0uzFohY/bXP/mJtfH5DNZWvhadFCMQU5M2AgEBBl6OSiCInZSawXZO1I8FlRwKQcJY7n99Y9PW96pq8hSBiyE44Md9sHU6rWA4Dx7EhGUIriVsXJI/SxIVeDnyHCJRwTr7dYiKM2DmOWFqBE68ibsHnCqTDWBK8vrifsTPIKtGx6bs4rPXbPbSJWspsHGyDRAjn8kJnOD9VFExMy3ibm39kSoqqjtbaqadgqgI3rG/NlGRqDhxSXYAdGPlgKeD0YErolJPPU+eCLY/hahIgmbsRZAVyS9PQmKfkrNK4SRRoShWDSodBERARbC+MD9r1cNjO6gdCgT1igrvP+IImr9nEpx90hqJZMZwLn1NRcX/l0TF+WsbJooJsFkA+q9JVCT3L41v+pSo8PPRz0r1dioU7M23v28//r0/sl9+8Ind/PgDW39w0xq1bbfFeEphzdcTFU6SiIgGbFRDRsgA/OXltfREosIEmgcLs1jFp/3VrJdJCBHCWEgZKW9gX9vJvSC5B355DvgD1hCrcjHYxfDZoYpSFpLqX+E2jRrLBGFEw1Ql58ESkvH8re9+zy5evGSZXMn++5/8N9taW7XpsbItTE/Y/MykzomdWsOmFhftVx99YOPFkk3m8QfPW7qQtfmVRVWuffrZLTX7AxSimTZKXZ6HFPz/CKKCtZOcZ6d7HPf9ZaIinieRqHjiuMo9gKpJkpSOFNEjhbxdWlqyUj5lI8WMfIOJCaisYE1KVCJVOp6+Hg8B3FBdGMUgEFmdzsB2q0f2aGPbagB7WF9QTdHHmiBn/+yd79q3vvVtqTHb3b7OnXqjZoUiQI/bPomo6Pbs6OjY6scNq4yMWiY9sEf37tq7P/+p9bstK+Vo+J1RjyD5xcf9KJDMjVbLduvHUlb6vHSCSNIKepyEZvNJAnM4tud20PP7ZvLHrMkhOcQ5FYjH4feCaGYYlj1ld3ZbtaeTFf6zfxpREcfI923JqYdnyhlyNRCRfE8AJNYUlrKVlRWbmnJhRpxnMcaKscqTiAopGAXweKx1nqiIYoEYO/BnkqjQnhcs8FQ9FZ518vXn44wY+6yvb+h8FFFBLBkaebrKGRAyZyvli9Zu9WxtdVOAMWA+IM7v/8G/kRXK7uNtu33nrnqpMJ9A5yWegOiQVZWvJ841VSrnsjYxVrZvvfGy5XNp+/TjTyyVyuu8o/8EVbjNZs1GRwr2xhuvCHwGcC+FhpgowrOofisVgfIAylmU+qxFxUID295Yt9VHq7KgW758RcD/n/3pX9ni0pKuk2c7OzOndQtQQTNRVMJUK6+sLNnm5qY16k379lvv2PMvvmTt42P1HQAsPqru2a2Pb9rLL96wxkk9EN+smZStr23b4WFdf0edCgBTLLnoitxhZWURcaiNT0/aeKViX3z2ud2790AiritXLtvc/IzskJh+6w/X7fHOjir19mt1y2SLtlc9tAKWMaGhsKrGsRlSJbCvD8gbPOaJackfAOu9+amreR08UyI5tMLhLMD61NXTiIwQgrnoRP10NBcAp0yq4njOqmIfeD9U70fhE0IfCTCwQwngIApo5iZWu8wt4kIqXrDZGKcHyMAU7zBmDnCTP3qeMj01pRwJSy/W0N4uVjFt9bAolr2RNxY2VLlNYvNRwr1goCqW0ckx66PihUTmGji3czk7PDi0ialpKZA/+PhjWd1QtXFYr9ve7p7mFTk2Y4HQJqqz47qKa8StO71HA4C3+iSpL1DoYcP3RSz5/4wVuUWMzTgzEMnh1NxtH9uVlQX74ffftnS/bc2jqo2NlBVPYxlEbL67vSMcYW5x0UZKFatVD1VlQG8YroPPYEwhaxgb5gp5KtUUNJ2tq4oROtutrSSePDrSOlycn7eJsTGbGh+3bA4yNW9/+dfvitxotHqWzhaDEA3VMdVhANrYJjPjOQsRL3n/zaigZjDYFxh7gG45H5DPyv/d82Oul/wZ8DC6Q0BEMI5yMQjnRrw/Jz+wG8Iq2Xs/kOsDgpPHxT2TOCPG4cOjJVTvSSQqrMXPPvYn8nPOfb6jKg+91nv/Ua2E7c7K4pw1qnv2/NVlq+3tWBtBFv1B+31bvnLFbt66Z51eSv73qOQZ98ZJ0+onTYGgzCmuSzhC4P5VBZTyyiKvrvWzhUoJ1p7mYrAGI65hLIUDEfcGsRNYAwQCTaufXZqxN65ftvbhno2PVNSb4hcf3bH91kC9RtJpAOe0BCuAwAJ0IfqC7R+fxY+8IbtX0pPDR4wAZYsQkCC0hSBgPXBd4EKQURAZ4ErgUOTV2MLRL4b5wVp2waBXY6lh/QnVGQMbH6enh1u90c9DPUWxxgwoehResA5rh7XQJzSt/jxYfzEn4muiWFfi2YxXRpD7J/N1OY6wLoNI2CvKgkA3iHJ5Vqw5hGSy9qb3A/aXCFoRdsY4B0Kefbg/sAvLixpDGtgzr8n1uEbOKVlkBwBf1UFBGMo4KXZEKBAs4Kk0YM9I9/s2Bjl3VLNOo2U5qsYKeZudnVDvGc7aZrNvuQJtFgs2PTtrjcaxPdras0w+Y016bGaxRXfyhTnPOhR+oB5VnoNHLDKuF5Ep4IWqynWxaexnGvvuktuDDUrsajiKtIaE0WlFyukcZp2yD0RnD2GI4FHths5ayMDnn33Gbt78zHYPjuRakQnzi/2Vaq7Z2Rnb3Nh0silHfEw1Tkn3wJhiDUbfG+1/pYKEUo93dm1ifExjTH/dsdEJq9UOJWwDy8QSkGoNERX0B267kw3X+w1R8VTo5Jsf/KaOwCUaO/Vo6NwR66+eCfJQpBEzfzpQzYYpcB01iwI+L99z3216EdBcCiuavJd8KnDzQ8JZ67I33yG5VANslN+hVI0KCzzugjdf9LdNcfdGtgAAIABJREFUMs7++V0tVGcUffOQMlvlw/6+fD6edjRzgjxQv4lQxk5ALJAoqNwVuKrawZUWChQoNeUwVGPYrGwRYCzVCJrmQ6EqROV7Ujh47w5tZlITSIunQ4/AV4RKUK1xyHDNCiCDUiWqVtrBqonXcpAzvg5seFmbEyyAXq48pcJBvS9SKRsplW1uZkaVFQQPAKw8U1RzKC9cI+SBIYE5yQFfkDCHtZoIC/VMCEGQAjeqTtSQDg/LUY0pn8XB5ZYb3vibcUd5hOKIoECNm0RSuN9pOkszIFQ2+JXS06Fn08sr7uUb1HD+/JwYkE9mAAhFVgUbEFVVAMaEypO43qKyRWoXCDKVTRJIt61xSNCeEvBceEJFhbyE8RpM9QJR0VdZoatTQkM/gYUOqvFZw+cX7V2itU+iGiEJVHCd8R5iVQSJMfMn0+/a/Oy0zS3NWr/dtL/5yX+3DF698v7EYqypRookhNwDY5+DKGo09D+BCkQFaysSFTSDJonhOaOcY66RRD7Y3FbTQve5PLUfcusc7jVamCQbkp6ipOfBFyWaodlXBBeSYLMHa6G5XFDBPKmiIiZT50HNp/07Bk1qxNv3fYvvJe3A4rVFcJTAFJXE2OSMiIrK9IydELBhfXbSsuPaoeVS2DaEdVGpKCFlfu/ubtv22gPb21q3+sGhpSCqEhUV8v8cbv6+9mNjcQFqYV85D8THvjlnz40w3sGi5XQMfr3TJQmqJT8vPp8kUXH+58Lhz33MWaLCKwO0T4aEHzXhpYsr9uDRhjfJU8CaEfDDvbvIK/wXgO14jeefe/KjnwQoxu8N7zGoz74KfIzvmVSqJV//JOA4eR1nQL/AGTyRIFAW92UyZvhaCJ4AziTPNM4Pzpqli1ftmedfsbv3V+346MAO9lat3agpKfiyycwpg3MKdodeEJGFD5UcSSBQ6waEgSorNSo5JU/0swAMDezJRIW84dOupNP7xqIXkln1n3ECLN7nWcA02HMlep6cNix2SwwlOEEpr9kjpbh7YsfzmfPVrZ/8LORnwz5WofLwyqVLig329g+sWa9bIZWy5dkpm5um0W5WVX77J31750c/si/ufmG33v/Q5vC+RSE3VrbJ2Rnts2vrG/bo0brO/yOUoDQtJaYRqPXlioqhZC8xgc7MlUBUDOdkYl9IVrPx8yRJnJwB5+e6dovQxyMSFdNjo7Y8N2epXkvWT+OVEStmIQ28chLglIcH2KsqUCya8tgAOSioMdZpl7WDestWt/bs0cam1QF5ABjSgDZZ+9e//wd2kUa6uYIUmdXqviy38kUS3LzmdZbqnV7fjmp12ZYAHpeKOVt/+MD+7m//2vq9lhVppJrPWpHXh0rF5Pnf6ffV/BzrhEhQJAkLzY/YZyFh43b+DP66fcLFCcFChXMyVFNqiIP1k1sdBnIgPMjk+/J3N+k8rSw6v2/F6/JnHhtof5mNTM6d8+TDGYA/2F5Glvv0tac9aASWqbGun/sLCwvDisHkvuTkRLRScCKCn8ez9TxRcVpp4rGDKhuC4CWewQh+ovVTnNtJUUH8nqpUfeCGwCj/jFYqKBL9Wlyljsr2tKLCKysuVC5aG/u8h2sCOqemJ61xfGQ3XrxmC3OzNjO/aAe7uwIpyRMQIOGTPTk5MVQm8nnYJskqtd+3jfWHdnFlQaKdv6chdaFszdbAdvaqaiDb62IflbPXXn1Rft9w84AgaUghbEkAqttUbfRt8eIF9WfhRbJEOzy09UeritOnpmZsdGra7t76wj759KaNjo3byMiY4hbAN4gOGmcyveYXZlU1gS0TynksPcZGJ1UtB2BIvzsA2bHRsq3de2hvfftbduvzmwJfl1ZWrNXqiqi4d/+R+h1ATFy8tKI4E2so/qT3AL1jvrj9uWyKXv/WW6rM+uW7v7IH91ftuecu2n51z5aXFu3G9RetVq9buzuwjz753KqyDkGvwPr32F79rOi9l06JlHD7j4zIF5qKYhupyovQMBvARf0EAWKVc4S8oG8usJIAzPPQKNwC3GJOHh4c6HP4O/lrbIgtoD70M1OPCoQC9Ftst4c9zvhMiHeeD9c1MzMrMQEAHoA1a2J6esYOjw7t3r379vzzz2vMmZsSseVyuj4RKrm87exs63e2trdkb4Tiu5B2Qdxv/+C79srb/8xaR4c6V1h7tf2q1apVt5rp91RdoByH5u/NlixReH6ofZkT2ILQc0W9FGjkXSyKLIk2ruQyAK6Mt2x9Q6zM2vJm2V7dXT8+dmsj2bk0lBeTr0qUEix61zbwiS+rKXu9VrWFmbJ97+3XrJSDNu5YgYawU9PqZI2yfGebhvAH6v8HHpBNe75C02UayGKdo6bGKbO96p4A8dHRcd0zVoRY/aD+397bF6moyLOHmOxYcQDX0mzWRTAur6zYX/zlzyTCOGogKiBXzQtoLxTAL7AvcsDcPfC9cj42h2c8BMoGe2P+zbwYAsmolUslj2uD0ITnRX4mYDmQEewrynuxjMZGLBC6TWzmKhUXDgbBGPsPhABfzH1IyaH1biAp4nMUcRTAWXAZ9dHSWe2VuZ6fajdVJSr/eO2lFyzVadqlpRm7sDBv97/43Hb2dm33sGbZUsWqtaa1+4gT+7Lj0h4c3BEO6jVZwzmZDfbCPKJaEmshjwOZO+zHXAe2d8wZAHvICno3cJ6rkXHfZEcNFgFB5s4IA8sMenZ5fsJef/6SFQZtm52ctEePD+z9z9csNTolC6+TE3qT0qA4pb4/wqdU7dK2vf195R08s+iUIeurIGpwwpPp6E2Wo5MFYyrrZa0Fr5Kcn5/T9R0dHurfPCvfd939gjWC0JZ7lJVcsE6TDVe/L2GrYtaAKfmYxB6efa86gKD2MsbQ+9Rt4/g8tzJ3rID3EZkS+i5KrBmsJ3ke/gycEOG1jnthIcbv5YI992CIk8l3lPgdkUGI25lnGeIC9c2s2DPPPOO2n9WqsAX2A/Ahr+Q67ZlJ1Qj3HvEiP9t57k7clQoujrmwuGALM1NkE3ZU3Vc/skG6b2sbB1bMmXrKsv7oh0H/UEjtu49W7aSX0rNGOCPxLrG2enT0NU9x9NC5QmNs2Qu64FfiWwSLskXzimzOBvX6UcN7F26xr6ovTejrpCblQ0uwnmzueS8sIbWmZD/oX35mpe24fqQ9cLJcEglDQ3LOZkh6qEN6UzA+stEvFGyRtffgvvdV8ejQ8YjxMY01ggTmMLgrjcMRGqxtbNnkxKjHDv2BTYxPaS8lhsbpRvbWuG60WnLaOGm29Ry0X2UX3vpy3phITL756zcj8Js2AuONhjY2LeBicRjcceByKLARsqgIxgh6WPzaNAmkAqjsDaqj93mwaglNuNnkXPnsfS3YQAiAosdcVFYlvYYpj3UC5NSPOv47bhjOpLsNEGXNqMU47AE7uBaUPyhZuH6VA4deCALFUeSgjKShV/BE9gM5qOhDdQXgcDxAxGajpg7NAFV+xngEX0AOaL7Y9BWwSoXgyZ43uHKGOpbh+qHkG5eXwQPY+LWfolPB/ooAJqFgl5pN4+1BBEQFza5JewkcmvWGmhSx+R03GyIaIG0InFBuoTggYOeaCHhJuFCqkEhwP7DbHKAcevjlUUosH0p6XLRaOkDwymMz5qBQIEzD8+Mjy6PKOoHw6ojxbTTqSjKkoFDD7Z7NXLigcYl+xfGZumLh6UQFKjqClliFEQ92ATvBU1QWIWK8O9as1TWHOFzzpeLQ+mlkZNwbqZXKIip6g46sn5hPEBXuEeml9jEY8MD+y0RF0ufZjyCv7kgCwbFslOvGVovyRjXNGvRsbmbKZhdnrH64Z+/+xV9ZoY/C1a2fCG74n7Uir1kOp9DIDZUX5easU7yXORCpqEBhNzMzp4Qgk3Grh+rBod1d27RmaBLO93St8vb+MlERf57cy5LAT/z7eaIirmUHS9yaJVboQBydJyoIniKgcf6zkv+OzyCCIXFs4/OIdhICikKgx/fi/iEVRRmiYtaWrz5r+dFxawu8oWn8iTVqhwLzCESZfyRAU1OTepq12oG1jw9s7cEdW73/UB7wUnxHoyQ3ifWvQPYMiYoAbkdSMt6TwKuE6vb8meGVGk8HxL7qjImBa3yGZwCvhPVTcn7G90s28I5jN/z94E8v+x3t7Smbmpyw6akJ23q8p7eIyr5o7UDiJSAxUVFxBmQb2tg8Oaw6DwJ+6b5DFclXjccpmH+2QXTymob3n6igiD8fPrNARjzxtYmfRSLC1T7h3glfo8VgQsWMLzXnxOLSJWv3UlLqDrBvO9qzbsfPk9PPCzZST7lZjRVb3/DMTNBnAaDUvomKWJUuvv6VnEY7NZI8zWEHNJNjJ6ICbWPohaKqPx8kV/fJ6/o8UXFKqsRnmZxXPmzeYSEU3qhXRST3WANRwc65rn1ZCjLX0fdTbksg8kzNLPya5ufmVc5/VK1aut2xZy9dtInxEWt1mtbotq0+yNv3/+W/klLv//z3/97GUhkbyWdtdHLUJmamh/Yad+7ct25/YI1mW4AERAXCiLNEBbSKykJExD91Lkku4F/J/Uzz4lwj5SSJl1yTcXyTc5IYA5WXqlj7XZsZH7G5qWnLWc+mx0o2QXUdFgayfHE1H7FD7DUAUeFJXmi5gSoRAtoy1hnkrNlL20effWa37t6Vz3Eql7aR0RH7g3/7RzYxMWV5mld2+3ZwUPXzv4h1CM08MyIquNej2rEdHB7pHMYa4OG9O/bez39qg35HFRXygg7KPcWLofKO++Q57x0fK5kjaXRzjCDkYCwTYx5Gdzh/tVF95deXST+9nLk9VMaexqDD/ejc+ybJiEhUDJ9RQsAwPHeHVYxPJyrOX/Z54mK4dmNcGG6V150nEHivSFTwd2wNsS3iK861GHvFSgr+HSsmouoXoBOSYBizJ6xeI5gR3y/+SdVxBHA9xj4VFcT5HAmU86QOr49EhXz+AWSwVTpHVMQeHPkjqpMz1mqhiOxZqQjYnbI3v/W6FdjnBqaGlI+3d0Scvf3Od4bV4ajnPYcZqDpoenLSdrcf2872hr3x+ks2OzdjH773K5ucnrONzart7h8IIOh2UdmX7ZWXr1uqT2PnluVKRWt22gKGl69cFRiBWAQP74XFJcums4rFPnnvV5ZJeaUL83p+fsE2Nx9r/qO4BcgFvKBHwebmlttdpFJ29eplq1Z31QsOG6/dnapAnI3NLbuwcsHm5mZUxdxqNmR/SqPsiUnPAQ5rR7I+fXB/zTo9ngf2tBk7rFW1f7F2IR0XFmft+vVn7cMPfxUaTDft1Vdfs+eeuy7bp08/+dgbj5opF8A/dWnloqVzJdl4AKECElOtRQ6FPamqkQOxxk4pSxyqs1Mp29nZFbDD66le43ekuJe9DGCq90wB7CkGSykp3Ftudzo6Pmb1I6o5qJBOizyXsAcxlB9UetYAXQA66ndwfCzQByQVe99iMW/HR8cCj6emp6T+R6T28isvSRFL/srrBRYWCvbhRx+LaAEMI54D3FpeWvJm1cH6d29n12bn5mxiYgT5lq0+fKhqikG3bxcvXbALFy5YsYL1zLjI4/WHq9ao1xXTQ9KCk2EdxVxgr15dXbPH27s2Nj4hYSHVbePM1Z095WJSIlP5LRLCrY9iNSLzMQKZjBv2vAicnDgE5AKox/L5WM+KM/flV16xL774QvcFaLm/TwNxGmQ37PLKlP3wO29aOtO1zQd3VHlC7jE1PW9WHLGt+4/UQ+Wf/fYPrLFblT3KSZMG3OOaryiBZeUla62TQLYwlBnVPbBGM4Wira1v2ezCos4QCI+RSknVGhBo5LuH9ap6LPzpX/7cAfMMwkICHIiwmvdV6lJlkBcJ55WR3piYMWPecKarj0+0dFZ/AAhG9hJXv3tfA+IQyA8qQLz/AmOM1RHAI+/lxK6TtyjuEZdRWSYlOBUaCD5lj+re975XOgaQCBKG1UdSkwerKa+IyShvl3WN+sXFHnB+PkJgYVW3ND9r/UbNjg/3baSYs0tLi1aqVMzyOds9PLJPPrttbRpWC+AuqNeUd7sayAKK/R/LRgfFOStYD+ACgOhNzRVIIMbH8RfWqPdQYF1Q5QIhB/EFwcSzklW1xJ00lWzbS1dW7JmlKavvbtrKwryt7R7ZLz6+b8WpORudmrWTRt2OjmtqHJ/NF612dKS9BMEqn08PGPYIEcxac/RY8y/ZdBUc8Fa/Gsi3YH0bbeMUTaTNZudmrV6veS/FbkekFEQjebVEkqFvE5URWmeptNFPAIskCCfI3kg6xPGCsPRnN9B1+vepfMK23EmMiGVEAaSHs4gmiL9dGBzPYd0TtkPhmoKFh8LPeIbyp5/RCERPQi+qgdauSEeAfFwDIHupfhKCz5pzAm1ubm4oQOTcjvGq5oEcTtxOfXRshChMOAVjCxdyhOiVqhIwohbVvRlbmp20Zy5fFOlBpM9a0R62wzOlmXfP8qWKlUcrtrqxZW0CXvJyKlgCHqZesaGnqz+LaDOb6E8Ycp94vSI4Uk5Ey24LV4qc411+XwNVzbCnUgGmvJb5zevDmIucOnby2a3TO5pPxBXYlqW6LVuYnbblxSX79OZN292vWQp7QhFWrmnhLBkfG5MVXoxvIMBaJ20bGxuV7ZOEC30sxbo6B8hLtnf3bGJi3HsADqgOLCsG5ufEKtjd835UVkJeNBsIyyGks98QFV8T9X/z49/AEZg4YSG4O7kA1cBKEtsJYA/VFM7oUyJNEOb+iL6ZElKcJoRJckGJmSyn3U9UoESwiOC9SK691M29+aJF0iAwqXy+QFEtei8JdqLBKxm86XewTcKH0HvC6QDj5wLtQvDGtbDRqsls8FxU5YbK2L15USzxUrVIaMbkG58DThyyUj5IUezkAffgtkrOPA99BRUdh3rJmBAGkMLH0TenOF6qPgkApjz1QpNYL9eN9ixK7bwcWsFyTkkEGyEZPYEnAa43+yaQ8vGlvFili8mmkGpY6T6IBNqxlC82qENxBHHFmPFZjD1JzFkAvhvcXbyKotnChxr2nqbnMOzeIM0Jiq6TFf2uTS0vBxWGW3/FhJlrcbWFf8VkOQLSHNxYaAzni4iDUMXyVURFuWy5ctEDg2zOLSgyWTV590CmZVMz00PrJzWE/zWIimEDr2Fj9FM7lQgY85nMRb447CAqiIwIqrL9ns2i9l2etY1H9+2zd39peRRjWDzpUG0o2OBZSu2UpblVTuXdXjU0JqKCZyZf2c6JGvctLCwpyOJ5MV9QStx+tG4NqjUCKKmZlCAqok1UkpBIbmf/GKKC5x6JCoKjfypREcGPOLZO+sU+NqfNaOO9xXWDP2oRomJ6zhYuXrH8yJjxREjSqKhoHNXU9E+ql2xWKi+CQSXKaqjZFVFx65ObJjO1UJKqxOKriArZp4e1e05lG8mKJx0Z8X2TIGUStP+qY+ariIo+3sbBo/iJn5vA9b6OqEA9t7i4YI3jusAhfKtJAgAuqa4CDOLPjoLt0z4jp0QFgdZXH5j/MxMVEQyMd+DFJg7uxTWms06H11mLFfYv1jTBfmV0BANzOzxsKLkGbK4d7lqXCsV4soYG95EAfNKo+VkMqBqq7xJp75CIAKzj3MXZOIx9JCr8NQDLZ4mKuO6VDKdQL/k5KTsmzhd6JgEgaW9+ckVFXI9xT49/ClTl/wRRofPbf0HvJ89/kskwhwCQpTAjoY5VCiIo/DX0sPjDP/xDNfT86V/8pZVSGVuYnrJyuWDN7okdnjQsP71sb37vt2x6esL+03/4D9arHliJxvDjZXnjIrwAJHn8eNftSRptJd4QcV8mKmKydNa6LQks637/AURF3JeHtk+JdXJmH5AdFg1pnazA1m12asxmJ8atmDGbGRuxicqIjXHOZb0qNqWS+p612dcKeDCXYB2HCj/+jk0OTUwHmaJt7R/ZLz/61DZ2d6zLs8mbXbt2zd5+57s2MjpmuXzJOt2+1F6RqEAkIgtNERUksHWBTJxruVzabn920z761XuWGnSslCfxywtIjvt7TMy1b6RSdtRqC2BV813t+U5WqCIhkavGdTEE338tosKfzpCUCxZvQggTBGuISPyPxPsmSSd+BD52/isJwHs8Gytyfn2iIvme8TO1ds8RFZEojWs+3hfnWqxYJtm9fPmy38rQQsFVnVGpGcEZ2S5QMQz4KqLCxT8x9onvEd/ndL9woI4z9WlERZK0jkBL8uyORAV7JQIMYm2JC9onw8raKHYBHBtpVWzQS6nqgXldOzywvnXs1VdespESzd0z9t5776m/BDH4Cy++aEc1B56jHY4ajXY6qrI4Ojywk+aRff+3vqN59vnHn8onfa/asIPasQg7+q9hafH6qzfMeiei1gojZQlKmij1aaJKDkV1+nHT+8KxjjI521zbsP29AwccLa1+FICdxLQAWXha832A3Pv37st/GnD6lVdftkeP7mvtY+HF9/f2Dmxz47FduXLVHm9vqWL9yqULtrW6Zq+99qrVjg4U6zJOVNXdufNQPXioKt7b27el5XkpRfHJ7rZbtrgwa9l8yq5ff94erK3Zwy/uqL9HpTxqb739bYEi7WbDHjxct/ZJQ/dYqzctnS+JCK8fn1iNChAJx7y3HsQ8pABxgcjedMqO8LKnyiv0QFHOoZ5uCJbEGQYrI7dKFAFVoEcAcZjnlgh7JiYnpLAGBEoSvW4n5+S2e7m7Glwq3ABO8w+qUkhdVEkT8trl5WVdOyrbSrnihISZrDfIGbk2/Nx5PffE2PHeqqKXOM1JbERgo+Oj9v3vf8umpybtwe27dlCtusKZ3oKVsl2+dNlWLl2wR3fu2Um9YQcHhzqLoLc5I3nGnD8QWYC1xOsidnIFVUg9fLRq1cOaKrUZMKxfWTfkEIB1jAOkIQQN88v3A87xUwJd9rKFgu1SdUQsgZJ3YkI5CGMKIEze1Do5tl7r2BZmC/a9t1+1Uq5nzaNDr8RL5ayQo1l71R4+3JQr3WtvvK73gnDpdT0WUkPrDg29i7KcYS5gq3RYq9vM3JRtbu7awtKiPVjdsJn5BQF21SqqdVOPFgRGPI+93R174aVrNjs/b3/6Z3+rPLQ/YNy9wmToBqFeHVjXIXZLCaB0gj70zVPs5LssexYAI89RvQ/C/OFnkD2yGZYin72R5tJelaOxgXAJwkNwElWthFyc/ZAx9Ca42Nu4nY3yQwlDwi4fqincYjtYYgeAnX8P7ZflAOEN3PmCgOHe2Dty6ZTNTo6ZdU7swvyk9U5OrFk/VmXi6MyMTS/M2sc3v1AfD0BQ8l3Elop9jlGG03zd3Si4buafMIReX6IvCC+AX0U2EDk97+2gZtpUuyu2oyrFhYdcofZ4yBn1p8zKXu+Fi3P2zv/L3ns1SZadSWIeWkdkRmpVWrXW3QAG2BHLHcHdpfFh37gvNPJ38YFL4wtpRhptZzgDDGYwA9Gq0F3VpXXKSp0ZWgua+3dOxM3sqgKwBM2Isc4xTFVXZkbcuPeI77j75/7uNVT3tjA3PY0nm/u4fncd8ckZxNJZVCvHhvtEgHiS19BRxxOJCj4DAr0ihUTWcGsOjyyV9L5hC6A23ITjPu6Aa7t2u74+ZueYAVARPkEshCJO1ei5nOVQMHui19PP8GzNe0IBL619CL5zTvqcDMOI+Jw8XgLNPeuWsXwelTHuy/AMl5HlzomySFe3x9ialz8ugaMyPsY5sRLlORzNd2coy6HTUser6imB74b5GC410BpFUUo+z24XI8xIEJDo4BhTZpxyMxgsTks2U+1zLvJVuNYY/hKSGJZ1o+xHKRDAENlkEkcHh4gNSeAPkM2nUGSHWiqLRCJiXYKNlixIN7f3sEMbOyWXsTPVd6fYTfJnfY//eT3v6N45pxIjpM0mjfeQwmEfAs6/kxAlZsb7xDWfpIIsA91hlHuxkVjWSWrP0dZ9kYMa8wPECDe2m3LESCeZ67GP3cMyhpz7TmDFe0rB4+RkAetrG3pm3Ic4pmRHnkhqrWV9TBEP30eC004L+0dHIiqUwSuL/Jjen+u3cn2UrUobPTpupNFoMFSd18ka/7uOim9X4d/9yx/0HZhoNlUY+gXAg0r+wCFQwAXS8oMOBabY4ukB45OgFot+Ft4wH1jbPRzragHR/Cd1EzgSYkxUmH+pbSzOy9QpO32xq+DNcNhaSKsV83iM2kGKE5mbA9dhbjRSh5HF5mbvOipY3HEycxHToU7ZGEZyaAMQWWOPlAvcSGEmNZfZZHkrJ/OoZAFs/24BR/Y6JnC1MCQ7BJmayIl7zB/UtazJZ5qMP4tq9UzbbfOvpc4RWlhpk2IhbPdX5/RwWGw1NzDrBDAg1bckaqNxweFUGkmpTX/QDtU1iVER4YE32V059ZIx9yQoTJVgAEoEzUYdyZQVDZGogQb8HbbX8lmwg6LTozclQXrLruChip0v3MgmF+mJyPtpbXmm1rAWRgMpPEgwtk2yzhRTJPgNXGPCKU18RsULOyrSaURTCTdmGUptYdpGVMTR6bcwNT2te8Ex9NsSFd6nOQj28bn4g5IBlSzejNziM8kXCgJfuGFGBgPMzkxibmkGD+/exvqd+4gNINUPC0Z2tvB3PaOvPxOWn0JWnfZmVADRs1dAQq+Drc1NLC4ti6TguGSxzQPU/dV1eb6+iKhQroDLs3gZIP5fQlQoME3zqa/i4HRGxe/SURFUXdqaZKCs/zxerRoEavgsuBb5wiA/M4e55TOIZXIK3SLYzu6jermkgo1jjJu+gf1Uird1YO53aigf7eHh3ftgrohfnzQJfxNR4Yhcf/9G3RUCfl+M1P9/1VFBooL2T8FnGdy8XtVRYeSM+Wrzqgk6XLl8CRvrq0jE02od5kH53LnzOCyVsLq2IYCqyqweb48WUNx7gO1Vm+cfIlHBPYBz0YOCZifjiYpxBxEBJo7LRDYl+5FWu2dhzf0uSkf7Ip0jFi09+joNfgfvnd+3/V58+nt+v6Y2RMMIAAAgAElEQVSCdsD5LvLEANMgYAhQee+BVAOJfBgdhgxptAMcD4Qszk3NRWCbRb8TFoyIqRd3VNi1mgBAxD7HldvvvHc7dxXOD9lCERBwxD1BPn4paFvHaYdmOetItgb8x//43+Hu/Vuol0qYyxUQlmVTHy30MIzFcOGd72FyfhGLS/P4+f/9N1i9cRMT6bgO35VGFRnaTchfmwTMEPVGWyCd6qRvdVT8PogK/5TtzyBoe9r8ywPd9rmtk8Kyt2ifOcDS3DSK+SxiGGA2n0Mxn0c+nTWBiGxpmDfGzkVTxqezVHBFtJcbyEEiizUIAYsurt+6j2fPd9DmmktgLxGVEv3CxUvIZkhUJKXMpn9upUYwNKraLBaJIRFlfUGioooSlccMB4yEcfvGV3hw9xuEh32kHVHBDI1gzRk8oLeohC+VRe4bRxyw3jpFVNhruE7Zby2vJ2aTM0FQVeuIChuvHIu+o8LPoxPz6hRRoVrMW7vpP+y3RuTHKTsj67qkTZIdiH/z18mfeRVR4d9z3ClhQhffdWh/j+Ly5cvjIGoXqqtOBdmMmtJXpKvzhw4SFV585OsbP17HdZAJizhvCeoaUTFWkHrFsf9937Hh93C/lvm6l+vN7u6O68LlWG2PBCtBoiLfyckCodns4PXXXhdo2O93cPbsMnKZFHaf70gRfnR0jE6vi0uXr2otIxBLMQPrLa51B/v7IgBaUtwf43sfv6/O2zvf3BZYtr1zjEq9JdFJp9NEPp/Ehx+9g8igLeK+UJxQJktEgasZHB6bhQqBrVxhEo1SWaDt5sYOfvnpbVy7sqJ1kGDG+x9+IBsW1myPHz9WhwGVuze+vqGAbRIVf/TD7+Pps0d675mZWd3rZr2Fnd19nFk5K3uKSrmMbCahXI43X39NqmSqRW2BiWJt9bmAX2YfyCI3HhFwKDVpt4upqQJqtZIsW6+98TryqQzu3L6Lp4/XUCzmMTVdVCfUpatXlIn25MlTVOtN7B+WEYrGUWcXWr1hojaJ4KiET6uznu/nr8WrjykeU/cMbZMoPuNZyoFI/H3WxFw/5Ckvi+Gxcpp1Ln+W6xp/38JdrVOA9Rt/h8Adu/74u6zflCdAW98krVSbAns5rho1I6D47z6PguOY10ygy855VL5OCGB/8uSZOiksB5DXyC6eqHbuATvwaeHaqKPTqSOdCuHP/82/xsazVXz5+XXNfKuq+EgiIoEm8jmkEymsrq6izfMcRXk6e1lNQaCVYDNFIeqGiMWxsLikz766uoZ0Nq9zKtd6Xif3NJIVXtwnKx4nqLBg5ogB8xQ7uY4CWmdpb0ilpQTn3JCi2AGTDFYPDejPXsAf/9H7iKKNg+1NNGmbO4zi/JXXcbRbwvXr36DT6+Dd99/Fs2frqFZJXPE5m4iq1enjzMqS6h8C4gTftnd2cfbCWTx9uo6pmWlsbe9h+cxZCWB2dnf1mUkA1QkMJ6zDf3puGstnzuCnP/2ZOmOOjmjfQzIiZZZXzaYU8jw/eovmulOL82zrzxB+/aIjAL+4J5JcVwgvLdZ0xiX5QdcAflbLJuG9JgjJ+85t2c6nIYn8WK7obC77LgOezcrMguL1fbkIuDXTiRW9QJHX4XEJf50GvJrw0G2I7sjMmsm6Ydm5OFXIIjbsY2E6r7pg2OviqFzB7lEZkURc4b+0bYxGE06EGFaWAXPBGBRPAFmiSIpThDkY9sPxzXmkHKo4MRPDOHi/RHBL0MEaj+SH5UVwfCn/gaHpwkGGGHY7eO38It67ekYZFbl0Ck+3DvHN423EJ2dRKM6o02v/cF/rRdwRtRRRKlOi01G3GZ+HnQn7+hy8Bm/z1Om2NG9JunC+006PHUN8dnSKINDLa6L1EzvJOM9ZV7E7gvM+rzWeBD6tp/s4ODiSGJR/z+csDNo6v6yeUmYbcxOVT5DV8+a/U+ji8y1bsiu2esdjXx4j8rXEqP5xIl3vOOIxEuEnzuZIWA+tyJ0LCe+DcDSJTCnMdZmbIo+sC87OcfY/H8ZN0RRf0+osrkq2Jsomi3Whc8HgnmnD1Gy/+D5e5JCMRSQ6KRZyuHj2DBK0RgqH1KlGe7eDo2PUa+x0iYvA4945NTuPzZ1dbDzfFVGhqoOYk9Ynw/tYewtLcPPE11fjc78TLDoSxuQsJEJJMFuwOucN563Z8lkoN9dVy2qz8xDXTH4uj+H5nAt7Luwmzojk6TRrEpoWcmlcunABn3/xJdpU8nB95R4qLKunGoGdX8+fb1vIuqu/+HpT0zMisSk8JdbGuUarQVrblaol5QORnJZFXdKcWjwpyt9nNxOxIO47tMvjWqVx8x1R8ZtL6u9+4g/rDuQbjRNWBP7ApdAdZxnhDy5iGRU6xsBL2xt9W6kKTnYdcKKKZbdANN+26FVYnHT8UjFHCxxu0lwsHfiu0CkGXQcOen5R4uLBxZ/FE5lGhtSQ5SXoS59XKRNIgii0xjYsvg+vkay3siQiUS0YVrCZIoegiw8Gt/c3D0BfxCjHYKT2N+Vk8J5oo6b6ggFULjxbZ1kFGvF1nH+eC+XRYkV1vNhqfVBdt4K3SQKFDWC1cFo4sLk18sjk56HyivdDrafNBrY2t/R3Kn/Ygsdim4ssi0u/6Q3DDCc1PxpT9dnb83Nyo2GBlYhTHdIeqRKsuB+rUxQAxOAoWj50Os4LkMA7NzcqQ6zDgSA1OygYYqZgJ/ffUoEtzepz8noti0OnJ0dUWLeOf+aeKDMCyYApO+ha14zf2OVZrs4YA71oH1YvV6xoS6YQS6b0uryvvpinDyLvEwMQ2Z7N165VSQ5YQeoP/R6k8EWCP1gHVdX+sO5/Vr/vQTRXjMYSceQmCiKiWEBRkTw/O42VxUU8u/8ANz//HNlUyronFNzGsD6OVZIRHA9hxNJRlEpHGv/cyDi2WERzXNOCY2t7G7MzMzqw8XsKOOv28HhtI0BU0DnShZL6cFLXqszPcRoQPU1e+DUiqFzzz2u8+nEisnC1tlsBYY59k1EKi3YX6HsaOD8N8JwgSk/Z87xstZXKRtZuEczOzonVmz53BpOzVHSkVZxQ1SQvyXAIKRGYbBF3RVenh26jI0/p7pAt9mHc+eYmWvUqQlRvyDvfhx17IMmFEI+sXMZA7WicBi/YAV7mfX7qk+h6fvuv0br9ivvjiQr/qqef62mbmSA4JzCZ4DZJYBLF0Qheu3oVjx7eRyGXw/mLl8Dg2+LsHG7duye7HKpKD3Z21GJshKShzKODoQ6J48/pi07+jJHIJqcM8jn6nAo0sHL72+Pu5D0LAnevAvpf9DrB633R747uD9cd1x2o1u4I9zZnNSXUk+u6Fbr67KGIFGoMfpMCx3XI8fMT3KAS2KwXXmyJ9dt+5uCdGBN6MQWH2vURJFHbj+6pWR+aukudcSSFKQTgfB0OsDQ9gddfv4TZ5WV8ffM+vvzqHvryZe8znvLEjbc9x8BKHVoD41sHKJ2DePA1Oyc7EBtHbSGf7DC0n1FPpWvNpq+uxi3Xf/9z/J62W7vnxclJzExlUcgmiTbIO77PTtBQGBffeBvFM1cRT2YxN1XE5tNH+M//2/+K6UwMCfRRmJpGs9fF7v6hDpdUfPUHYfll8xrsOm3MqssjADX7+eQ7F0/cEAZ/B778fOXeyn3TWsUNZNecsA//wo4B/zJG9PDg2Ueo3xUAcH5lkZ3ziA6HKOaymMwXkM/mBFjJrpOHbh04zc+W+4SUpVQxu0BK7tWhWBLVbh+/+PJrPGOQMdWfYdrTnMGHn3wPxakZ1RoEkLi+0/qp0eKBy/YjgWVUtQ4h/3p2qBAIIzHx689+hacP7iM66CJDMFdK74h1BVLRR1FHJC4yigo3gl0EBet1y6mQrYd/BhRfBHKifK2j/fclHRWj5xRYK0/Mb2f95O9zcJ8fzT1HPnyL+nhFF4fvtvDPXvPDqUGt+dYO2149aO/vP+vJDcLPZ6szTn75z6eG5jBrcdbB44wKTh/uiVNzC/bqriOUh3jfUcF9z39uv88THKPqmXUIr9UTDWOgz+b7OMrDbGRoUWTiJQMDbH3k2LD5yjo1SM75eeVFKDzE7x88HwGvAoKceMqCgs3iJ9NMYzBgFkIaU5NTUrvu7jI/qYLvf/IJZqam8J/+5/9FNmdU///lX/2FAOGpqSkpcxl8zC5BBgIXJia0Fh8f7OJHP/o+Yqk4bn35a2Ryk9jcPkKpUlPtSFFOJh3Hxx+9hVi4rw5M7nsEsKq0kuwPMHPmDKp7B8qGY00yv7yMVr2Ju7cfsPrWWk+wWyGZAjt5D6kSZq5ACyWSGpubembNWhNvvf26LJlS6Timp6fQ6dASaYD9/UNMTkwJkOd8p9KzfHSED957B7fvfIOllSUcHh4jkUxL7U7wkTWwwJxUXGAbASXaV83OFJErpPGLn3+G+bkJLC+dwfvf/wGOt7bxkx//GFOzUzg62Nc8L05NY3p2Dm+8+z7u3HmAw+OKSAsRn+GIbJKYY2eKUbPkrddrqgkKEwU9V3mQOxsgjlUOTBIIBLA51ngmUXe860bvdnoC2FkiKGC33dbrEgTnemFCNLPcVYYAhWzNhtZI/jfBoUIhr1qflkW0NGGnButt+rPzeXz40ftYXlrS2Nja3NC9ppqVz2RpeUVk9q+/vqG9iF1l3jOd75FJp5DLZpTVQ4JmZrqAQj6G5YV5FBeWcPvzL/VaBO4iCbP+onCr02wjnUxbTRDjZzFBH9dpBmczd0Fh4QzJlTo/qaBeXhPHWq3elIBP9jzKLAwJqB2Dj2ZxYmcZduMNZWXCXAvmFWbTGREbAh/bbZw9e05nESrGdcYjaE/OsdfA/HQKP/joTUTRQbdZUxdSt8PA3xBufPMQe/t1FCZTuPb6a67boKvsqGw6p+wnZlVwvFsns50DZdFUyOPunXtYWlnBxtY2Ll25qt9jZwvHte5zpyXyip0X77z/GmZm5/CrX/1Kam1ajrG2597NFyWZw3WLVisSxfF8ymynHjNAjHAguc4vA+EjGiPen5/naZ2vOh2NX1POG9jpaxVZmEkASXsYqtGj2r/4uTgWZVWtfAzDGwQVuyXd9l1/HrM6kc/f1jkDzS1I21TsEkiO8qRMsGWtR3QzMFA3Hg3jnTdeQ6dyhEQEKO3vIptJYnZ+HvNnzirH4+effobhkOp82iQxyDyla06mUyJZ2O3k6zKSDrwm4hzWpWIqe+73shhisG+D9uDsELGakgQI55JChKlOl23sUFk3Eqr2Ojg/X8Qfvf8aWsf7OLu8hJ9/cQtPd+uYWjmHHWZk9Luywml0WghFKL6Lod00ZTlFhUdHh8IieJ9k/RS152N5qiGcO3/G7MxbLewfHGqs8V4Xi1PCTaRGb9bNSirMNacuYQX/m8AvyQyuFRongwEOj47N1jIaxdz8nMYFX4dZMdy3+J4cw/xZvob20CFkDaUpzetnHkVAICTyirhUz1w5/BkpuKsH3UW8Mt8TE/yT65Yn4WydtOfFMxRJ4PEB07AmZfgwjF0dO5Y3apmyBPdTIinNy2So+2pYGbNHWmaRFjVcgZ+Rz4JYz/HhgYjaRrWh+jMeCSHUHWJ6KokrFy8izfUwzeDnHnZJTGxuoVJtIZVNSThYb3fl+tBilwazzxQcbtfnxYn+/nhCwWzrrIOHd84T2fx8xPRoi8R8FD4/zisSMfx5I7PZlcDQeMMk/ZyTBZrrNDNIiVZ6Vg+RJCV2l0lGkU3EFVhfLEzg5q1bqim6Bm7Y/h0JYaIwoS49vp8XaLPe4lqfjNPW8VBkhbr6+n0szC+g023j4PhQ488OBmF1PdFCMs2uEJItQ5Jy7Pa2vcpIaSMwvyMqThXE3/3nH/4dmGy6gweBeG+tpIlvE1dtrJpEBtwbkMBFIQCuuXXQWmq56JFRNjsGa8VUyWpWDkJszAaHagQtum7zZgGhQxZff7R4Eiwx2ygyo1zoCZRzYZ2bm5OfrDwDWXxQfa4N0VQKLCp4QOJrUkGlhVttvu6gI6sL0zVYK6e3H7CFW50TrvPBWzH5YDgPsHERZ/HERd5AT/sMXOjoyUiG3QM2IizUhmc+yAbCOcsKgkMKqIrr4OjzQfja/AUD3C2kjYsww3t4HxR0Jk/UjjHPPVP8cAPml5E1MWsxpVc6q0xuXgT+1fEx0ELKe6ICRz9rShArdltO0WHAoZFTfM2E/rSsCbteqaDCA3R73NioMKEayMgKAdbqiOijuDTjOipIVJg9hBEVfD0qqezo7dXxniDwKpOXExXWwUMwlSA/iQoehpLJNGJJZlQYUZGhZQUVV7QLYDh7i8q0GY0FHh5GuSQOPPIghidN/KHaX18QuD9NVPBatAGywCRRMTkhYI8HWt5n+vwvTM9gf3MTNz6/DikSEjEjz0gycdOmfywPXPTXTTEo9kCk1piosNbANomK58+lBuSh0Ns9cGysPt9Go+2tn04TFQ5ADeSgnAbVTv+3H+dBsPskmKtE81Gnke82UkHwOxIV/B0PdJ8GjYLXFbz3VpTYepHN5JDMZDBz/rzUiZzXVFQlYgn5Ges+txn43hV+yvvV5iGnK5McDKJD5HJZPHpwD9vra9TKKYgsxJZwHTZ+O6LiW7uFA7P9PTxBHPyORIXUhwFy7UU70/8rokJrtBWDUYLBtA85cwYP7t/F4sK8Wu8Jt+4eleTfzZC0qekpPF9bl1f2qGvO+Zpr/IioHQNwvtXWA3Q2r+y/vKWSB6l9N85v2oGDRIUHvk6PGf/fp8mI4H+/jKhwC5UjKgI2fW7tUDfb0ILf5B/K4L9oXHOXyhuzYeJOaW3BDGetVSquA+/ln+5VpMuLvudB8Eg4JkUtx72ts87vVUQF19ywbAnpXBh2YXtzM9N4/dpVXLtwDpNTOVSadfz8l1/jV9fvYkDf3yFVckEDSAPdffFPOyF1850Aht1KwNwB5Sv4vcX2Y78vu9ZEpwKzwG2Nc5IsAXKDbexSfEWiAh7PLEwin0mhVjo2C8RoDNMrZ3Hu2psIpScRjaexODuH8sEu/vf/9D8h3m8in4jIiovdAzzA3L17T4BQudrSAUDr/+gzBDNPrADSPXaPzHdMjp7gS4gKA6atW9Hu2SmiYszHfWsweDWbII4BbR+juHDmDMK0g+q2kU+nBZaRUJgpTuneEJRj3cBagnsfD0MiKRTm6eYafz8aR6XVwy+/uoG17R2Fm/JZfPi9f4X5hSUdjvi6CQZc9gcolY/RaJQRT3D/SqqOEVHhvMbpr0u/boZnf/HLX2Dt8UNEhz3kkklkknGpY/k7BLDYfSElW9wOlezUIVDGDpcmw2VFBDuC05HdWoXdmPP38jRR4ckz37H5snXAZ1T477+QqHCdL6fnmubVS76+TVQYIC3bAQcE2Xg4SWrZZz35ui8jKoJEjWEe5levjDTZ4Fh3BYH4heUz2ov92qzMMZf9NuxabccvDwbw+xRInCYq+DO8btb/sotw+hteI8cagU8pBt3h37o7WKdb3XGaqPDP0a/XVHweHu2aR7QLrbW600Az1nT8s9DJo1ppIJ+zcOyV5UUUpyZEVhwfHWJ5ccXqZoGTIQt3p9rWEcisY+X/HAnrz06nhWrpEH/553+mLqPbN27Kf/8puxHKVVmI9vvsxkjgg/ffYqqLvKM5bnVGymZRPy5b4GcorIDsTqstu0l2pt9/8Ay1OoVRBlKWK2WcPX9eQinWi0+fPdOZZG5+Ht/cuoV+d4BcOouPP/4AN25eRzaXwhSzFCIUr1Sxu72vDgsCzlQdrywvYdDrSKU/NVtU1xNBVGrFNjd2FZDL9U1AaZikYBS9Tk9gXXEyj+JUAecvnMUv/vlXKB0fCnx98/U3Mb8wL8urjfU1HB8d6YgUpc1HqYpkmvU0A0DpMGXPhtl3JCZ4xuBYpzCI5z51srtuC6nMBwSXGwLEvcKYdbp2Bh0fQzrjcR3zNr18hiRAaVujgFdmoHCtcvlHBNF4XiL5RIBneqponZ7Vqu1z0bCU0YN+T2siQSOenXh2JBDJ9ZJnMHabUBymcaGMxayIJamjOZYVoEoxjp2V2xQAkghQXl4HsUgfZ5eKWJybxbWrr+Hu7bsKxmbHBP8n4QzP4J2+PiOvodXvqU7l2ZJjn10c+wyWHkIB1QSGE6kk1tfW1dVSrdXR7vYwQxtbdpeQ9HJdxcH62a8dBCkprhOQ225bDh474GiFKkshCtfiGov+Z7j0djsNoNvE5fOz+MEn7yKGDnbWVnUOjUSSKM4u4vioii++vOEyuBaxubmNTrev1+r2QrrXJJbYgUuwzsDVMI5KxwLTV9e3cOXqJTx5uobzFy7qnu/v74t0YQ4Fz4nKFKnXUK7UMTGRx+bWvgBqqrC5hFowN+exiSY5D3kfOV54EyWUU1A0r8lZYA3tXhC0N0Io4uxXLCha7gW9nsYB90/+LvctczugMNBcFTjuuZdp+6YgU+9h4cACLIMByeR91HUfso4fZ/fM++/zDr2dEF+ba53U2Qhrh1V/qQQcRlRwvOSzGawszCpf79qFM+i16qhXatjaOUSz18aAXSnNnrpOCIKmUxnlaDB4moIjhRGzI0l2QSb4MqEqgVoj/4gb0MrRhIskzszeV8Shuid6I6JNKnaKX/i5ab816CEWGuLquQW8fm4ehxsbOLsyj8cb+7j5+Dmys8uIJAnOVvWMQzHOEyPnuI5MFAoak+VSWecI29cofDWSSuD2cIiVlSW9l7q14kl1I4m065tYlH9XDSxxKLuLalqj+ZlZx5BINZB5KEyBf2os9Xpa1zj/uBdx7bZOal6jvQdFtXwNEhncA72lnJGrltd6+nziS4cTZ0GHhWifdaIC63C3L4H3IoFs7NjcdXgKSSNXm/J9OeeVY6dOXAPemRVkXaVmpe3dRvizwhCU82PZUtZVZBgfx4as0GibmjFhJM8NmUQcGXbKJmISCtUqDYkWI/GwrAbZOTY1zXyPrNa9dqeHR8/WsLGzhy7lWTwb8j5K4GZdJ+OzvTmyONez0ZnXiya4pejzE5NyWbgm/LRnpufqOit0ptSZzNw8rDvKanB1pbhCxtdU6uqQQHGAXruJRBg4t7IkMpri6XK9iUbb2bg5K3sSXbxv3Cf9fZXFXjIlsRq7N/l5tE9FIrKAYvcj1/mJCRIQlofCOcoamGs01zTDwIba09j1U6vR7j1luOV3HRUvrcG/+8Yf6B2YbltYmbhTl1VhbWMGYNgiZ8pGFkj+ryIhvELaqxxdrgMPMhayMxDQLaWmIx+UHyG1lmtnldXAQMUZ30MssTscWZiVBWGzkBE5oKwdayPXwumsgngp6jBgp8SAC2hLG4nUBk7dLs901745+lyuOOA1SZ3mQhT5d6pVWHxpgYuEFCjG1zIvSgLNAxVQVGJxwRazPehpYeHnVbusDxznJiZ1O0OmE1LN8E9uuGSvpapkmDPbpTstWR1w8WSoG6+FryX/0P0DbdQqdBi6Jz9BhqATbOhr0yEj7PMneB1cBFlE8IBA9po3mBu+Ch4WWvGYCiXeY7VRymbJWlV5LQo+d96cClPnxu+ICiNnzEpEuQsxCy+noQeBTf6+LID4P+el/SqiQl0ZIQOqThMVCgx195X3JOhlbR0VY6KCzH+zUtWYoII+mhgTFSkebhxRwda8RrslooKvx6LEPzON/gDgdhIIt83Nb2IeuA/+jH7fhdvyeXmigtfKtn0+g8mJAqYnJtCuVvHVp1+oHTYcNtCNOxhDULnJ8nAmz8tYSMFM/GKYtrzAncqFHRVr62uyl+JmyOfL/7HAfr5/KCLDDikniQqv4h2TbN9W/wYLqCBIElz2ToI2RlTwmXml5uhe/o5EhX8/PyZettT67/vCOhFnQCLzPZI4c+4c5i5ckvKFhYonCFnY0vKh36lrbaA6hwcMduQMOlR+D+SFT5XJ/u42Ht+/Zyqf/wKi4sT98Wpxr8w9Ha79/yuiwrxHPVERi4SxMDur8be9vYWLly/p8NciuLK2gXa3j2Qmq4DL7dU1AR/+GQbnjE4HAaLCA2Z+3mk9dvPHk4P6N3N/CYC7r9p8x2oiDwCOO4HGvsR8hdOgo3/vF33Pv6N+h11cTnETfA35wXItUzcK13BTA6bTWUwVp9RNQb9wT1RYwF0bz54+NQWQCyJ/0ac7fa0vn4f2HU9U0PppGCYA7Pd161Dgs9X2OuyBzzcVjUuRf+XCBVy9dBnTBLq5Fkb66IdC+MdfXsc/f3pTSqge7GAX/Dpx0OLYDhAVXjXuvcN9vofNX2tP9/dcRKBvXOJBK9BREbQUI+jE/Y/1BQMOX7uwjN2dbR2sM/kcCrNzuPzOu8gU2TERRTSewsLsHBrHB/jZ3/41Nh/fxWSaVgZRdb1Rncx9dWfvCOFoAsXiNO7fvy9LhOBa+LLP/K3n8wqiwkITjZEwAYQB19bqcmKKnLjHnsBnT0FowMDaOM4tLyqQfdBpI59JC0yg8nFxbl4ihEqpjGqtqvlK+wTufwZAc+82UYdqiVAUB7UmPv36JrYJRkbCmJ6ZwV/81X+LRpOH8JzqFnZUMCizXCmhWi8hHrcORilURShYKCpBNNo3EJz49Of/hO21VQV+51MppBNxpFIxeV+TCt07OJA/P5Wd8pgn2adutwF2dg5OEBWy4gqsnf7vWidOdTf4w+xpEOBb8/u36agIEBUn5rx86V/89fsiKvxn1Jw7RU57cN/WOF4Hs8EM1DerCLNAYI0w/yqiwlkOeOsnvifrIlo4mh/4uKPCwJsxUWGWpMZ6cR1jTcV92HLjrE4XaetIuVcRFbZuRnBcoh3emKjga3miQnlcsRjeXX4XTx6tCiCjMpw1eig8QIp2sM5mlRYJZVktMAvBsiDMCsisPaiGVz3c6SIRZzD8EP/uv/5ztFp13L55C1NTc1hb30apWhdA0G7zzxTee+c1DHttqSgFXvEM0u0iV5gQMERQmV7Us3MLGNJCpzvA9V/fxsMnm7h6+YAVRx0AACAASURBVIJq7b39faysnJFqktsKbXB4juIz3dx6jnw2LxDt3Xffxp07N5hfrZBvzrFatYHt7X2cP3dBdSLPTQTMKgzGnp1GoZg3gENzPIatrT0LKZ6Z03vk8hk9G17n+toqzp8/g2erTzE/P40333oDu9t7uH/3Hg4PKjizsoD5hTnMzc3ovLG7s68MmQcPn6Afoq89P3tfoJTZqDrBlBeFOCtejhmemwQiMeNoGJL1DNd/1mzyo6f9h+pYByjR8ihBa7moziys7Um+aMl0PvQGpI59xzkWuQ/wDMdRKQ/6mFmZcK3ja1hGn51h2H3BdZ4CDIXSMmidwLazY1XnRzis7hR2i5GZI/BI0I0CBJ3V4jGR94kYuxQHCNFetpDAbHFKZNLXX91AYbKIequNnf19VFstWbbOTs9ic31DZ890PouNzecaG+wsk5NAp6cw4QQJ5sFAhMaTx08FivI++HOwec7bOd4yFkyU4Al31QSsTHjGYAgrO+WZVzkYiIDmuZLnS2ZUEMBeWFjAweEBBsyFGnSMqDg7h0/eewMx9FA63NN7ZApTIsBIhN1/uIp4MooPP/xQljm0BmU3J60CibMyj4L2obTP4vrATsgHj5/i/KUzePhoFUtLCxr3V65ekyCRIDIJQ56Zl5bmsL+/qzG9ubmngG0KtCh849pAO6nDEoPj03SsVDahQniZj9Ft67VM/JfQvyl03Ts8OKcFjj0bRwRpzarH+/xzThKg5+/KErpHcimje21daSHZJYucI4bALAy3VnN8qqvFCXDUOcGwaZc5JKGns5LS/jcYqhuI16LrpJ0vVdXELrzIxSmvlUVANX86halCDp1qCZO5NOaKOXW80FHhsFxBudHC1s4eLB4jIqKCn4V7RSqTRqPVULahCEet2eZAobEcslBs5kwQ6KY9HAkvBsSLBJASjQQQnRTozMEut5Tm0YDgM/cKdrl2Wnj36nlcWZlGq7SPM4uLuHHvGe6u7iM/v4L2gLkAVeEJfSrIUxndC9pWW4ZgT6SaD8ZW52CUolHLaeNzmZmdUh2tfEyFMNM6kJ0LRmbRZkcdBf2uCEtPhPAZ8j0y2awC0vnF73G9MgwiprHDOohrBYkK/rwkR8o/IGYUkcCNJAXHAW+LMAsRC2NCanweMZD9hV8OTPfnVp9TqnrNZU9Y7WhEinA24kT8nutaF0HhcuxEmAUIGgHiYeZjWmC8cDgSx3USLLSAIslM8V9Ez1J1hvbxiDom1XUxGCKdjCPU6yIZSygvbXluFslYWLhcpV5VduHxUcVlxyaQzuUxPz+D9efb2Nw9VOeu7J9Y/4p/MdLFukjsLMfPwPe1zlP3pegPO9Nw/vB3iIvIfst1P3P95pzlMyCGaI0mlmPjRbuyceO4lUuKWbjZ2m9ZNRLkdlpIxqMI9Tq4cHYZ05NF3LpzR+HgXbr1ySKepCwtFKf0u7u7u7pQn5nDscj1an//YOQ2wX14crKIZruOo1IJ01NTsk80coWEl3USjeuprsYex22jYR1m6iT6jqh4aQ3+3Tf+QO/AfM+Brdw8gopq5TSxsLFchHy+YIFclbKKOh3uAp/ZA/wGKNmGLsCaCy8LRapgaB8ggN1awPmzAnrVDm42AdbVEVJh5g+UfF8uKCOFFxcpF9BGUsQrRwhOsy3QFGq0XTJ2nwsN20G5EBi5YZkB1t1hizIXeykaeKCj0oLFqlQ6HW2w3IiXlxatCMjSO85Cl3gPtp9vy36KCyHJEBZE3subrLDaTUlwaME1b0OSDiwMuWDyUMUDjvmDAPkJ+sNWZePDg6FXgCzMz8tTX5sz28Lb5n0p4kP+dFBbIe89PwOLfRXlVHiR1HC+1PLL9M/XMf8WemztrGSixbbzwMZWVimNas6vc2B/J6jg7LD4c+bvx82YwHRDAF0qxWKijU6PvoDmpc2uisnF6VG7rVk/GUAj5atsMGxM+k3b/n2cX+GV1/77Bl6y6DZwn8BXs95Aq8YihDYraUTijqiIxZBO53T4oZqE7fu1ZlObBt/Hb2TB6XwasPTjMlhUBIkKHQLcNdHrml9svxxZP4nU4YbZk33Z3NQ0Bu0OvvjFL1E+3EdIbazWtsyDDzd5FspSBsQiCkvkfMqJcGFHDZWFcbR7PayurdmhRc/f/kfl1+5xCV2Rj5yfY6LCwI6IswKzOfmiYulFYJAHJz1Z8yKigp+R99SDRH7dEHDpfC49qHF6CT39nqdJIL3WKaujEWgSppc+iQoqo+L44MOPkZmZRbXWMBWGiL0O6o0aGrUaup26tb3m8yrOReY1W+gxzCpJ384Wsukkbn11HU22+cp2xuarB9vHIOPYtz64Sp4kKgyEHH/GcffAaZDtRcDai+7Vb9qCqGQiIRx8veDfT2ZUWJHoF3oC8VyiuLTSm3ZhftY8Z3sdXHntKvb2DxSeWanWlYGQzReQy+awufpUIZ0qsB2YPRovL1AJn553/hl7/+DTRIV/TU+q29wbZ/z4ucg/R8Cu2+f8wXE0X19gm/XSg4Mn9tUtSKDY1iz/2cbPlTS876qzNuVMOoscD0XKI3LhnxhoLSCx+fD+PSlLfzui4qQlzKhu98/O/YOuR3szMyqiWv+tVd26ZCxYlKQuMJHNYmVuHueXljFXnEY+lVSbMpXsw8gAg3gYv77xEH/z00/RpGo0bGpAmwnO8k6yJ6rFiT9Zt4CthAYWWL1gbfFeJGHPyNZxHYodkDIqNLhvSU11iqyyPgTLznKf5dzStAD0SR4UMjksX7qM+XPn0Q3RxqktYGlpYQHdRg13v/41PvvZT5BjwF80pAC89Y0tXcvM7DzC0STOnbuAf/zZzwSY+K/T8/LEXDq9LgXCtINguv2OgUg2ln9XoqKnzq7QoItCNoWl+TkBpsNeR964tPVgXVKcLMpygaQs92/WALOzM5iYLGoec30jeMvDGe1G+uEYnh9X8NmNm6g02wjHuYa+j/fe/x62tndVDxLQYkaFiIoqCZAj+YwTdCJRYR0V0JpAsoIHe/YQ/eIfforDneeIhwYopNPqqEilEzoAc588PC4JBCRgIo9wUJDRkZ0MLeVo7+M7DEhU8Ct42Pf392VERXBNGM+XQDX7CqLCHuv4PYO1ga7jFUSFMolOEayjdfF36Kjwn8+vfb7Lx4A0A1G94o7KYwHwrvOW18jah91uU3OLmktesUiwQbWWvEB8veUy1wjicb0/1VExmgus4WWZwnVmTB559TprMNaYvtY3j25fdxjgEZwXfr020CSCUtkO9F5cEyQqfEfFYmwJc7OLWH22Zr7bPZI0HSTiZmlKP3PaHvHpcWdjeDUtfOhNrvvCse/UsFQkK6S218Kf/ekPNW4fPniAyclprK7vyG+fAcnMcZicyOCdt68hGaei2e5nhLXzEDg4OJSYaeXMWXUDDSmA4DeGITxd3UKrYwpWdXk2Gjh/4YLqNX7u5zs7soggSPns6aqIHc7hjz/5EHfv3lT30rnzZyVuatTbWF3dxNtvvY0vf/2V5uBrVy7RBxeTE3l18U7PTMv+xIDkHZHk9SYBjjTCzJoLDVE6LmvNnp6ZRDodx4MHFGZE8cMffqz8iwf3HuKbb24o0PjgsIrFhSKuXXsNs/MLqFQbuHXvoYQKzB/g54owP8KtzwKNef6DZcGRJPXPnWcZjgmSmY0Wz1JxjRWOVa4D1VoFg57l2qkjXkIe22tkreOIJv7Jcdxq0qrFbDw5FmRRLBV7H0neU1pmZDKay7xXtHsxEAmyGDp79qzGMkVoVO7zq1wuac/kOuZBfD5KjoV4Mi1bGJ1pZTXTNDELeBYMo5BN4Mq5RZHjtJ1ZX92QmndrdxdH1ZoyA2i1w/MQxUfsAk9mbazy83BsUHBEAJR2IiSz1IVTLmNubh6lY+aCrWn9pMKXda+ppM06hecD/ulrUFt3DEDm/eFZVF7+4fDIRpgkN4ExzmEJ9oZ91NtVUNzeqpZxZn4SP/joXeRzGVT2tlEtVZDJTyCfn0QoEsNXN25JwX7h4kU8ePDYAse7A+TzE+ou4jifX1jEk0dPBOgS6N3a2cHSmWU8397WnLlz5y6WV84IQK1USjqPzi/M4Hs/+AT3797G6rNn2NuhrRo7HNgdFcIc86cWl9HrD/HXf/tTkUbsoKIFlOX2sZuXZzDuKXU9S+at8H7wvMSzLW1WvMUTz9v+zElQXNY3MRMhck0TKakuRetO5Nk5PzGpMWPWUkNT5avYMSzEdz6oxqGTgHAYW02tg8388hUMTEcJ56GvPxkYre5Rdt7zJS1YXpuLyxeLhIa4cuE8EqE+osMuNlc3EIsMZGGXL04jPTGJG9/cQTyRkeCAwgCu3+y64r4ZTyWUmWZe+97O1NZr68K1So9kheyhZRFq3Sn8eRJpppYnRmFkGNdjdRmRUCDA3u3gw7cu4fLSNCp7m5iemMTTTXZU7CA1PY/C1CwOD3dRKpeQSCXUUcFxSnKGZ1y+D58NhZmym+5bXqhshgfWBZ9OJ2RrRxKDoC6/z5/nuOfPNVv2nJW/lkzoebVVYwwt4DieEBYj4iORUIeV8CmtKZbXwbWbc5P/ZniZBdWbVVjSiE7iUR4PE8DvCRUPujuh7AvOIL5e8RZFrox2Nor2Pgaqm404MSzhXy77xCyhfKYj1wDLVZGASmPerMT4ZLkOc5jaeSCmOUmsiveP452der7ToNnpIpdJq3bkus3uXXaDU2rcI4k3DCFJu3WEkU5GMTUzgfnFedlpddpdbGxsYmNzG6lsVt0ItVYHDb4Hj9VyFXE5eupOsOvjGVsYouaBEXfm+OJsv51gwtcxxNzk1AKSMGnDUVzHnRHhZsnm3Tq8HacnRjwZIgt5nWlYJ4S0BnbrNZxZXtTnZs1B26phKIrQqOOJFpuzum9Hh0cjYYVsnxJJvffR4aGeGwl/jhvWuyQqjsvHIj5JFKn7fkCyqKP1+LhU0nqodWPQl/0Ws7nU+UdB8XdExeiM9t1f/oXcgQXuRu5LAL8DdDi5uSESsPfEAw8q5vdp9gTGYLrWdQcqcOHgwuZD0mJkvjvtUYt5EBzSgiPQ3AgCXon50tnfvSWBV4mJyY6xm6FtbXYRtuqZ0oAehDxksMClKmpyYnL0c1yIqGhQseEAdW9VoQXPKQksq2JgbYskKFpsaSTDbCoMUxHQ49uKUV6PkQ1UG5CY6ZtaQJ6BZkPh28185odsk5yFljYMX5iw3bzVUDGTyeWMJHDEhdhxp2QjU63A6y7ZVGsvpPqlXK7qObGw58GIKyoLEPoBqsWai3nHmGYW69YyH5Vy3NrJLGTIe2qKAErE1UbO76s1WMUvixe7l7KTope6CicLyrJQIOue4GdttfmZuLGw6DL7p/xcUa/DnyVorhZW+mdLAUCyY9wSGSQpDAS0Qk7X4awJPCnAgslbP6kzxbHRLOpp86QiMRZXy74KTgLZqRQaraaKU76O9z/2xUFwmnvyxAMEwfc/Df76cU7gkV+y1eJmPlGwsECFVHUFGBQnCgj1B3j24CGePnyAyIDgPoFKiIASEeGABh6Ad3Z2pKri92QVRnAuGlVnyNbONvK5nMaFf8Z8hrTkIdtvB5SxmtG39Pr20JeB4sFui9NAiQdnTy6J1lFhrddGbI7uqbNuCariX3T/RoBT0DKGL3LCQiZIl47fgwUmlessCtgl8cn3foBelFZmVIWyGK2j1aijxeCq42M7jIaAXLGIniN0GtU6+t0+0rm0DrZLC3P45tfXcbC3i7C6e5y/vw/6lfcvQQi3Po5ASLuuk0SFtYT7r+ABUmPnlBr4Zc9lDIi/eEMKvm6/Q6LC7L/8+BwRbC7Yz7+K73zQM+P/qZ3YlLIcXwzTLJeOMTFZQHF2FndokxPmoUVySRQKRRVaz9efolopuYOWs/YbDQa7T35e+Y4K/1mDJIH/HAICWAgHlEfB3zv92fx9N1Kca0bQZseeycvubfCO+p8JkhGjvweICv5OsLvA1r6x9RPXHVqREeilp3SXaj/tscDM9LTG47MnT7Qes8vh9Prz7adse3ZwbBlR4wOCx3NC/t7MIxhaBwUPfNwHqTgmqJ3LpTE9lcHM5KQsemYmi5jJ8+9RKVL7wwi6oS4iqSTuPtnEf/7xL3BUr6MfpgaK8if7LKfJHbs2I+JOj1d/nePrp2LKDiICFJ0aVPsn38V3cfJ7ruHAOYMY8eLeJ58J49q11zE9v4y5pbPI09+d4oLhQN7Yu7t7WF5cQj6dwv7WOj77p58i1G1KMUZve+5Ja+sbSKazuHDxKubnF/Hpp59ibX3dkTJG+o4O7W4cexDbt/n7z8X9z3+ZmMPb3vDzmu2E72zT67qOCg/EB8f16DVdkCHYbTrsIp9JYmF2RqQFAUp683KusmYhCGXWYn2BMASN2EXIQ6MOoPQ7d114rXYXiCawsX+ET298gw5t3GZn8Cd/9ieYLM7h+fau1laFSbKbszcQUVGrH1tGRZxdHAmpW/llRIV1cQy7bfzsJz9GjR68tF1J0fopIb99KfUA7O4fYP/gSLljBAtYZ9LrmrkAFkM2tkLi/fEZPyPhi1/fTq2hp0nt4PPwe7mew6kw7ZeRlf79TszJF2RUjAiFF3WBOcs+8ygff53s/jhp/RRc0zX33a/5Nd0sKHjv2fFr3trKq9Ih3jIDaGuTLUzpEK9abjAwNanLlELvJFHB3+X32VnL3+HXaaHGy6yfaLNDMNx+3gd7f9v6yZM2/DPY/ca6u1I9MsDUXauy5Jz1k3IQCDDWM+h3h2jUmgKj2U1B5TzPCYhaJxsDfwkoU9nNjh2ClazRGZwsz/5eT50SVQJ29IePAH/1V/8a8VgIX395Hbl8EZtbe6jVmihM5FGpHGJudgLvvfsW+t2WupbZeXRcKctuNDtZRFlqcAIOOQVlH+7ui/j97IsbeLa2JVCVmRb3HjzBJx+/LxCagPSdu3ekBGdterB/qHMGIZcP3n8Hd+7eRDIVw9TUpGrLcol1TBWXLl7C8XFJnWHMhmrWajizsii70MWVBeRzBVk//fr6NwrqHiBsodFh2p5WtYYS8CBpvXJmAds729jb2UH5uCzQ5aMPP1adv7m5gb3dHQH8yXhKwCs7BBKZggKQCQyzo4JnOW+7QTSVwivmEtBilcARzy7y/+92tSaZQKylcwx/RjaAIQJoLYXPW7f/QPsRxwnHpFkvmYqCgI/msssv8mOe9bZEWC5cW7kgPBcw7LpJsDIpUJXELufXmTPLuHTxgkhr2v3Q2o7ALBXWPDPx3z7/4gtsbm0jkytgGCIAxiDtuOpL5s8RLOaYoLAlFmKocQ4H2weYn5sVUUPCd3JuDo1uD+VaXUKiH/3oR3j44KHyLyLxqAJXFxcX8eX162i1uhJ/sa4i2aGzCm1lXYgxzwIcZ7xmqrgpvhJIXiPx5fccRzxKGNbTudm7DKjrifPK2yR1mCVCWyWzUmvSHhUdZJIxDNpNvHH5HD546zV0G1XUjo8wM82cP+CgXFMw/Ob2rp7xD37wR3i2tiFSjIAix0WlwuyCnjIwnj55qj2KexXnTXaigK2tLREOFAYsLPJPdtKReGrh3Pll/Omf/isTtXHsH5c17ymokz2PlMsp/PPPf4nHT9a19lQkUDJ7MZ4xuU9xXvGHpZR2QKzGFgOlu11ZO3Fv8esi77Os50gsOmtkE1lZLgHPaQTDea9l9euU1cwXUUA3awRdHV0HCDKarZIXaXpLG6sHfWajszFy4cYeC1E+I+1E3RnDrICUnKfxO1mwAO3K/g7efeuawo2rpWM8fLKKw3Id/ShwWGpZaHw+h2iENsyG6ewd7GPA1yVWIktsZ0cpe2qK4oyssSBmc5wwLIMqfqtzeB21Zktz0mzIEqo1KcbUfODnRh8fvXUFZ2ZyCLVqmClO4qvbj/F4p4JkcU41yNHhPsLRsIgT2smKCHDiUtbI3FuURejqTgkee7RxY9ZjTJ1i4bA5bMj21BF/ZnNIsVoXqXRStQYHgzqZh9aJxLMjb4MnHzineG+TzOVydqUkXTm+fEeF4QdedEI3C1rEmVCLryOMQWPDgGa+Htcl/t6LziHBmkVny4AuSSB82Mh1XquIWNaCDp8yYQCxFcOh+KVMNAmBeDJh6DjFSRQhWScQu8n4JVLEuVe0my3DEpyYWMJhK1jVKassuxivo4d8JoF8JoPZ4qS6KZrVMva2tzVPudYTs+JYWFpewjS78nM5hWd/fv0rHJYqqLY6CMcTshpttg2TslrD6m2RrboPZnelz+o69vj8+FziCd7PngTMwgzZYefrl05HQjtl1A4G2i943z2xYZ/bIAbLgLN6xX6Gdmh8f67tA2RiEZw/u4J4NILV1XXUSHBRjOysoziXuBZzXtLiiXNX+S2AyHFmiR4eHanDOZ0066eJyQlU62W0OpYDy/W8kC+g2exoXPN6j46O1SlmQcE2TlvNtuo62R9+R1ScqKW/+49/AXfgSpahyydtnOyQTPsZ73dHtpYbJttnbaKanxuBfWd1RODYLYw6aEgF72wcXMAQ/30c+MPWODvI6vWc5ZJN47H6UkoBtyCxsOI1+EWXf8oWR2ynbZRkdllIsj3UNm8DogSgEPRwrb8KC9VL08+O5Id1PlhRYioC8w8mCM/cBGuLo4rQ2qoNfKVlggKS2PrGBYhtyM7n3lte+Q2Id3UMbrsOlnBIpAhVEfps/IzqPHEljW8XJWMeOHCSPLCCzNr5uQnoEEASRO1v9M60azFAhUFcbV0ff065IDwU0AqHtkjaxIww4KGACzw3ES6iLGYU0uPCPr3SWs9ZrXm2+ak9MMJ72DLPx0gI7S6LU95bts3xffvIzxtRwWsXaB6yYPHfJ1HBFnYSFbxGFgtRtYdTCUHFTFafneQFi8hmh56kDBWl96nZAIyemSPvbKyM7Q7436eJihO/ozwWUwEoE4Tt7EGiQjZkHVkwMHivUamgWa1h8+lTdBoVqf1ZFCrMVq2yNl6YtVKl7QCDqZz3ojy1w2GUCBY12B0yoeLJExWlUhl7pbKICoFkApAcyTjKCfDBlicV2h4gC4LH/t+CQI0H7cZL4hD9dkPzIhh6rtdRiO9J+x4/Rl39c0JdGSzWTNA6BnBPg09+rjNQkxs9i5Tp6Vm1j9edqqbdqKHJ/9UqqFcr5jebzcsHtTg3p1Z+1kJHB0eqBSani2jU6ypKbn39FbbW15h8byp6qaQ8AO/Apt8DUeFtQux+BP3wT246r/qeH7P+NdhNwa6KIOg+IipUuNpaeRo81s+r5Zv5jmxPnRCxw7WKhwEC7gweptKZaiOqVqk85WFm7/k6Dg72dNFB1bNdk+UzaIq4Q5u/1uC1Bz9xcPz49me3yDnFjV2/Hwf+swTJg9F7eFuhwBz3sJ8p+k99eZA88Kfe6xRRcfK3mGPiQkAjRg5PThRl/8CA5ibtxQjeUcU6PY16tYz1tTUV2gxJDn69DGj17dD+Z+0Zjslefz/kIU2yQv67UR0WGbY8PTmBKXmpcv9ie3cUiUhEIXFThQnEpehjWz8EVMTzGdx/to2/+emvcEzbtHAPYdr8sO05EJrurycIrAZrDf8cgqSKb533KnHNMN/27fKHNDbUpearBavZCWLZYRtIpob4s//qL3Dp6luIpydwUKpgfes5soWsWtHX1lZ1AGDY7NxEDtWDXWw8fSTFGJV1AhSPjrG9s4+5hWWcOXMOGxsbuP+AAbj2FVzvf9Pn+n0RFR7A9fdMvv+OqGBGBQ+HkTA7TwaYyJN8Mosmkto8LCmU0+WMUWGteoDiENmXRDWPaetIkODe6gZu3H+EcCKFt957B++//x5CkQSeP9+RJ3ohT6IiNSYqagzqJZDBoEAvQjCSgdYwPEi1ahX8/B/+Hs1KGelYBDmSFPQzTsctwDESwf4h7/uungMVZKGoWQ9wvnSoQNe0sLU2aP30uxAV3wL7A3vKaaLiNOnnn//vQlQYMDDOJRut2y8hKvyctfd6NVHhgzb5k/5QbfOwL4ENx8i48zImIJxAQSiaGNk38P18RwXrGp9Rwev0xBrHiScqgnuE/xlPVPiOCl6PB5OMqLD1TB0HAj18F4XPhrP3Ul3piGj+ndderR2fICqkIg0QFax1pvoMlmZIb1ldzXyNRNzAfHYMsK4uHZWRUGYCbVsiIutYHwmgFbljFiwC0Hnb+x38u3/7bwQBfnPjBmZmF/H02QYqNWZTZNFqVBSU/MEHb6v7gnYvyUxKPttcnQjM0OaV9U2tWgc1yVRbM9vg5td3QQGrrHcZbu8UrFoD+0Pz5M/l1GHEMHkOH3ZUvP3ma/jss1/K/oZA6fT0DDa3djVnzp+/KHCZBUwhnxY4ubg4L4CbgNzm5nNkMnlsbOxYvgKtADFEKpNCs1VXJposR5OszQe4fPUK8tk07t25i431DZ37Ll6+qGwM7lcEpHef71mHSqWGequDWqOFeDIjaxrlc7DmlDeTKWQJVHNNYA3OayXwzg4IKV+daIxrAXNtRFQo98TOYroHFEN5P3EBfQmz1uFrk7BKJjVjNIdoceLEcOzwlCJYY8/AS5Kt8qrvMEuPVj0kKwjamqqY9+7KlcsqU0RYlI41T2jR8bOf/TMeP3mmrCnu1xTlcUvimONYYld9XLmDURTScUykY5hg+Gw6jUePHgnkC8WT6lhDLKFnfPHiJRwcHKDd6simh2A2z7c8k3PM83PPLyzo2n2NlMvn1FFBoolAndmEWFCwcgwFPo7t2sx2zSvjKQ50ALybAzbHrbODZ4xejyprnheBtjqUwug1GriwUsT33n8H2XQCRzs7GEh1EUN+ehYHe/u4dfuuvNUvXbiMg1IZh+UyqMKenplDrdYSSXLh/AXcv/9Az4EPjfZnU7PT2NzawoVLl/BslRkVF1BxuSvdbhPXXruMTz75EPXqsYQ3ujftrs7wJCDj8ZSyOv7+J/+Ag1JNexEzp2gdqHB2hgJLGkeCoAAAIABJREFUXU8bJRK1tH2ysx/P+v6crmcaM8tl3j/+PJ8BnwnXJZ9JaedYIxx8RwU7HiT2IdBJfIBKZwKevm5wBAM7YJQJyfrFkW/WlcBOCiOc+V4e5LZuC5In7VHt7OshV5UYoZZM4uKZZTQrx4gMewj1+7IZZqAxc8WoXr/z4KE6nkTStXsmLnBzkFhLuUarLfvc/CKZw3VMuZkSuZh1FvcYYR3ChQzsl9BEmZ+G14zuTc+AYs7PTrOBD9+8iGtn5tEtH8sG8t7TTdzb2EdmdhGRVE6kq+yZYiFEE8RpuurgpNCH94xB9xzPIkOdcNELZXmPlpYXJZI0YjuCVsPyN0QeUMme4rnfhKfeVkf5oMQneL4mkdlgkLfZYtFe1KRb3MeM4CcwTlKV5x3t88IJrOOFz0vkRzis8c49R92A6jTznZl8nbE12Kg2Ue6bE+647gLRXATN3RhkzStLRGWCjQVLvC6zLjOQXkSIE/Hw+nw4u+xeBcITj7OaikNTr8fXJhHs8CMR+SRw3HhgV4judb+LDm0PdbCnbXJX4P3K3DQKmSzmpnKySmJnYIfWi5WmbOzYiRZLJjA9Nye7z0qjiTozeljDu44Ka7ke45PjFDhb1yWWdnihanDXsU0RqBEVNit47epkcjlyvMfE8VRd8fNyjeA6KUGv/budNT12aJ17RkwOZGHK/7FrKZtK45tbdyQA47V3SWSwlghBJC/v93Hp2M5ezBmNmCU3X7tSrmjd8mLgmdkZdY41O8QkcuqW5H7HxZHjiGOU9YoFtbOTkJ+L+CP3LSPbvyMqRke07/7yL+UOTHUJkrtNSGmaBljLBihOGyBjVn1LuTw+eyxwfbhOTwsvJ5OAWxV4tmGb+tWsH8i4SoGvvAcqoGKyIFCR7kJTteQ4htTUhR6gc6yqFPxUD5qokYsN30t+iANaMXVVBHLD5ES2ELWu+dE5IIzXyc4FFXRS/w+l4CFzad0VPDCY/yHVTCwwRBxgYDYE/Fxcj7loUcGTTKnoZjF67tw5RONR+c4dHh6pUA+C2/5gO1JLKB/C/Oz4RYsfhTTxfUae5w4gV2C4qT1ZtEiB1Gq4e8ngZNsACcRb2I61hfI5ema52bb2VD4/3g89M/2OMfoEMklaWKhSHyyAWfxS3eTBDMvZ6Gij9T/H58YCTxuwNhjaDVgHBUkKDqpu3wK1ERpgYmFqpCRg+x6Ly983UcGDD4kKfnHBj9A/UuMwhlQqa4enaMxYaGUTWPg0n5d5KRuAekId7eaBH5c60DtQ1B/W/QY3AtSdNyzHlicq+DNdtkHzMKzA9S5q5bLAwU6jgQFtiKTICot0M19QvbJavfk1kc/rGtX1hJAO1sfVin5mcrKgz8WCgtdfKpdxVG2o6DTyzfwZvcrK2428DPQO/vvpz+sBBa9qH4OpQwW4ybPUFVV+zVRhpAJkXAwEo3h9gJx/39FrjsDjFxAVI1mpeZPy8MswbT7TlZWzIoQa/a6K3lqlhHajjm6robA2Hs7TmSJCsSjmlhaUZ8K28Z3nZrE1OTWpg9K1yxdx7/YtERXsyPD5I754FPCuU4PvqPBHiG+r3vXZf8uOCvvtAIEU/OsrSAy9u6vUBP6QqHChgR4MGgFDUrCfvK8nAWaTGpPYm52bkZqUFgnl8rGK91iMoXIEx8NIZ7KYKFjIZ/loF9vPN0eFX3A+sWj3BFVwjLxoHAbHnZT2Wl3dfXV3Z2T/FFAu+89wklRzd9TNcT/XTxMBL+oM8D8zAi9lNWc5FcHvjesDdt1Y67wdaCMizt55513ZDjx+tu6Cs0Mi10tHB9jZ3rY5cyqj4sVEhQEOwY7xb3dUiDWVfSHVTtOTeWQzaXUnTDAUOZXEZKGg/XIwYFhhB6mE5SeRrNAexfbl4xp6ww7SxUk83tjF3/3TFzhuNjAM9xEhSeWICre4jDoPXkVU+Ps0+hnn8euJCmomPFGhPdwNUf7Rcx2JngzW4ZFjiiVBvI+//Lf/Hu988AMQByKQ9+TZKmZmprC0UJDCeGFuHjtbW5hMpzA7mcPdb27im5s3TJ1NP+RhCM+3d9DsDOThTFDBe816AUSwEy34fDxxMfq3QEaFH9/j9c0dfp0Q4FUdFb7TaQwU06aHNRp9gSNYWZhDPEqNIYmKHCYmCrKW5Gd6cO+eagsRF5m0aiQPTpOopwjj4aOHWFhcQT8Uwa/vPsSTzW1MzM7jBz/6IyyvrKDd7qujgnvqRL6grkTfUUHrJxFgJCpcR4UA2kYd5XJFB3/aGjJMe2djHZl4RKGL9HFPp2zNZv1C5e36xqbmuFriWTsKSO+i0eIabh2jJmgxMNLvvyfWiVd0VPj796095gUdFcFaP0ha/DZEBX/efo5rliPWXM2rtfAlREVwr+T+zLH4rbniLNCC3ReeqOBrsw4zv3PzZOb6w7qAh10SFbKAc6QBr1MiHQeSnSYqeJ/4PQ/OBevaIFFhwIf/X+gEUWF1ru+oIGhn67/PqPCv4/cm/yz5mWp1AlYN553NvJJxR4VfW/OtnIQvx0fH6pSdKhbRVncxjECLM4yZ66rZX3JOE4yl4vTo+AjPnq1qLVcHLj3puR52W/gP/+Hfo1ot49bNm5ieZtDvc7SaXSSlyOaZI46PP3oP0UELPXb4qBva6nWO0Wq5pkwFdvKSHDre3VV+xcP7a3jy7DkWlxfQ6Xexf3iAK1euqrstHo3j+pdfIZvPyxrj/sNHulc83/zxD7+Hf/z7n2BlaV6+1FSG7x+WpGC/cvUqdrd31E2xuDCj9TKXTSufIZ+nnzptlVJ4/HhNNmqTxSmJkVJZdjc0JUigbdHFC+eV8bO2tokPP3gbZ8+tCPT+9Fe/kr1EcXpSY/rihQsKKadCfmNrG/cePgGz0piHxjBe/gwBFp4LCODLjpP2Fcclnav4miIoHYjj54rPJWSA9NB5TmouOYETO8VZ35oFiNmIsjbh+swzSzqZEjkjtXu362xQrLZnvW2kiREjVEN70Rw7DZkfNz8zjVg0LCL7448/xJXLl3VfLOibuTlh3PzmDo6Oj1XvKKCd5JiCaoeq7+UkQJ/3WgXpZBJvXzkr4ou2WY1aFXsHR5icnsX24TGGkYSs7Xho45nMhG9hZHJ5BXzzPhBc5f30Qc/emoXzm0BVrV4bndusu9EU1/ycXN/92UZdlX0TALCbUvY1IcgamK+9t3cw6pBkndBq1JDOJBRYbYBzC+F+C7lUCO+/dQ3DbgtPHzyWpW4yW0AuP4F79+/j0eNVETNXLl/D6sYWWoOBCIvCRBGl44rImDdefwPr6+vCGmifQytR1pYHR8eyZXv89BkuX7mKSo2Coobm4xuvX8Ef/fEPUD86wJAgdKuj0Fl2aNCekv9jDgs7Kp6ubbs8EqiDyrsqqIMwkVTnCe8DQVdbfyyjiSQ5z/o8v5IEYW3D+2gd2gZIq5tHYs2+cAJbZ5Juv7JuCSqo+WwMHPYBwfZM+Hs8I+vnnLNFULDlw+b5uhJ9OjcGW4t5rrYzlFkK2sKrTg/Z7Qwxnc+hXW/inTevYHtjExVmnLDzJJVAoTiJJ2ubSLAOKBTQbFu3HDEU666MKeSd9jvK9XBuFZyXFD3w2pWPSOV7o6E9haA2MR1ZQSvHs4t21wSd/B5rjn6vrfOq8jAjwLvXzmExl8GgVsXrV67gZ59ex+pBBemZOfRCSZTLDLLuIZFi/wX3MiASorWS2dwoOFtkAjvcaJld0/zmPaKgita+Ihl6Pa2dnMPchyQwdTU5O0qIvZB4ffrsCWp1s4Hj+s7nScKU1pUUvlEoaI30Buob+M1uRMso9SJbit+8G4fWP3UC2vrDseBdIfTMXCfwaH93kv7RacytKRIJO4yKIh3tk47o4v5uRITdW2WGOjKf/yb8xp13VJO6LmdfF1hHhe2VvouZFmn+GcsynQHaTrCqdZ3OJsJRrAsvmTaRcCKaQJcdRByjtF+n6CmfRDYdVdc4u8Fi0TjYuXtwVFbnzbONbVQ4h4g9MsdGfDk7q20ejeoh3nlvI+sJF5fT4R0aeE9EvLhOIL4On2fQJUDfc5m66giRC4phk7JH5hwS+RiVLbvWTp1vrWuFQdrxEHD5wnlEQ2E8evwE1JzFU2lZpg1CQ+FkzJhlB83h0aG50zixLK1/iTlRjEDskYQGhQ9cf1iL0JKMNYwEFLG41hxmXPFniAGx/lZwvMSCCWGYXOOJ/X1HVAQr9u/+/i/iDky2WPxbQa0ihCF6VJX3qMxgIKIpmC282VQrVKgze4GbPCcYNziBtq5DgQumVxbwYKQN2SkePThnHRrWyutJBwNb+P9ci6TWUyuovHJfaiPX0WHoLQmVuB0Ch+Yzy6AsblKFXF7XzE1JSskEfZCTFswof/qmCmxO9FwuI+CYf5c9TNfaB1lkiKhwu4bsr3gw1oeFQJ35+TnML8yLRCFTzN+lryI3B26iPLRby6gx+97HWy35tJIS4zsQOM1Chc9DHR0iGmwRZfHLTgce5Lkp8Jr4A5a3YUUUiwzfCWPBTq6zgiHMoZAKQQvcsUJYBEW7owWOz5Utflwc+bz5uUkuUXlCMoabnt8gLIjVVER8Xd4PLpDcPLnxsW2NBRhV11Qz0H6A7bb8O1V+hcWiro1Fzkjdr3Y5EiQs6k6CfrwXvk1SxYGzfjoBJPJeubHCXAgWCq1qQ5+LgAxbCfmmXPRTabaDEtCK6uDOQy/HkFcKeOLIAFF36HagiP+eDkcB+5nRIdutCmMgyQWD0yMxnVLAsIpcZ7fBwzcDEjlG4yw21KFifro8ZKo1u93RwYfPrVk35QbbpL3ahv9erVRk/cRiZmIiN+qm4L2j7UarwxZ6T/75DgC36dN73sqckRL9VYubB3c84ebHXxBcEUDSsZCtk6CL/deIV3CohgeLbTCPvbzNe36clSDg0mE2NgeDIO1A+a2a5wwcVJh2WtYKHD/NTg21allrAduHB72u8hM0nghYRNmSek6Kx3aHeR+rutc6OO3v4+rlS1hfX8Pu8y0cHey7AtOKPrsnzvZmaG32tkhY9o1X4Xgl8Mvu7wg4O9HYEtSRhDA4mUE9UrwEiYYX3fN+p2sE66msiHGBPL4qU+Tbf2uVtVAD5CcLWDl3TgXTxtq67gtVNNwrrDWZeUYTymHgb7aaVayvPtG94dz3uQj2vAkUuEObywiyx+/GZ8D6KDg+eEdVwPLnXKBgsPtBeT/BotypeIPg5OgzB6yfvm3xMn5V4xtdBoULWxzdINd+Yeu1I3xMCKT/UZnKNdNsE6MC0N56+y3dq5v3HlsrOIEsWXzsyxdb958dFQGiKThmXkRajMkeH+JtAHh4mNDBNZUM4cr5JQNh4iThzeaBHtqT+ZwIbSrruOYM+j0B0bT7IIBNQIm5AeHIEOlCHs/3q/jJz7/AHpW+Me7RMr090WXgRs7YhkrT2g/sALMYJNTcOuuJXu9Nq9vv7Bb1HJxv7eiZeGspMYCczmF88NEn+Iu/+m9QqTVx4/ZtlCplnL94Du+8+7qCIhWcO+ijvL+N2Zl5HJYa+Lu/+b9QP9pHiqG4DtDZOSwp2LHV60v5Sz9j2XLpOkJaV42w8AoKm+86b/rVLsS9z/7LFOr+Pqgfx/2+D9O2+6Qxf2IdsBEwGqcD+zvnFQ/ztBpZmC7qWYb6XUxN5kU2eQuLL7/4Qs+TpNRk3sgLdo1weZ0oFrUO3rv/AMtnz4io+PzmbeyWa7j25rt494MPkUwxZLUn60H6y9NGRsG92mPKqFSP5XfMGoo1AwFgfjaCB+WKs4WKxaX+vXfrtuUx9XtIRIbIMUybllGxhH6H/sXNXkd7Jg/CvBEEfejz3+pQHMP6yAJJHYfv7pnZXOrA7hR2WsNOkbvB+XN6LgU7Kr5FPhorFljTfWj16XE93uesSh2zqSOiyl2Y/ltr8kvICBdK/rI9w897r+r1JJnqZNVcJAfCBqLRBiEawfIK7Yay7ntjGx1vfRnqmzjJEy2+k1nhx7J+tRr/9JhWbTgiK0wJTJKfBJmsGZxS2Idpa6Sry2vcVREk+VRfRsKo1cuyX/SCCK/S9V2jHLuzoRl89MHHsozIZWh/mRMIbV20FMMQNG+jUqkhk7L6aX19U0A5x/OGOtm6muP5ibw6Xp88uoc//ZMfIpmM4dbNb7C4dAZPnm6gXm9pDKbTMeSyCYH5vUYVjWYduWJBFhAkootz80iEY+qWpU3S5NQMYuxa7nRw//4a7tx5hNwEyYi0FMyXLl1Eq97UPs2O6FK5gmaXJAYB8ZTgsbPLi3i+uaYQ+nwhL5CiVKmLSJ2amRUo3mzU0WnVUStVcOXqJWSzaXU6b25uo5CfxObmDnb2DjE1NYPD0jFm5qZFbCl/i919xSKuXr2MSrkksJZdfu+88zaWz53Fza++wpOnT80vnFZZ2QnMzc+jOD0nr/FSuYa6LLUGuq98hlxreQ4UGTYcqruEZ0cBYP2+Mhj8GYZzgWcLs9EJoU4ynCCyC7Tl2thqMODa6gCuNxSLca9gXcIzXq1KpWpb894EWS5A1c0yCdZkJ+UU3/Su73fBpYb18jtvXkU2lVLHLclenif52nxvdXrl8vj5Lz/FgwePTI3Lc14qpTqInQwkSrhfMfuA9jjMdEiE+5jMZXTWXF99po6WAaI4rjXVtUaAi+I4gp48R5EEbtB2hYJBl+vI8UvCiZ+n3qjr5zgXZNvU7ytUldcqosPZgpC48WuL8lDc3OU6x/nIe0Uff4KwPNvz7Ecyi/UVrbB63SYWFy08fXdnR3/fePYQw24NH733Jooz0+jXGzjmPtnuay8JRWMKDKc48ZPvfR+/+vxzDNhZwCwGhJWzwY7lxYVlbG09F1lCUJxZJIVCXmfVmbkFPFtdxYWLl3FwsI9+r4Nup4E33riK7//wEzRLh9qLeW41MsAyuLo9Cmoy+Lsf/xR7+4c649F+ULZTAtFJDDBr0oN9xDzMp57rF+8/9x0GRZPg67m8Fdp1+c407eMKtzZwmusGMQV1BhNHGdKCxsKVe12zsuTn8y4QBn4a8GkgtpqgRt38AlYJirJed12qAl/VMcqzsp2l1c1NsaYWXVej9nsK037/rddxtLsre8viRF5dFhQAbDPQuFqnqgNtdkB0+1hZWRL4T+smjgmKkDg+OxQsOnEk6wV/D9StlkiotiDAy3XZgugtA5SkEckjHzaey2fV6VavV5GVzTIb0Jp4/43zOD8zherODq5evICf/uo6titNpKfnEE7mUTqqiTjsdBsIxUkO9RXaTYKV6w+vl/eN4+ztt9/WnGD9yrnNscruNtrk8DNxD6qUjqVSl2vCkDWxzd2VpUUsLy0J03rw4IEIDtos5wsTuhfsPGF+AwkRWUKR7KbdG/NPlMvJ9ciF43F+aW/g+ZNkS2UkyGIHmQkrjAi32mXcMe/3R40b2XsZ3kHwXBbs7KxwVt4KaZftloU9cxCZZsoEw96yin+X20ngfXylYR06djbj3/V51G3W1trO32E3K794PiBJxeulCwhdC/i5qf5X5xcturgedXpYWpjHyvwsioU02o0ydjY30GAXVZOC4gGSqahEQ8w2iiXTuP3gITa395Uhh3BU+6dEHCIOzYJJc84VQXY+MNGBWTSJSbSuTVfsWX6FkQwcuyKp3WfydQQ/ozBE1y2l++7CtnmfJXySXbqvh3T6FBkYHfbxxtWriEViePDgIdq9oYK028RQh1xngbm5OYlIiQvqdUR+WrcN9wnWxvxsPAOSGJmfm0OpUhImxbFDnFWWj2GbX/w3dj2LGHT4m5+XfD3WSN8RFS+rlL/79z/YO1Bs1UeHX6oKPDBCpthCs0OaKGYX4A5ojqHlRiUgUgWWWUpwdnKx5QbOjco8Ru33fPsuv8/Jap7SI+GlW7Bd4JdXtHsg04HushniosQNntdLv/Khta0ZR0qQIoKYsg8MTJDliQfJqMhJ0PKHCpFJU/ikUtpM2AXhPSi5LrItS8C0OkOcgs91P0gVIK86Y+65YXOT5EakIFQHTHEB1zWx2AjYBflQQC6iApxd4BwLEU8+8Bkoz8C39rFDhKwvFTKptFQVbDX3B1V1e8jKx77IiHuQn8+QXSdBcFv2AH0rlPwCTrCei6ZfvPmZqHTkWGAhY36mRjLI17PT1b3koY6boaCbkNlMEbjhnzwse6KCBVZhcVIbCK/JAExTKHiFSVC16JV7wUPxbyYq4IgKKwqMqLC2PxIVvHfGlEdVbLFA9zYCXs0nOEJ2DWN1IP/thN3TKX+YIPMvEIsqGA9VhUJSlFDZz89JNYKUXp2ubIV4OJa1GtsKYzYHFF02hL5/tM92cAZUme+yqaqsA4RhVgpxd50LPAh5KyuqOVj0s4hnAeAB3xN/CgjxPqRmzfCqryBR4Z/VafCbRTuVVp6oOEFEuBc/cQ2jtYDAnyMrCDC7riSPWQsPdVUWiRyNfa+y5l8iPJgmdX9SyYyUaJznDMzsdGsYcJxq7bGigYQWAeIOOObjmJ1ZRDpbECB3eHwo0pBACQ9KF86fxfPnz9FpNeXPrEOJs/6xenNMVNg94j96+x4HvuteBxe9k3c6WEwGv+PvlaBQFjwvAfFPP7fgfT9NVLzqGZ8G7fl+LMJmWYCeP6/7t/pkDUcHB4hFTJ1oxGsCk5NT5pmqgreB1WdPbBJJ5WI0rZSTnPXKTWDBfQr801YyJgpOEhWmXOS/cdUXhxLsrnBB7cHP56/v9DgMgpTfJirGrxAkHr817vw6EMiGGIGRVNiGGUTOz8quObMbeeP11wSIPN46sO7FaAyZVAr7e3vY39tXTo8zSBtdRPDaT4OrJ0gYEo/ccxlyTXXhIIF4KIRCNoz33ryMhbkZrYP0bWagZToexUQuqy6Lbof7jZEVPMjNzc7JS3Vjk10xYaTSMaSyGRxVevjxzz7D6v6uiIpRCPSJuW0QbXA9H4OxQWppfJ89ic9/Ofl7Y4D+JAlsyqvT8yYZi2L57Hn89//D/yiv+NX1ddRaTZy7eE4dUhyP3VYbrfI+qvs7yBWm0AllcOOr67h9/XNESK43mupcy05OYWv/AM/3DiViGBDQcs+HHu8kKgi+jDJFFIzsj4KWY4GQ2S3yy4iKQD4NzALz5GewQ1rwztjfA/dTZZBZ3AzQRWjYx9yU2XXx+FycsBwJAoI8gN++fVtjb25mGhPsqAmHFdhLW4zZuTmBp6urq1haWUG928XnN28hlMzho+//CAtL5xByitDt7R3kCzkBPepKHXiioiRve62/CVoqsG6kj3ENlQqDjCkMSOve1GsNNKplHO/tYHtzDeFeAwnmBmgeZLB/cIBStaIg3UQqpr2Nv0c+k9aHDdllmmL79Dx3N1P7RKAR4cQ9Pj3vg3PrNFFxcq7xWY42HAMcHOlqdIQj1V+wuHrF38ln7Z6zR/fd7518z5PWT6dfWj8rHtnGle/0MDsJ645lvRlTDpMRzgwLZpAqn523YmINaPabtBOjMMkEI54A4fc9UcH389aw43rAPosvQfnvfD0qwU1depKosM5DA238dQfngK9reZaoNyrW3TvqemXeGm1fzV6Dn++Tix9jujhtSnsFrVYlRiJBQ/FGOEIRCJWTliNF4Il+5LLodGHgVLvrntBOFgTGasp8IVFx78495CeKePxkA40G8/okycJkIYMP3nsT4WFXRB1PPaEkMzIilrPQB9L8/BITmc0tn8OtW4/QaBLm6iOZSatOI7AhkiIaw+3b9zE7T4vAhgBGKsIT0QjefectXP/sU8zNFDE1NSWgbWvnAEelEi5duYJ7t+8IgLtwdkVAO32y+UxogUUv68EgjAcPn/CEoG5mfk6SJSQTuwpLjWK6mNeOeuXKJeQnJ/DX/8f/KZBxbmEWb771ljI19nb31L3SrLUEoDXbBDaBSp2WHgSxTEku2xUXaKrOIhFzrGHt/Mj9xtuDcg3i2kFwjOdNhdayTnDnS52FRCDbuYU/x/HL8F5+z0hKcwXwoJ9CbtsdhZISvDNyy0RYJBbUxU//fQatRkmStHHh3Bl1FVLFz44UqsYJ1PFz8/ryk0Vc//VXIlQ5filyI3DJL+VL8ZzJ882QoFwC2UQcF5dncXSwh4lCVqh0uVrHuUtXcOP2PamI6xQs9foo5HI4OjoUkDw/v4DJ4iS+vnELy0sLUtOyXmW9r45UDCUU5Lni6Kik+UmRjlcU8/jpbVA4xvnlz09cL6JqP+TRwERLXGdJdnB+8N7wrEEhQ7vdQDLBHIk8omECo8Dli8uYzGfx6P59HB9UVT9ce/0NkUZPHz/B46cbskW7cu013L3/CHVmuPT7SGdyaDbacmu4duUanj5b1X1lHgXnKgWGOzu7WFxa1v5E6ycqj2PRENqtOt566yo++f5HaJQOFc7MM6jOVC2uXVSZU+wXx9/++KeolGtIpjMC8kUm8IwagnIJSQTy2ZNUVw6lMgQI8FoXOM/hnEeqUR0hwDODumdcd4MXG5Iw4pcCkyVe6KPZ5DOiOCWu8Gt1nEqEaLZQBoSaKl72x1G6FdA+qe/IKVO5m02eZUN6QSlfjMSiOtKIiXh7HK5dGGIilxEpFuGbDoaolY6RSsSwsLgkYunZ+gbWtrZlz8Rsj0qtpnnPecpnLHIxHtf9V70FkoA5jT/OH/6byD8SP8qGYe3YEWnEzl1a97DDSPu2E5lw/IXDQxG1Ilq6XXz09iUs5LOId3uYn57CP332JXaqTSSK8wjFcyIquHb1+m1EEubt36BtnwD0nt6DuITISOIxAt1JzNNysqb9QXmfCrdi95UJXvb2D9RdnM9nJSSleIPkBhXsrJWU3RSLolSuCi8i8UKSj2s0zzbszOMzl+qdnfrt5lio45wOuEZxjeM4sD15IMEPHTv4Wl5QMSIrAqHR1o1j+Jnmq872lqHK+2gdFa4rgPZ3JLvULW/qGJYTlt/DsWPnJQlNfcHk/pQ1VMSLRA33scwnc2Nf7BOfAAAgAElEQVQgpiOQX8HuzHIheULshuJZVaOyvmJ2g3Ar1g09ZhF1kI1HUSxkMD8zhUSEYra49tpGvYVmo4tKlVlpdSQyWZRqJDy6aCvjMCKiokOs65QNpOPirDb+f9h789+4ryzL88YeQUZw3ylqpSTLtuR9qezsqurqwaB7lpppoHswmPlp/sMGBhjUTC1dlZWZdqV3W5KtjRJJcd+XiGDsg8+57wWDNO3KzsxudBXMhNMWFQzG9/t9y33nnHtOjzBKz1YdQJ4bGXG1WAsxN3kevv55zSaSJ+BzInyDtXzM+eA1jmlCVHiODTgi62WGD9Ls2Buv3tTa8N2jJ1rD2/I89zB1njckGVZlIioC6QQ2IUyVPLaNTe3f3GM+K3lRm5sb6grndbKoS1P/OpbJWsD4JysJcStjlGfIuGJ+UiP9RFRcUHz/9K1/2ndglNY4MbUeUOZeiX7YqVU9tJpJz0LtQcwArkXPoAhtWRxCtLmT7RA2C6kWmvgseo6BAOCoeGch71lAvZ3KNzSdo+SJHTspQihoTyvraUZG9CN3MkQ2UGJPM1q0dQALjCwLKmw/isJLly/bzOysitf79x/IF5OFgEWC34tylH8DYtIGTosaoLbUX4FZla1OUArBmKpNnLC4Rl0euPI5lJqWTfk0LJP70rXFikpcQqvwi+3JnFDLbvTcC4oNCoAIpqG8ib7XWpxD90kkGrqdGvJDZNPxhTkuxuqaCWQRSgMV+SE4SGHc3RZDVyLRUSGvvFC0qFVaCpgjsexcO+wv95siGeJCKp2QUQFRQZA2BcrQGaIi5pQ4CYCK+HchKqK6SjZJbe9EODm6mKjAQ19jQy11TlT0+oHGeyySJNqSBeIstg/qQB3bbMIScB7s0M+fIyoG8SzkMBBCpsE8UJpw2OCzEFSvMHI2/bZZPpPVIWltZdUagId8E9A4oAGRyHHFJvPB52880PNtkVcUSuEaznxOviev6KgKdp/o3q/zAGkvUSHorMf+Kj47xgDWT9FblZ85D66eBxf15wjCB/VHtHr5IaLClTHh01JTqA01p04KFHD49XK/ab3s7yOUnALaA7NUvDSbNjI0bFWsydrYE/TjG+PBdwlvt2ZtOzo6FFFByB82OPt7OyoOyKlQA0gAq3SNXQCml6gIauk/AFEhxDtgmE4MXiC7vmBMRqIiPovzz7n3mZ8H7fnY+IlOX7pkkzOzepbLiy9tf2dXB9cIoPYXB0QOCcDj0F6r2NKLBQe/sMP4gxAV/vicqPBsgi52yPd7iAoN7zAn4rrbe51/CKKC94v3K97b+EyYVsoMAAhTDZ6wV1+5IxsFHuL9p8t+sGX/KZVsc2PDdnd2A7jtGUvx63cnKrKGg+3IUNY+eOc1HQhRhGI18c03921idMSmRocFPNca7dCBWFNH1/DIiM3NzEplhlpxaKSolvjjWkJExXfLS2bZ0FHRowg//1nPz/0fqpp+jKg4vy+cEhYudujRo1uy0xLA87//n/+HzV65YimIs2TK+gfwy6UNvGOdVsMONpasfrhr/YPDVkv028Lzl/b5J7+x3bUVS0Ikn1Tt0uU5S2aytry+betbAHOH1mnXLc36EIkKqTlPAew/PFGhBV63LeaPcGZSQDahjBAV1rbZ8TEdwHPJhA0PFqW+HRkeVSfY5uamAlYnJ8ZtoJ+28rq9JLdjYMhGx8dte2tbns+z167Y9sGRff7gW7v+yl279877ls4ULZXM2kmjKrKWtZX3BrSLRMXR8b7lcgTxhjBtxCKQEpWKLOIE8hX6VEPWa01rNU8sn05a5XDPFp99a1tra5buJGy4NGDNel3dRdglpnKejZYvFGUx93J1zQ4Oj3v0dWdHk3ezuSVGL1Fxfp/yvdEP6Wf2uxCmHfe2s3//uxMVMQPolMR08YsO3eeIinNXdOZaz8+l+Gethz1B7d6FCiiGzWlWOQjq3Egm7PLlyyIq4oGeesFVwU5UYP3U26kRD/ZdoiKseQLculZW3k3heiUfq7yXgkbpzg5j14mRi8O0e2uCeF0AzbV6WZ0Z8TyibmUpmrNdW6s/ef1nRrthf6FP44y5QV2FerrZRu3cVHh8p+UgB+Q4Y/Vgf797H6gPRsbGdOAXCJM1dSb05bOykUqn8/bFl+Q1rFqpVDTrNK3Un7EP33/LTo4P5HneSSetjlo6kbDi4JDVyiciRbFIJHCaewLA/stffGI7e2UbGB5QDbq1s6NOOzqLEFc9e7ZoeFbvHRzYIV0WHbfRuD1/w54/fWyl/oLU+RCN23uHtrN3YHdevSMRBQQrNiu1SsXGRkdseGRQ3aOAZB2IikfPLJHCCiyvs0+ZfArsbXNZq5arNj09buurqxo/d27fsomJMRGdi4vLNjJKRhUWkJN248YNWbxsrG0KjF7f3rdcAeCzoiw4t0Rq+ZlMtRJhox09H75QwqtWRO2ufD0XFkXhVKwJAeY4Z/Dz6hZvu/DNz5Xk3XlQstS+9ZqejersSlmf1fMtHDjlBwQoh7oVIpVny3iChIZZoluF/RrgFoDt7t3XbXJiQuccQHTOXw8efiebX87DnGddIAMhhwqfPAkI/6osoJKtps1NjtrM1Kg6XshIKldOrGlJO6rWrdpoWzqb1+SRLQ2gNWdIrHabDQ+a3gt+/PKSD/OrTWdAUfYhlQpd8nnt44DeEewMec9d+6BYqyGEY5zV6ifWX/JMu+3tHdVuEGrqgiL8uHKk8UAIONZ9rQYdB1nLpNp29eoV++yTr+3Rw0fWaiXt1TvzdvnyrA0PDdjz5wsiC195/TX77smCHVTLOksPDI9a5bhi2HddmrlkT548tbGJcYkJ6LRAZEin3507r9qDb7+1m7duKh+qry9rteqxvf3m6/bOB29b5WBXXdF0m2PPJH11ks4YwNM++4//8f8W0Ez9R06E2zpD4UNUeLg241OETQAO3Q+exwDJWnehYCChWGuifU5c3zj7SyhA0G7IlGBcIh2IodrMewmjZHkUcu3c+8AFitSrxnnfLQ4lOIz4iNZXz+ykRoxjlp8mC4hxoH2u5+8zyYQV8zkbHRqQWOzWjetaN+jiISuqSX4B5MVJXeIj6jm6P3gvSLaDw0PvVM5kBcwLbAWXJd/DTErw2BUqAWTIJuVzA9ryGmzE6H7QvQydJ8r3aNY9VJvvd5r27uvzdnVizDrlqo0ND9vf/Opj2ziuWmli1tqWs4N9HC/IwTuxWptcFgfcZWHdwCYbFTmhyw5AqyuLz4kwVeJQv0fUSMopkPVxQnUO3U4QUZDD5LXR/YUzAfvGwcG+XBbI3wP7grRhrZLTBIJNqdnJn/GMH88xjWQfhAn3paF7RR4SZICcD47Kvl+GGkXrm0q7015jAHXlZoT1SmB56KSga07zOthBR+sxYXN0mUbBC0RFDOgOHciRqNAZReHUnhPKuPbt2s+7LlR1PYZne3inhXfNu327B3eDC5ILAwGXlOVZOpmWaAzpLRTzQF/Wtjd2baiUlcUsgi3IoZHRMY25ZrNj5VrDHj5+aruHR+qokPBHGKDXuk7ORaEfn9HFOeqnD3l8slYLYuCYERJrIQ83dwE1X1Gs6+cH78YQKUOnQ4auIre27/1H5GLolEilE5ZRfpXZvVdv6V48ffpc2S91thc+P51++ayNjgzbyXFF4w2xMgJtLomxxr5CHhG1EEQFX2CQ+wd7IXDdxxC1NsIevnhejHcs4MEfIGT5Ym7xPYQRPxEVZ6vnn/70z+AOjJYPVKyqcYEwaYHUHiTEhGLww7AT4EWAEUXAgwffarEXsJrL2drqqsBUhX2FDoEIgifSTFrfJLwgcFW3AEaAfthHsYKurPW2X/87FicmMRuQsg/iQqOQYVrWvFj1w1hDSjyKOin7Q7sXgDULAq1SkBQoydhkfv3xP9jjR48tnc3YW2+9rWDNb775RoWnfPxZdGqEisFiozjx0GppqNiACrCiHpQEa67CkJwIWsfrbosVOyhko5XP6T6y+LGYKABcllYdFYQiDhTe5QU9LGu8Xi/0aV8vqPUSUoNCO4aBeXEDSeJBYPxZAWBSnLdUPPOe9QYBXKZ7EQ+RvIb7qzbpjmnz0OE1sNO09vFZ4oblhQlFIcRyUq2QtKSro6LVVEHAvqo26nRSlhDYUoCVnycqPEfDiYro34jq7vchKlQwBl/c2g8RFbmCWyAor6LvDFERgX8/VEOAeVEVC9NIVKjQOjf/f4yooMDoLxW7ZBgKLDYaOlq8RdwPOVg7ERzJXOo0W/IXZ1ysLC1LrcI47/3q+lJqQz/1/I/ggT67CqOEbJEiENALbuAV7T97caB2L6AdwYsIisTPEn+2O2bxbS0fhmwTLzIuAit7P0+XqAg3VmtAOJDJaYVxElSyKvBjq/QpPmipTFJjmDmFwoDCUm25Cl1MCKRUQHmw7uJ6xsfGbedw1zJZCnCKsZSKJXVhaX1pS1l36dKMLb54IYCPPwOcdKTUiYpuJ3UvJir+cB0VAE29ANxvTVQ0mhpTcWz/OFERguCdgsAYVl7Zl69escHRMa03y4vLCk3MgjmpUExbaWBQ9gF8QN7/pFa1l0svdNiTyY0A5dOOCop99z32A4XIYFlC/VhHRQhiZ9QGVdEPExWn8/f7RMXZbAd1DF4s9O+uSVzn+Y6KeD9jwXtmTgi4czKL/aqvkLP/5c//3JYXX9jYxKR993zVNtY3tYegosVOS+3hwtKCQiq84e9DVND0MDqStw/fed0mRkYEmAH2/vJXv7ZXbtywyfFhHdzSuT4pZbEAISwZFerlS5ekcN/e2LHxqWHLsWa2s/affv25ffHdd9ZMehhz74ronzV2VJzaiP1jJdOPERXdNTmoweJB5sJ1pX1ixYGivfLaHXv/jz6067duWUfq4ZT1kY91cGRrq8s2Xsxa62RfgbXt7JCdWJ+9XN203bVVW32+YPXqsU1PjtnI6KjNXL5hv/zoU1t48sgS7GmGetK7KaI6zifX799R0QvYnr9nXYIGT3QUbFg/WVPdOgOFvEC24VLRRgZL6nzAE/irr76WUhgfZkI1Cdqulk9sbWNdHVAocl8sLupQPjw1aWvbu7Z9WLb3f/6nNjF5iT4/S3TSVmtWbGV1VeAYdg6oUalP8BA/PqaWPLV+UmZPxy0ndfDHAhMRR8dFK40q3vXY/FetxfsuLtsafuX4sKeztrezrQPy0Lh3rDZ14Ezb4tKKgKzTlJqzd0hjL3QOnCcqevdy7eFSOgYxTHgb5rc7e/liEPc0/+vfj6iIv9/zoQJgE1R70bLg/Gc8H6Z9nliJ8+IiooKu2whIYN+nWjuTtpmZGcsXSroit39ANe32krpeLFoCkBs7LGWLFPy2433RethLVIhziVaIXuejJhS4HJSOUUhxUZh277XH30992mhi03oUiKVWEEG5h7bAlmzG/tXdf2G5TE5dEwAOFKnHx2XV4rWaA/13795TOCoiKlSxUZHPmQHQAMXwvTfu2eHhgSwbWu2aiPiTalnATF9pyBLJnN2//62yA0aGSiIq3nv7noBTauFENm354WGpXtdXVm2gOKh8ikNs1uiuKGKh1rAnj5et0UxY/0BRJBJ2dABOleNjBXDTEbq5vWW1RsteLL/sKrDfuPuaPX/y2Bq1ioKesULb3mENO7DJqUnZNdEZMTU5bu1GwybGx6xY6teeurmxZeNjk/b4yYIdHlLbZ+RZD7BI2DZZaVzr3ddft5GRIfvNxx8LvJ+bm7EP/viPrby3Z7/4xS90PkTIxTyZmZ2zqekZG5uYso/+4TN1O2EnQ3elALhEQl0AkGWeQYMlaF1gDGQnamzmA+MvWmGwoLpNrQeGQnYVlJ8HcNzQuSPafwHSs8HymViHeYYuDnNQC/KIGhrrP+qFGOzLmNSZVN1GObfLqp1oHxwbGbZ00qwE6ZvDNsQ7eO689qqugTPkRx//xl68WHTyhxWYPIJGXUTEYKmoMyK2OX19eXUtJutV5Qhdv3bZFhYWJIibmbtqjWRKOUhkfExOTsnXfGX1pXc7cv4eGLCHDx/oszL/OAuS8TE2PmqX565ofhGkTvYDKnMAb2oInYUVjh482gXKIRZzkZrCXRMpK5aKAsew+aGjSAHIMomnvuI5ZO369SsiCSZHRrXXzF2eESGxuPTCVl6u2ouFRcskM3bt6jVlwDGG5i7NyqIHsmFrf9+anYQdVioCJxkbzAvCtB88eGh9paK6RPjKpjLqyhgaHtGcnL85L/sdbJ/qtbLyYN55/y2rHOxLbAARgKiSptxkIiPLIkj1v/h//9IDbjn71hsic3LklohI6Bg+8eRkqHsn2jIFgFj2ygF/kB1eq6X1IOb6cYZQyHloBGYsR9W+BIHttsY2Yx8ijzVc3RwAxAJdIwjrorOOurHR8sQO7FMBWCTTY0eMuiixCHa+1TsHeza6JF08mZSIinb9RCA8eSuvvnJbn3nv4Mi+e/zY9g4qlsiktL4U+vv1WdlnwXzobmGMI9RTNxEZJwpoRmDgxKP2gkzAYmQb3jTEUCr7yCEN85+fYc8ix1OYu/5MZ0XL/uV7d61xeGATg4M2Nz1n/89f/Y1tndQsXxq1RKpg9Sr3rGVt1IdZrrOlOgaXB7rDZDFVb9ro2JhtbW3qGUAOcC3UKBtbKNbJxvEMVdZDkZoSq7VV487OTotYHEawdlKVyJG5hn03AlXwnNgdJjIqdIpqHw5OIzWcIwSgu70XGAvrGXNV9uFYYsXsGfbVc0RFrFmUYaGOGrfrlmAUtX+tfmr9hCg2dFAyX+I6KDJDJIR3XUB+ewUeTlY9do3RXrcL9CMw5plB0MaOXxEVEDPgXF4bMO45WyvXJcm+m1b3EGQvz0IEFwKnUskK2Yy988Zr1m5WrHp8YBur61Y5LtvRsZ9sSv0pm5yatmyh3757+sIOqyee70TmprpJvDOut+7383XI36GGgviOriISUjtZ7QIMF+jG//Z1L4q/3PGAf7y7ia5+BMkpjU/wIYTbzFUIEeFzjG8FrTN2Td1o9167pW6TxeVlO8ZKN1ewdC6nmheSe5hu5mPfVzx71qkzxi+4JAQse1wUCyOugminG0gC8EZD9q0Qvvwsz4J1TGtXsIISudTwca+Q+PTU+z9wjP3Hjl8//f1Pd+C/zTswXQ9en2ECM0EB+FBwYPswPjHh3n6HR1LTbG5uCeAgOJoCCWAeBp5iioVOALlIBice2FQA8SkWpX6hgEThCvsZmExV0JR6AbjnM/DFAsLCGAEa5VOELAwW8NguDMNJMS0GNJHURkShBtuN7QEqQiY2gOXCwgupC7ncGzeuC4DAXw5fcBYFFh2RBHh5siHgDQpZQdELqK8QHroz8LrkOgkkdC9ehXpD9Eilx2JKa/UpM8vGTtHDwQrfbwpJgAY8ULlXWE9JBSe22xdHFdVSIvmCKwImdDbwedkIVTB12WcPRld7m0ID/X3EGHd4PwdM+SzaAFruNckC7x01fl9FKJFbUaupQyTmk8gflqwMinOFo7dU2NMhAKCby8P4HsuWqp/cjxO8QesiLmhVVUbFNIrrZHi2Tlx5m6h3oXQVoxAwIVQ8ggWR3IobdPdgK2VVULZ0zIkzWkRRlxBSFKyflPGRKzgRl0jq73o7KqRiuKBYjMBRL1FxHiDrjtOgjui1foKowE8YQIiDV2wfHih6qJJUXs2mHR7s2fHxvrp9uL+Alwym1ZcrOsDqpBu+fDPy/3eAz1vPewmHCF5AUkTrifMgWCQq4vteBHx/72dix8O5QOh4TyhwICp63/MioLX3vkbwBkVifO15UFjHz0S0/fH1QFYdzDMOFlnaVrMifSi4eZ/D4DPcqJ/onqoVNlgHMK/GR8fs8OTYLIEVGaQjrb4tjUcO76wnABcollUwcHBpNz2PhnkULF3cPosB3OOkmXDSNXas4OXv9yiWkKdgWe+zO79bxPuhn7zA2qj3Pvd2/fD9CCRxiND1x/HTk3/gBevpWOqCYbFbJJW00vCg3ZifV6sua8zS4rIsyQBs+R2sS0ODwzoYRCYFcOjl0nN1ZGH9FPDDrhIytrK7xahnJalPQnaBF3cT6G9C3oEslUJHRSz2z+SYuFype81unceecnoQ7L3X50HLM3MtrL9xTDJnI5immdgF0E+BOsfvKW696EbB9b/9h39vG+ur7j9dHLNH3z3qts3v7+5pbZadUehUuahy6O3g6H12/jlYC7ih7LV0fmUtl0jazPSgvX33lo0Qkj02YS9frto//OYze/O1OwK1x8dGLJnN2fLSkmwPp6emBAROjE+IlH34zUObnBmzQglgrWQff/GtffzVl1ZtVb9HVJy/p/EznidzVLb3VNUiEHu+Ee9v773tfUYXPi+RSXXLFdJ2885N+zf/47+14tCQHVfYL4s2OTyiLrat9Zc2MZCxjFVsY3vHask+6/RP2ovlLcsmU3a0vWNPH32r8T00WLK3P/iZ/fqjz+3BN19am1b/lgdFatz1WC5GokKOPLIGOrV+iuvxmbWwx/pJyt9uh9TZdaJ3jOm/6WBtnhIVUgCb2VB/wcaGh2xE3urDqt8+/+wzdYeiCmZdLOSztruzIyCXboqBoSF7+uyZlM3JQsEWV9dtbv62vfHO+5ZIERqcsaSl7aR5rK4y6j187/H3Z7+ks5IcgRimjTAjnfR1ANCJdRP1egawETEKBz/yvhingGfUCI26ba2v2ebKqlXIPpE/b8qGISqKJYlkUGkTsLq9vdcFG87Pj7jeAcyft366aC7FZxjHEo8rNsfEe346zs4TFVHd7DVsbzPi9wi0C8K9457nPuOnQoGzP3vW+un8Phpf2ytO8OvE9inaeLowA5KCvZJMtb7+QVcRyqoAGx1Cab2joo1XecgzikQG9SoWldE6Rp0XFxAVrN1xX+8lKhwgdj9zrcHdesVr/Eicd/e68N76/SmU7Gva12U5qnXchU4KCc9k7U/v/syWXix57k6+T9kNgFWIe+j0gUy788qrtra6rvMMORYvX75UB+b62oasyrB4+hc//9AaACUdLBu2bHNj1V4h56E0KP/7vf2KMioeP3pkg6WCDQ3k7b2379rR7rayLYRw04XcbllxYNAOdw8EfpQGhn2uHB7pGXz+6QNbXNqwsYlRq7dbyrR4++23tPWRW/bVl/fVtVBrNW1rd0/bWLHQZ3dfu2Mf/+rvZU8EmA/Hv7O7b+WTus3NXbGlxeeyKxpEiXl0YNPTk7r+XJ58GPzSM/b8+bLbsJFDAICS6mj+YVVULHiH/OzMlE3PTNnD+9/Y4osFZT/ce+MNG5uatNWlZXX+QWBjbVOt1Wx8csaOyidWwc60xnmMPBQH6BB3yS2DMRPsamInPbWw7JdiXlSw5eS1dMQQ0sozpJudsZHLkIuDSj2lcw4AGbWfbJ1y1PeAkkEVHOzHOEcCSiIucatdJ+1kj6JuY88GVMdyp6WOFKYr6m/sGF34UtQcHRsdFSlD+DoAHmdZ1jjmcrT3Iywb+xN2M+ycitmUvTZ/xaYnyOfr2LcPHlrlpG5Xb8zbs+UV6ysNi+AB1J6cmhBAuLt3KBIHO7H1jXVtC96JxDpY8E5R7lXbyVQCfw/LZY1r5hdgGH8P+MpZmH3I7Xc8H4E6WWHEqaRl8074cS/WNzbN2jKeVQconYPpTMKuXZ2zoz0UwKaumvf/xQc6m7ZOWDeaVjmq2NHBoY0ODVmTcOEM3Sh5hXP/5vMvrc45FuvdfL86IDjjzF26bEvLy6oZKZuxw+TzERybL1B7Z4QLsGdh+wTh+MEHb9mbb961avnQ2g1yKyRj1vm91YaIQoHfsb/4i78UwEwmCmpwrGTUNdYmQ6Hhorzg7ctYcvGk+9wLwOQ8y/k6uEqwG/PfjFdqtNh9Eb3wPcQ4BBenEq5MDzWAy3N8fZftD3sF9kKye6JTgcxDFxl2xZzBT1/1vKzE3L7Y3Sy8Q1nduN1NLeQltZs2MTIs+yc6Tqjtdne2bH/vWKTT5PSsxsTy6poV+osKAIb4R0jQtZrO5tQJKaAd0ZyrQnTNsl8TKejB73JS0Lj0Dk9IAcB1dblESx7NV36krYwJFPiEab/z+rxVdnaseVyxiYkpe/JiybYrNRubuWSNRsLKhx52nuTFGRc7co6TtWzIVdzbOxQRymfEsQCilrlN/iPCKWoanq06HPJ5nddYt3KZtOpxLPE4Z8uyDVInmRK5PTw6ohqZ2og5Xmu47ZGI7rqr7yE+sR7HVhtsgdsEZsJ6wf4DeKzc13ZLtZbWLVktuV2j75N+RomgO+/BGPCMKUSjiFrd9kv7Xjj/ucjCcTIFPwfRlvAL2W4D+Z92n7ttUhCJha4E5j6AvncW+LhnfEL85+guCKQSNnjMda7NcbaELA3JWkGPIrwPUXKro468HNZQYF3JjuVSCbtxdcaFNKVB/Txn582tQytzj0oF2z8q21G1ZhXEN9yOlIePx1K4W+MEolnkTMD7+Oy65tg61hVEOB7i1rB+Jndyoqf3Wmc2t41y60BfG3EMkaCR9VLi5CDgaGPLmLQsxXa7Y6/fuSWscXF5lbYtZbvxpIRdZtI2Ojxs+/t7qpv07BIJYZLKwq3VnHAnPyWf95zUbFakPAK/YmnAyogW+vusfuI2Xqzr/L6IZyJw1RrcckHyTx0VP1Th//T9f9J3AKIignb9xX4p7qanZ3QQhUBYX1uzF4svrXxM23VWym/aZFF7sImjWqQYYWFTJ4Y6AjwrwQFvNk9UA64o0CElBD9FYoKFOC4iKlaDqkEhoxxSxJo6oynv0bBo8/s9/I+2XVfpsSnwvpAT+DFTXHIwWFxa1qEES5iJiVEVgHRPrK1teH5Cqy1lia9bznhT3DD55cOYDrY0APvyPHRLJDHsGV9AWGC1gcvbr2NLyyvuQQeBQXGhMHInLtyXnevDKoENDu8+zwthk9Lio03JraO00KIK5z4H/1MOjjwjilDUHvLsVdiQ4vUAACAASURBVNF8rO4NSBMniwhby7knKy3sQbmiw+lJTdfNgSAWhbHYUiEbNlZUTPr7ALixkFNoUjDxTADfeRact2l5xnmX564gbREUWFR4+71nVDhRwWFGxWEIb+RwTbEUwVbuC//9ByUqlO+QEbgEcaB7F9p24+/qAmPBvzgeouOYPYWZz07/LlkRg+DDpsnYiEQF45pnocIKz1c2dQWGt12NdFJ2wqrVEQjPIRdlHuBaN9U9Kt0DtKsNORTCZwiTAAD85xAV5xe0XuIj/l383nlVfi9RgRXC+dfHP3dB8QDOxEOq1EMhTJvXAhjp70I1fhFRQSGh4gkf4ww+6ByGsgrlg2ggJ4H1AO9/xjtkZNR783MEWB1UCRykUCDfo2gVWUY0dFiiwJXtRLIjwA2FEu/P89jd2bZOl9j6r0NUIKXqVUycJZZiSJ8XpLqHAQRAVSiGNnxd+AzCwceB8AC4YyWWTdsoHWnXrykosZeoSAmYMhVWFFDBd8Whsk5LwZ/Vk5pZy/NtolWWVGBxfApRVH9QyEvpAQR7OpocfjtLVPT+5HkldTwExGv2w+hpeN35sf6fQ1T0qq69IA7UYY8VGst2O9FQgcqhYKDYZ//uf/13sg4DrD2qmosAXrzQGrAv5WDomlK+ycXamN5n1/u7/XqcqEDpJKS2lbFsImmTE/325p15GxnE6mfCvv3uiX377SN76+5rNjJYVFgmJNSLF89td3vHZmdmpaSbGB0XUfHFp5/b1My49ROQmi3ZFw8W7KMvv7BKsxIOAj25C+fIuN+WqOgl8HrXDj33EKbdC+Je9LwAtCDFcoWkXbk+a//9//BvLJHJWjqLXdGYFTMU9EdWOdqzfKJsVt+zXH+flSbmrJWfsI8/e2DNesfmr123+199bR/98m/t9u15u/vGO/bVV9/apx/90hqVQ+u06qFLKLSgh8OQExVuOeZEBU8RUsPn5PfWzHNExXmiuJeQPnPtyhFAQOGhyYBsZJGMDpRsaKBkxf6CRBDs98+fP7fh4RHZHPT3F+RjTdgkys+JySmBFOubm/KsX1hds1S+z9758Gc2PjlnlqA7kxbzlNWbR/ZyZUn1IRYtHLCcqDi2oyO60iCK6Q7MWTaDAtpV7Si15Xme7xNRgfqY2oBcDZC2dqOlwz72WY1a1Z49fmSHOzuW7rRtaLionCFUp/39A/b02XNbWcU7WxLU79Xf/60SFReRJr8LUdF7wT9MUvhK2UtUpLF/CvskHRW5fFG1NDUo9U8kKiQOgagPFhCRqPCMCs/SYoxGEclpR4XX+j/UUcH6F8U3/xhREdcL/s3PJVMdeTc7uOqKcEDXSLLw7w9vvGXPF57L/mlkbFTkw5tvvimQAGCXnxEQcHCkgz/zAdJtZnpagJJbX9VUT1NL8Od6HduyXRscKKoronqCbZPaVO3B/ftWyCZssJS39995w8r7O+pcSOYylikU7MQ6UlOW+opaBwjUTufy6jg8ODqy33z0pdVOzK3NMmnblXXTbTspV6xRgzBCvNKycq1maxtbugZqZrInHt7/2iZGh6XahsDbOyzb4XHZ5ubmBNRxRkklOlY5OlZQLrlnAB6AbMzj7757ZplsXophuspP6id6dgDMuSxqUrqlyzY5MWbTszOycHz64FurVCvKDACEmQpE9vLSiu3u7dvaxrYd15qyztrZP9Q9Qk3MM9RYCvsiFAJ1Ah3r1N7qXg/gp9f5Sc8KxHqHNTSF2Kpt+WAfBrgoAVlYSwEMPWfCz58ApwjmAM6iCpUzSoSn4hhkvKszP5W08smJznMtFMSAd4D3GToOQqUPSJvP63rc6iat86Ofj7yTOaqgIY/ITmBt5OxH923KmjbWn7diIWeDAyVbXVmW/c7Q6LiVa207xj5ra8cmJiYFXu/u7Qp0xyKE+nNjc10ZIXxG5i6bCuMagD2ZcpAVAB1iiHVZxA40cLDD4j19/4SAwyvfw8tdN+iiCHfAc3Icaz7ANO4DdW+xP2ez05N2UkF81LTJqXF778P31KUvQVazo64GguAhdxh7pjN7xxYXX9qjp8+srzRgx4gzMnlZmfDZb1y/YQvPn9vE9LQ9e/Hc6s26DQ4PCYcQoBdsi7Uv1OtWrR7Z7MyE3bw1L5U2NqzVckPqfZ4NY5vOiky2oI4XxiUEjtwGAiiLmAlCRJ7/IvpRontOJOspz5Hcv2jXg9BSltIA0zrvuz0MZ3Q+k7rMQ1cZz4ef5+wg6x2BnMGAKIgQAP5lIZVwm2rGNnlLMRw3ru8uUgz7m4oAF0vysyKbQkaFbGqDX7+uod20/nzOZqfGdX9mpsatL5+TDdrRcdnWN3Y0phjz2L+R4YHFYlR7A3byGeXUEMLqmb9xrWVugkOImFOWh2MAOv9zXkUyl07b8TFdbE5au/izoTnZUr5Kwpq1mn3wzh3rSyRsf2PHs6dabWPkdtLYbGXMGu7u0AA/QKpvEA4xOxXrZg8XlspfodpOYrtS3oF+YQ1gJLUTrWsQFeAVac4sxX67dGnWDqi7ZRnVlvXY/sGhrEOxDpNlY5JnwfOiM9DHjXCPRsuyhawdHB26jXSdM05C6wr3ELKQc6Jnk2Cj5g4VvWIcCWLVcYJVtq+XEpaG4Ht10gQcIopIqdtip020Q+Q+qcMj2LLHsaN6s6drVOfpMMjcsQRSwB06ZAMfQflwnonnRwQA3Ed+XnicwtI9O0XWS7J+SqkjijMytSgdh43qsSVaDZ1rEh06uEo2PFSyQn/BnQuSKfv6/kPbO65ag7pC/pHBtkvjOoRkBxtrnRBjEHmos30VC2eEkOPGtfE8Y71y0ZnJcYdwpoSs6RHvxawrETbBFjPVduIF3gxmlY4RiIXHz56LqDBEjpAGslOvy3bx8PhINTj4nFxHWgSt92vMQoIztrj3fDHmwBrK1bK62dU1USgIn4uiPsYQWBKEhboW1c3nGB8E208dFd87Evz0jX/qd+BawkOSAPKmZ6Z1IGRSLLx4bgsLz1UMsbCgKkY9wqETH7pLc5d0wJG6PnjcSd2UdtAcgJ9FE+8+lDpuU0Q7oFsosYlrk6NVr7/ffe+UheFFJl9Ks68SYkY7d9InYejW4LUqGNVlCNPM7yzoAH1p9pIsdmhf5Bq++OKBDQ/32xtvvKHXLDxf0MGdLxZ3PBgpnCmMorc/n5eFgr/T4gzok/SDAxuKCt9k0vr7ilpYFEBEAW1mj588sS+++FZsqDZ0IATZiniInuc8nIYfqhMgbDxSMASFkTpPVIw7MInNQtw03MPQO1QolCm6WQgpYihCAOJlg6QCyu/lcflIRIWz5F5AiKiQ6qzi3RrBeiqqAug24Hrl80gRUHc1hYe5efFPR4kUAtrSvUUWWRjqSgq2ZpOQOA4dPOOzHRX4nvuhN26wXkj3di78oYkKVJ2MWTw4GfdHZYLE6MQBgMUv1wFC7Vmhu6VLVATixPHAHmN0CYNPldSOVAXaJVhIXURUDA24wkDqWKnt9qxSdn9kaQ5h6JtN21pbt72d3W7409l1x1UZOmJExUBQaXjRg7IU1djZbosuEBisny5ay86THr3gYa8KMoKlEThEkUeBcv718c/nQXK/nacZFRGePZ9RcZ6okNpGyi8UHWlZKBDuBZFADoCP97oOb1jsyGcSVZ9APgetR4ZHbLe8b/lcyQqFkiyg6KhgcFNY0yHE/CBMELsuVDnYp5TLx/b82VM7qbh/5H+tjoozIbGho6D32cW5fR4QVVt2T67KRURFfJ8ziv1kQoF7s5fnbPrSrFpzuY+xowKigjFGqz7ray9RwXqwvrbint9BBRuJitA57d7Q6tgN4apdK53frqNCAEhYT/0/fKzHKdrbUeEghauge0Hf3nF54fd9gLsiKdrCnLuXFxEVXEon4epf8mfwZ/0P//4/CFgGiPrk84fyuMaGECXX3k7IPrnA+umHao0IGoYr9vuPci3hYdqRqBgdztmd+Ss22F+U9dNX3zywtbVNe//tezZUKtnE+IgVBkr2+PFj293elf80eyCkd3++YJ//5lMbGOyz4Ylxs1TRvvz2uX389VdWbQJ6nLV+6rWnicRQJJ17x+X5jgo/J5wlZ7QGad31UMfuV1hzzz8vV8Sj2mvbxMyI/dv/6d9aX2nQWp2sjY3PWj6ZVc5CrXpg6faBZRPYTAzazI07Vk0M2i//4Wv5bd+cv6P651e//DsbGx202ek5W1h4ab/6m//PKke7ZtjqiJD/MaLC9992B9uI0wyBXkLGO+H8PWJLfpTC9ZIUcY3tjtVW7ELlgNUU6J9LJYOasmT9fQXtaWsbG1bGpmbEw3cJPcVbn3uA4GB0YlKCAQCdl2trdtRo2OtvvWPXbr1i2VzJOkY9RkdF0moNiIplkcDURtQk3H/EEQC6qGg9IygvAQsz8/jo2I739y2P8p3sAAKNZcdR0+eQ/WGTbMKWuj5LAwWrVo5t+dmCHe7tWLGAQKYgX/uBgWF7/OSphCcCq/8LExVeu7mXsY+zH+qoiDZOPcMzHHq7a+oF4/p3ISrOE3WxJo7g/uknOEtUJAH98NzP52Tlms5gReChxBK01OuqyzV3m8GLOih8XfBy1vrpIqLCXaxO6yBqzWj95Ou8dwlfTFSc7Qh1JWQM6G4rUBcAKNbLAoTCZ2ec/2z+bRsdHrPDw7JAZQEjAQRAvICNDPUtHbWAqqqJj1Bpe4gqdTPChkuzs7JEk+L78rQtLb7Q3v/g4WN7+9337ZNPv7LZmTl9H6JiZmpYa2jrpCz1P16IWMmNTU+p1t7e2tEZACUzdiV75GUVS/bNV4/V4YXt0v7xke799PS06vZCNmfffP3ACsV+fd6FxUVdE9f5/rtv228++pUU03S9YUu7sb1rG5vbduvWLVtYeCpxy5W5S8rQQpjFGjQwVFK4cDqVtZWVdTupteSST43PPlXHJiadsoO9HXv37bdlH/XtwwfqznjnnbdkQfHwwUOJ18ihwIJibu6Szd+8LWVss52wv/7bXwj8zHCPg48742RkeFjAjazi1KntliLcY+o2wF1ex7ohyw5ZyThICwAGEUoXOiQ047DY58HYAPRsw5wbuX9a79bXQke/d7K6ICwtwDCq3wHCZXerMQRRw1puNjY6LHB+b3dbmVGIxxgXsqDiLJTNSwgjKxjZSnkIOudUt31xW17qUvb7rNT4TZubGrfLU6PWOqlaqdSnMXB0XLWJmVmrd1K2f1yxw7KTgNSayv0jt0AWwBCEZZECshHOZd06JIcIBwCLuduwvYM95U5xBoQsYR0+OiSnDyDMO9cho7zLHtFg2sdaX8EKfXQRI2xDiU4YuHcmu41yw4r9ZF8ULM+Zrlm1mZlJe+/Dd6x2UvHnhMVSvSU1texQw/W36m0bGB6zX/zdLwRA1sgiyeTscJfOlqzN35iX7VMr0bG//Ku/stuvvWq3X32l+2yp1RAk8rmPDvZ1PsJK6+4br6u7Q3hDBdths3KFMPppW98kZ4NunoxVa3V9H+IGSzAIoIOjA5FqAwNk9LgDAUIa9ivGBLY97C0KaFaWCYSEK8kZc3xfa1mrJTtf7n0cSzGsXYG76lTLKvyWexuzNxloYBpAq7yHCLOs28UU8mSFeBeSMi6C9Q6/m7ElUkP1HXWoEwl8L/ZCKx8g2ZF1GfaO+3vbQmFxnIC8IJtzbHxC++ez54ua/5CndJtgAc779ZdKnjtFV2NUmIeO0WjFw1qkE0/Ix2DuyAqKTrmQeYqFN+NXFseo1EVYJKx5Qo5nRja8d+Yv2/zcnK0trdr9bx5a/9iolSGUqRNaZvVjiNWExkcn4w4d2Ipx//i8PH8yIJxwdAvrahUAFwEowkqwIXeYgDTkc/IswbE4BoyNDdvN+RsS5ihfNJdTl+gaYg2Rno5VARbv7h8E0WdeYfARI2LPeL74QjgaaxN4lgPLECFFiVWZq6ytBGu7I0CkBH1/kxVWEPnGZ+8CVT/bsj+BQylvgbwLdUI6ecJ9VWekuhSDZTVIjILdwzPqAeB1PgziPu/e4dlVXTSWCBkkwQLJ93hfcyNGFV1O8tgsZshV4R7VrQEIHyzjICmyiABHh+z2zas2OTZiWxubtrW1Y6tr61auNLU+9vXnbHh83JbX1m2/fGJND/VT9hvX6PgeQuYe8WrIUvXzWBz7XvUIfwjivCgAjpjZ+XNCxKzCQO7+rLAXQsbpjqo31MWoLJ/aiQ2wPzGWrWVkwdy+dVOdkMwly+SMy4eA5lkhJJ6dnhKJBSbG52ItY89gbeKZksPG+uy1UVu4JbU0uCqCBtYGCA322oivsheSQwQGJzeUYOUHUfFTR8UPnZJ/+v4/6Tvwr29ct+mZGW3OHCjxTFvE+uGoalNTY9okOKgRBsOmMDY2Kh9L1BpMJiYRhR6TuMsEt1yN4cExeJWSReCbrtrURGjA4jobL08+BanBzratUKBAcJWu1M/aYEJwdg/o74d651L5GdqkuQ4OA3RPoLxjoZufv67CjmsjUFKgPn71ubysEWgbhKDpL/bJ49YVALTSiTbVJlBr+8EmbhysOrQ2UgDhAY1/8sbGht1/8MDWN3cF2KntGV/44BHKQtX1AA7qH95HuQ4JwiJ984cplW9laEFjIULxxX2MIYIAKCqyQuu+/h0W9Ague1uwF/v8LERFvuDXFw+oHE5lQxVsrxQ2BlvOc0BBFJQV8T1QwbjS2pWhAn3VLQHw1vQAYmWGcN0e1AZopq6VQFSUJoeCwpjiIaih1L4M4OKqhgh0RXBLxEUABt16gOfiY8SBOW/VdWsfk39ureyqoX6sn0KQZFrWT3nPPsnmRE6VK8cCLxkPjFGRZryrWlkdPPd7Gj3BA1h22kHYXQMiaBU3zbiNQmANDQ9JIcUGRlHKtbExMfalBKnX7fBw344P9nTQ4XkSAI9inywA7Ml6rXviL405FS5K98KFG+O3xq1xULF6x8XZ1ke/e55R4S//vtq8V5V+lrjwDNDuV+hG4lmhlkMZe/4r/nyXiGBud1sxudchGC6Az1EtH99HqongLcnfSTEnpZQXqmpjJyStkNc/eGhSBHDwI4wQxQuKhIZCHBlTkHgZaxhzrKiAUQ5Srvb3+UqhzTjn8MecGCgVdViku+L5wlM9M4LV1QET7r2PSe64dzD0Wj/5tZz25HTvSY8S36/Rn6GeY7xhFKXedHDaS9PTyhqqNe9N4N7qPnJPO9aq+wH6B5/JOWCtO76wLCqV7Nr8vA2NjqmVHqJi+cUL29pYlxUABdjQyLDms08eEHreoW27O5u2t7sr9XPsqNDfcJHdQtSf5Vmw9kzfyOkwO0+4Bfm6j10Piz2dkD3/KXu4UxDtvBo/An0XERW6lljsR5u98PHi+/QSFfxWAfLKVHFyhDUYguvP//x/FrEOOPLpp9/Y4Oi4PXm6YIV0zva2Nq1SPrREKvjm9zwTV/+cXXR6x87plboNjdtnsTCmNA6GBvvslRtXZP3EAePLr+7LZ/29N+/a2NCQjY04UfHw4bdS+tycn1d2E8QcIZef/MPH2heHJybN0n32zaMF++bxE6spN8c/19nPc3aMnyclNKzPjDnvBuqOuzjuw2ukdjrLYXT7yvQ+PX/HEOC+j4wP2Z/+2R/b5OSMtVoJm5iatkwya0svl61tdWtWtq0v5Qq8W/feskRhzD765IG1LW3XbtzRI1949tSajZoNlQZte2vX/v4v/8J2N9fM2lil8LNBgNDVqXlHRWSO/S7wOicqfF6f3i9sH5zzhmDzV8eZL2sH1vTwb94zHsYAg5jPMTCZ410+m7Vx2T4U1VXB2rXyckWHYew8S/1FD/y1tu3s7lpfcUBAxf7hsR0eH9v+0ZFN3bhp773/RwogT2eoSbB1cBFErX5sa+vrqrPkL5/r805AiIrDPXXQcnhSfpkEDmZlfInpqMhkBbailuNZKusqKMxQ5OLpz+cCiGJNp6OCcZjPuCgEC0oA3qePn9jC0wXtl9z/3q/u/AgLTfd+aqM6nTsSFQThSNdsrMtD9GZW+JNQHSL/Y1/TzixGWuvDEzu/Fvf8Ts8S8b4xnythDVfWWlrrlsaHat3ucvM94u57xJzsEBhDbj0T9TC8uwNtKFw9Q409EsHE5NSUrA55sQ7lqaQO5fwjJWoQToiYlcLcfb1ldRP27CgmiTWDi2q4sFPrJ9lZBrsdgBXVtKGjWHWH7lvMxwpzo6fL0tdR7CVaEh4hkuIzAaAyJjhHcG3U2vemXrHFhSUbHRu3Ql+/goEZb8svVwRKAYZjNQNxgAr3ww8/sF/+/a8Eti8tLdmVy3M2NDxgU5NT9uDBA9nf/emf/twWFxdEZJ6cYNGSseeLL5XzsLy0aLm02fhwv9199aY1TxAmpSxb7LMEZ4UgnkBBfkhgd6uj8QswAdjwN3/1a1te3bPr12btqFyxeqthr776qlvgNlq28OyFXbo8Z6sbmwL9y9WKDQ0M2dUrl+zRw/t2aWZSz6tUGrS1rW2FM/Nc2YsJPEbVv7+7azfnrwuIZgo8e/rcpqdm7cuvHloimVEXJCD77Vdv26NH32reZcijyuft9s15hd8uPl+QfeulmVm7fe+eHW5t2bNnz2x9bV3A3cDgkGrpy1ev29LqulkibasbW/o+nevK5JOYqua1aSplh4fHOnthywk4y7XJrhdLjKA452wJGFOl7SSoZZkd6vypebc46xDjoClrlWPV9qxB7GuMG9YhBcATlktHTOgkgBCplN3ahrUA4oz1h+7biZFRy2QAFcuqc5gPvI7XlAYHZJ/F/OB75Dbq9zdb6lhhLkD4EEqOtR5oKwTJ+FDRpkdLdm1u1oaHB+3l8pKCjfPFQTtpdGznsGzlak1gH+dRXACwjJq9dElCsI2NNesvFuzOnTu6hqdPnoqgwZ8fqyOCtPcP921kdFjrLjkQdJ2k0zndX8gTBIM6H2j+uU0ygBnPpdluaNxwv1kPjg+rwRkhadl0wkZGBgXss69WKkd25eqMvfnBW9Ykh65W8/Wi0bZahXHHvsSZPmX1SsOWXixLcVxE3FM50XyvlE8kgHvnnXdteHzMyOz75PMv7Pnyks1du2zXb1y3ibFxd1Cgs0lqeCyLKzY4WFK4vT8XOofSIr6o2QlwFuie77PFpZe6F7lCQaI0nXs7batUy7a8vGhLSytuF5bJOqEj22i3XukvMCbL+rer893e1C2EfM8BhOZZADxKEZ/Nar+VsA4hirI4OKsGYYy6K7wWZLxy7pclF7iASDrsgvxcyPc4gwvARHQRyCZ178gmyF/DWQcbaledu3ABkh9idajEZ+9o/q+vrtjWxpYdHtW0RkH87x0c2MDgsBXIz6lURDRIQBpwGN8bUvo+c5HrZz4xliAcoy11BNElGAqkobqpQmcwa4QXQwC4KT8rqZOyae+++brVjsvWrrVsZXXDUv0Fq7RaVgGoxe+/7VZXdJV1dJZLWL3quaMifrQVu90WOJSslshDpXuPsxtjU3ZHni2q/SKVkPiMWuj6tSvqgtvZ3FQNw/Mf6C/ZwdGxng/dagoXFzHl1nXcCwjuErUTeRftlm3vbFt/f0n7mzIdqlifIZjLC1eLOZ/gZNrzYp3AciircLf84qFydu61P1eX2EnNOx9ChwDd2J6f6ESE8Bx1TnhXgbAzXBnCWIo1Q293BOOL17m4zJ0seJZOWKZk/RQznDgDcB81PgOGR3g345zPAdnJWAcTy6VzVjk6sn46i8gTSXes1F9Q56KPG663re6eTTJh0xnb3j+0Cr8bjYTO+N4hF/vgovhOIgfDocTno2N0Xp+xfotcVGaD5+ZFYcTp2c7ribifeJefF2MeSh+7n7D949zkrg5YYXLdN69dtdnxUWvVaxKU0rnIPFrf2rF2Im3Q3WS+cE9436nJCXVU7B+Q1eprL3UQAmeuTzmXHSeHwIK4Pmz+uBZwOdY16nXtYRy0LeEZFaw94K8Q/3R2IfDO5/R+P3VUnDkS/PSHfw534P/6sz9TQUVAIvkTLPIo1ygAN7d3vcDHV7JQEFDH4Tiq7jkgAB4zAeMCAdMdN3PlMdDmpkXY22PjwskiGjdCea4VUe75l2wrMEuoMfnyQeHu+RCngLz7IdIqNTGJxVO/yJSlxUV7ubKiBXuShbHQZwcHh7azvaNARwWooWwd7LepiQkprZn8Knjx4iSIj8UQDzqhTL50dQCOAkDPe2fSHjaOHdbK2po9fbqggxHsfSycYbvVdhYWVnU8sEgH+xW1PxJYpYUf2ybf9HQ4QwmkAHIH3/g5FjkUA96q76HjfEWvzOilGb3w6ExxP0wHYyENuC6eQVR+UIjzu/lMfE6Btnj1CWvkdzR12JOFgDo8KOArGg/82YkTt+OimExmU2qfxvopnUbNUJf1E6p2Bbl1mjY4NeJt+wpEp+X2tDukjT1UAKsiSdH9N5V5UPidBxm9DNIurfFGcSWiApC6v9+JioQH7uFfrHbQbM5KJVhrFBnkqPSJcIvXrwO/edBkdzMMvswXzv3gmx/BallYhVEtomJkWOMNooI2bQpeNidvvfQwdLxty/t7KrI89NnbPjmkQ1Sor/ncVwQKTlXkZ0OxVZw4Etb9OgN4KlPhh8O0fwgcVSezbk1oJQ1iU66FriAdjOKcDmr0+FnVTtsD3PUWUrEbJf5s7++X7U8POcLPqSWZeSYriJTWDIpJPe8MxWtB6l8CCmnZxbbODzYOGmnccGgLwXAxY4GDj6tbEurUQo0c1VbKpLGObe2s2/rqS2vXGirARbAJLPflw8stzaawnsQPfwri9j7OOHZajnF38xdiZw/VTzO890WkUvee9XBpsQNA6rieLoDfZv/S78DfeXTMrs7ftHxfUQdkQBAAjM2NFbc0wmqmWArZFJFJgdAgxJD1d0vAoFSy8Z7oQTrJxFe81xHM/cHPp8DW6Dnak63xA2Hw8X2kSusGn/tk6AX9zhIVZ58Pzzbaj/FzvR0DgzjutQAAIABJREFUcX3qHet64vFAgvVhKiXSjL3qX/3rPxNAW2/V7bNPvrbBySn77vELSzU6Vt7dsnr92CzdMmek/Cuudz/2zE9fewqE+gHW1eAUspemJmUJAFHCnlWrVu3eq7dtamTURkdGLFfst8ePvhMxeu3aNQUMojCD0P31r/5eewHESjORsS8ffmdLK+s6WMROh4s+33lgtffP3kDxPfbBZ0wMNQ7k2oUE0rn746sRBx3/4cGhAXv3nXfslVduS+0MONZqJmxxbdlqrbK1T8qWbtQsk0rZ7bv3LD80bb/5/FuzZNZmL88rjJPg81q1os4S9r6//6u/tLUXz81aWBfhW+zdV8pW6X6e+EnC7A8H05hB4Wejs+t0XCO0mnbY8xNGttFpJ1wEzH29lW9xeLYoJvneQKnfhul2KORsZKCkmoR9o18Ea0nEE3v85s6OrF9QLm7t7ckDH0V0/+Cgvf+n/53CKdn7URB7e5J/1pPasepE1tdBgMg8wEBbIOHh94gKn9ccrACGAaZUf+lgHn2j3fs3qvN5xnxWaoODvX3b2tqQj3Qml7G01GgFW3r+wh4//FaARUKj7/SrS5QFopYl5vv32UnRqGmU9KLHXvB7tcWZ8em7+tm57qpIjdlA+Me/7927qOeiqKB37ZEQgoOtwls9W0w5M12yQq7HZ/bvM+Ms2n70ACC9hKGujd+B+CaVUlgv2XNYy/A6DuQC4RRM6mIiCYjCvOM1AqVEVODj7XZmvUSFkxRu/XQ+o0K2ibLWdEqIe0Xgtdui+ViXJVUAHc6vIZo6qbZU6F2iglyCYP3kJEza3p69a0+fLEi9SrAwn7W/OGCbW26bxM9fvnxF4xGQ+rXXXpN4iXp6fW1V4cTUWW+9+YbmDfXsjWtXrVw5UmcwREWjlbCFFy9tYmLadrc2rD+ftlIhbR+8e9fK+/57ICra2MUmkyKjG1IQFzxTIZWW5R/nhKePluxgv2r5YsF2D/Zkw4Q1G8AsooK11Q0B4zv7B3ZUOVENPjAwZJdmJuyLTz61+euXVddAfGxs7wn4vnT5si29WLS+Qs6mJ8fVSXVNWRaoxd0aqNno2IMHjyydzsvCiLUyk3ef8pMK1paQmgM6M7377puWy6Ts2dPHtrG2LgLjytWrqluphda3tm1rfcPWsNVstK1Sb+of1haeiYOUWqzcax7gs97QMwJkjeNG5yZLiDQhcwIQmHOmupuTCfnl88V5EvB4d3dPwiKyVtbXN/S+AMVt/sd5qtttw7hMWbPe0L0SOGcWREke/MvYA5CjDiGjpF6lW7xt1XJZdSzz0M9bTRubGBdIKf99MvqUmehknwfkIhTyEG5AsuEB6v26FVJmxUzHXntlXsKWA2p8pnQ6a8e1lh1WanrGzFX2GNnsYk0zULTLc5fs5u2bNjo2pO4Xui753bu7+7axsWXLiysiGDhTQwxh28TcyqQRXqHYh6zkUp2wdJEXCmF3OgBsZd6qH77JOYQOlJzWIUSJ7VZNnRSlgZIdV6oCwu/du20//5MPrFnFArFhzVrTmvWm1ap17ReyKEJlXznROf7p8+d2ojNNIAUwH+yY3bx5yxZevJCq+sateXv0bMGWV1etUkY8lrHpyQkBnHSBsm8BDFI7sR+T3cH9RiTHZ6ZDtU1nR6uj/A+eaVaCwWBZzDkhBDojNNrfP7Anj5/6cx2blOXl/t6R9l0AW4BZfifAMeuv22d5NgF1tGy/AnjP7wJQjHtbJwHpRcegtmiB6jrHB7EMr8tCtghw9bML84nzOmdpdVwEgJ3XAiYzXxiPssSWAtu7EZ2giO4LPDOsGpvWbuKBX9afCXcnBBqrIkhROqroNGE24DBAVgWZTrLPljVYVQQWmIXnuoXOJHIY6LHMMT7oOKcrxzEPWVV3HCDXOa3t523WHdZFciPBAfK4GaQTepbz1+asP5O3o/1j2dt1shk7hmTFFouMGwk9TWOnlcFqqmOdOt0fORETbknNvfI5Sh4F67ZbZOPQ4dmlPHesr+gypduMNX10eNRuzl8TscjZRKJO2TZhwdQMuVusRw2tZ4gL6aTiLHh0QNhxTvUIawD/II7s5ocy9iTWyEiooe6xIAZljRJYH4BrjRl1env3VLQ8924WPzuwN7MvyqoRwWrEIdibg7WvZ4x6TqdQtJ5uA++i8DHSPbvo94d1s+3rtIgAahGIsqZ3Svg51Gtbx8ZCngv5d9gFdpy8U0YkGF/LbAhCvtWy2clRRTYhWoSwqRweW1+xX4JNRAF0k1frDbv/7SM7IMeBVQdckfDxEM6t6w7uB4xH/uxnRT+/q4QI3dV8xmjf5B0q3D/HHf0fJyq6fw73xQVlQSQZ8AyebxqbL8hguitqNbs6O2sDfcynfv3DGH6xvGyPF5aUwZPKFayOkwl7fSYlXLJ6UulagqlGFC6hZHgJFqIsid/HvrcNwZ1IuF17lXwtbO3o5mNMOykHsYFIWhlxYG+42ORyGrM/ERVnjgQ//eGfwx14Y3BIAD8TF79+FoS9/UOxowQmA1AwaVjcpMRTmIwr4ryVj40KsN2tmGS/QghZaG3SISfhrWvOJAcQvtn0zU6B1fL96Kp9sYtyzzYH/liw2KTZlFBGx/bLK5ev6GB1cHxou7vbCspmI7p1+7YWYCb8y5cramXli+/duHHDajWK3oYWEfw+BXIa6puswRK7qtMXceVQ0GJnKDVQndBNwqGOw3nFvnv0WB6cLCBsBTDwCmq2jjXwsI5+g2GhFegdLJ34TLE9L5IY7mXnm1g8HPom46Crs97NEKDtC64K9BhMzkJNd0UmIzW+W2pRZNGKRgF+moEhH1gp5PzAyn0F5OWeqguGNmS1ozprq+BsmHWpQRwsUTGDssHaCgCiICAzRN0TaFbrtGa75RP/prgamBw+JSrwBg0emw5e1B3e724svsF0Oyp+S6KC9ulG1Q9mUjoFX2UPLCq4Gi+Xd4/fhqsEPQCr2kNUMMZdicM/vWDKRXPfAQFXy8bOgF6ignAuNhjeBzac+w1xEYkK5l61fGzlgz2r4zdLuy2kWCol+wTaBDuBnDoPzghkDbjmeWDmD0lU6Bp7AFgReqh7Iu4TgDNAAg7cvYBO789G8K2XBPI56n6averoHyMqYnEVfShRwvEc49xxBUNaaw0KOb4ATmo1CjPseDJ+QAtqV91zfH9lP+QFBeAm6yDzgC4yEbAKGoNwOlYGAwUYRbqIxtjREvgKvwd/OKICEiMWPL33RnhAHAMB+5WfbVDZUOz+GNjbO6Z6iSMAwvGZWZu9fFUhZxyCISAWnz+z7a01y2bSIozxCfYDKhfuh4p6rWL1WtXVhVL49BAVgHodB8F8LfRW53+UqNBAuajz5zzwe3aW8r6N0E59/r7F+3kepIzv8HsRFUFJBlFxY/6GzczN2Pr6emj9T9nbf/Rz++u//ZVtLa9Z/XDP2u2qdVLY2vS2KwUw9XuK7e+vROoG6gHC48FENimAH/msDveQpajw79yct/HSoIAIgrIfPXokRSoWKHRSAHCzDz548I3UyhAVu0cVBWTuHZXdU/bc2nM65nvV6f7dHycqTgmirprpdyAq1NlnHsJ5Y/66vXrnjg2PDNnExLhUl51Mwp48/86sXrHhfN6K/f02d+OaZYpT9ukXj62TyNjM5evWbCVs6cVzWVxI1NBp2z/84hf27OEDa9XL54gKB4EECfWA27o14f5obPd0U8S1VCKIELjpAgkXJ6jLoKeDqJewkvJa1nehzb/dspHhQXmg92FhkMfiak1kFOGwIwrYHpF6eY929EbLdvcPrYptStsEVrz59jt27fZrrtZt+KEYUFk0TDKh9Q4rA9ZY1MR9EBUduiaC9VMaUCUfOip+N6KiTzYJTlRsb28pCBjgAS99gLjN1XV7+PXX8vL/YaLCAchuZ9q5TkHvzgn+2bFb91yHVByJ2rfCNHO5ylmxQFxLIuh+fm+Of47rW++eqKEROq9YMyVIYf9R50DYCjn5n/udve8R1YZxzvfO/aig1PuGrlLyGyDdGdtSVaNMRFFO2CxEBeronq5WLp6/5/fEwFF+x0VExfmOCq45EhUCDDB1gKhgH4niiNBZ4ePslFg63YP4AC1ZX3pN5Fl03ycq7tk3Xz2Qtcmrr70u645nz57bltSufba6smp37961l8svtUdfu3JNXQGEWa+trKij+ejoQF0NB/v71qw1FCC8vrEmUGVv/9jyfSV79HjRZqZnbHNt1Qo5Iubr9i//6B3l1qSzKcv0FxSObWnI6ZwlswXbWlmxocFhAfQovlGT/s1ffmSHBxWbnJm0asPzGiBS5AWeTNs3X9+3qZkZZU8cAxw2GjY+PmHTk2P23YMHdmVuRuMSIc769q4A2rHxcWUiKPT2pCL16ejIoPX1IdBy+65OO2mPHz+3ZIru4oIdoS4eKIqMIXcHscxbb7xhS0uLtrr80ubnr9rrd1+zo/19e/DNNxqXUT371nvvClRF1PbZF99oX5DMDKA8Qy6eB9QC3jPOOJdAVAyPjAi4ok6G/I7nR+YQgiF1U2AlQ6d92m1AqMNYy+KZkv1MQdxYHfX3i8yg3i8fHwUgt9UF41krqbcFwIVMsXjmcRC2HbLqCMut2NXLc+4AALgoQsIFZXSsbEvAl9KewZgFWJQdGecUbJrqJ7I/Ys9gjeHap8YG7fLkkE2Nj1o+m1IHD8/DIBOM82VanTo3bt4Q6Yta98r1K3b1+lUbnxizWr1qR4f7/ow6HZuYmLC93QPr6x+wWr1p33z5td1/8J3tH1SsWMzZyMi4HezTmY8FTl4AtYJhJXijroVE4r0IFccdwccM4cPMCQLX2X8B53MZz6lg/djePVJXw4cfvGF/8q/+yFqVfe2BkHGNGtcM1Ahg6gI7zn0P7n9tz5deijQgTwM7JB2x2wm7deu2ffSb31i5dqJ5MHXpsvUXB1U70tG0trqqWgQLLUQTdFX0Fwo2MT7uWEKargKEWB39bq6buYUYjc49ulIiWM3YIBvw6PDANtbXFCBNXg2E+wfvfah97bPPP9d4JhxdXUCNmjCFEgIA2Ze52jy6K3A/6dB2IQjdPC46k8ggdMXT3SJP/9AxzBoXgVbeX1bSGTIduLcnmiNMMre6dIcA7WWhPmZu5OmkSKeFyYBJyJ6njs12w+oad01lVHEeIoRc9/G4ZcODRWWQrm9uCecRTtPuWKVel70rtQFW31wX95/303zDBSNYI6v8xoq76jZjIlTUwdBS16Q+v+yM/HWAscx9Piu2gFjQcj8QVVy7cslWXixZsW/ATupNO7G2VbDUZL3gDfhcmay1ISHYP5ptSwbhBNcNGeQdRJ5/Kuu0KnZk7sShz9VqG/mr+/u7um8QFePj2GCOqIMM26NSf5+AYUi1cgVLOO962d7ZU4cX9/+k5qHxo6NjsvMCh8FGEVzErb8QhGJT7riJxEnpjPY/2agFzMSzuLz7kd8Ts1AkDK3TtRdiwoO4UK9FSBqyThljdODozB/ILPZscALV17ICix2gjuJHgjZaDDG/4tmY9YC1LpJRLhrw9TpmJ/B6agNKJLmhsAm0WR9cACH7KtbWOoR+3fqzeUuR+1rI2uTYoE1PjKlDA8stCELCzE8gVNOIoLO2e1y2E8hGSBKwKjpu694VETtGwuFBn8HzOII9dyyvOTvy/ZALyrX6GudYWvcsF85QOhf1OAwwrBz5A/choyhtacQTdM+lILqO7erMrJ2oi6xqpWJe+SY7ewe2tLpmrWTamspxawlvogsFISxE3eHhQcBQ+1TDusNMwwn3fF5ddHzl+/rk/ABQJ7v9KhkV2CxiZwYW5fZzp0RFwTt/lPGEDVr5J6Li+0fin77zT/0OXLaEVHZsHLu7Ozqgjoxi79RnGRQvtDKhvIDNk40MFieEIqXdAzbh7bXupZjRfytLgk1CNk1RXOyHFDYzZ8Nh6lngTwQA0O3AzztjSwDjsTYBLUj6DDVv72LDb7Vtb2/PNrb2LYstAItKLmlvvfmW7HWeL7ywlZcvpXxRVkbCpCArFgfs+AjfRRjttvxgaSOlMFZgE6oahVxTzLtSW2w1GwehV21sCYpWPipLuUUYKfdmcGBIxaJrVrBHwPO1bamMkxIxsFD2K1InOGutELJwINQhFjAAT07uJ76VWthp40Sp4YuuiILg0xotInh9tJdik9TPSqV8Sv6IQMKuHAUoIASkSy7fDUxk0WaTHh0ZDnkVrpZAJaDCDC88EAlUCnVvQ+QzKdANyhxiBsCfdt86lj9tKYg9n6ImYAyqHbKil6iQqk4KQj/4Erh96gd9qiT+fYgKlCq0BonJVhCY308KZ0AddYKkYLApfHo7KlCquNowFgU/BGT2AnB6fbAw6iUqAAic6Glb5aSq4gp1BhtSPKhVj4/sYGdLyhkVqBxE8wXZDG1ubPw3QVR0wQRlXp0SFVLrUzwEQIOCsBdQOUNyBKC5lwSKBfDvQlRwz9Wumsu5CgqLp2oM+fVPgVqOcYui0nEqf+aQa2zwteBRykGKA2guRxgtdl1FjZeY4xLboV0VlbKV5Re2s7FlCVmXBRArXN+pC1EAnbvtIL97R8V/DlGBwgW1kNZNBVr+djtWBL809/M5m7s+byPjE/JNpghr1bGEeGY729jAFOR/rznSpnjWSubrfaOmdQHLvbaC4nyV1BgKB1p+RyQjf1uiohe8PS1Ag4VOF8wPti3h90WiohcM670bvXP8/F36fYgKPo4syDIpe/fdd6ReXVtbE4GaTffZWz/7uf3d339sCw8fW3l7y9rtiiUyLIinHRUXfc4fepLniQpeF9V/SZHegIVwRMzVjs1fv2pjpUGBQ4BC2EowTybHJyQMIJB5f3dPBTQ5JXTV4Cn79cNHdtLkABWC73q7SMITVtl/rmPivzRREX81ew4HVELCJycnNPbmLl+ybK7P0qWslasHlku2bTCTFiEzcWnG6olB++SLx5bKFuzS5XmjIdGJiqrWAYIWv/r0N3b/00+sXj1ULkQi0XIyQRpSH9vnrzmC2d5R4U8u5lFo3P0jREXsxPD3dbI4EucCC4KXNkQF7eYcCne3N1UnIVigWwY/e543Ao6VLTzqm8qbSdD1msrYzVfu2N033rA0RD55FDWvN2Sn1nGiolI96iEqhjzEsu12lfv7O7JVEJAiP333RedwCughGw7EKT0HRWqa044KJw8Kgag43D8QUYFyFpKCfzig7e/s2jeffSHFs3VOyfA4r3X/fTMJftDfJzCdqPD7SAWiA3/gx7tkUJhg3YBFf7IiwE7XnLOkIOvf+bka/9zbocD3un8OishOykla9h6BeeEg7vXQ90PDL5r/58kDtw4JoIQUyAkbGx8TUHymowJghsBIgBJZl5zab/J7znZUnHaY9hLabj91NqPie0QF4EzoqICMifuAAzYeaOteDDwev8/qVoGo2N2V6CmqPc8TFW9M37XNjS2rVE7s7r03BMQ1Gm1bWV9VTYAP+d3XX9d6diLL1hGF7a5vbOpcgG0OnRV37ryimou5kkknbHUdq6dx29zcsVYnaasbOzY5MWkvF1/Y2DBrQsv++Gfv2dLCdzY5NWGZ/rwNTE1LpLO37Tawg+MTtrfivucDQ0MCSZdebFizkZRoBcsfACzEYrKLbbm1KUTH2sam6el3AGNrNjo6rLmNnQbgbaV6Ytu7+yIWp2am5a+eSSe17u1tb9urd27Lnx1PcAD/6knDHj9esOPyifZ0zjVYwm7vbmmPnhwbtf6+vN2+Na/A8MO9Pbs0O2PXr1+3sYkx++LTz9R5AvDHYY1sqplLV+zGrdv2+Vf37eC4bLU6YqmcyMyjo8NQe0N60n3tVsKMw9h9Hz3a+XysFy76SbrtJqBVu2WVY84iWFOd2pD5cPFO80J/n0BBVK6opwWyy8Pbs/f8XOTd6OQV+Nrmal0U75z9AOE5t167fsWODg6lKI5kH68dGxuXxa9+Lpz5yOtgUUdMx9hC8MbYJVCaKghFfqt2ZJMD2GldV3cpHWaQAjv7R8ptqLdMpPHQ6IgNDw/Zez/70LLZpPJLDo72pYyHBAPspStHQHeHDjeuiay9Mf33k2cLdv/+AysfcX5I2eDgmGphAFbmMGdbOusFOrf4jCkJ6mAlXBV+opB5amTW68P9PdUK/QSBF4t2cHwiAubnP3vffv4v37fG0Z4l6ZQnw6PetGoZGyjvbOD8i+Xf5PSk/erXH8l3Pl/o1zzSGG8n7N69N+yrB/d1nasbG1attS2VzdqVuTm7ffuW5QGjy4jH6rJP0zMicyKIjgCZj6v7duPGdQetFXbs4ezYGXK259lg68OZi/mjXEeFAHfs+rUbdu3aDZEA+Od/8eWXXUESa6m6zVIJ5d1dunRJ2XfYcrFeRIEd4wPrafZaxhI2cZBX7ImOI2TU1cHnIDB6fGJc91qCQIVpt5R3d/v2be92UQ5JTp9VgkNEo4D1GM9lMgLiEWYWshmB+JzNEQllhZ8kRXgcHx3YIV1a1tF6wRK6vrJhu7sHyvAhoL5y0vR8zsFB2T9hYcP5fW9/X/gA783+7CHRdYHtfIEb6PwfMgV1VvUeT++iCaHujEeAY2UrqEPP7cfksoHt8UBRdnt7WzsimchRrHVa1pDks2M5OmDUHmsicpsKlXY7Wzp1sPPWGsn7iyR0a8Vob+tEheMmIkgrZSsWC3LYGB8nw6OkrYZ7UME2TkJQSCRwioQxr7EJZNwwYOhUwqIMNw1qI1xAokiUrlW6BGQ/l2XNcYtD5XlWIVyxJ3NRaPDoCDa0LqCN3eRytgiB1tr7gquCLMNCILfIl5AtBbbEKYezncSu0dYodIhQNwp3gpztsY6VuDSItiDm/Nzqn4xxqS5FQHF1XbE2OgEXHUJkv9fN8uyg7ZMdF+dN7NMJTEe+mmzR/eMutP19WRscGrbbN2+pqwJng6WVFXUMrm/t4lBr5XpLNSnEnepOlQDe7RJtruJxwgUPLjKONRt1S6y/nTR0N5eLcBvlfYRaTuNG5bsH1vOezH32GgJwGHOQindv37KNlRWNJfI1sKgju2R5bc3aSQgWdI50SDluBMHJegV+w7jnubFPk5HEeEUQofqKvYpsNzo/9/a1XjiB1VJWBa+D0Oc5QIJxLiNXhw5HyGutVWnIlJ/CtC+qi3/63j/xO3CFYMMAYnF4YTJ5eHJoA1PwVmgb49BjKOsbKuS7FkHxcIGqAOWyWG5nXaMnIxtptDViYrmlUWxlSwuYVceAwvY4tKDw9+BmNk2Kugm8sUOo84sXiwo6u3zlimUCObK/tyelCgUmExrFC8GRE5NTKh7xZWRBHhoqKWgTAgCFNBuUrJDICpAiPGAJobVMXnlcV+VEHRrkUOANSosgCxKFmS+eDri79QRKSA/QjiBE7ExRuy2LigBTVyMo+DpsSqdew95S7F6CDkygtuO/FaaU8nvovoveesl1yx5KvyPaOCV0yIek4Pl5doVvOhSMDvI6mw8QQNHUV+hXyzIFqNToJ96CxvN0y5+k2GZCstkgKeh5rrHDptFCYQCT79ZPFCkARxy4SxND/vO6XidUFKwrVZJnVMQDcDx4O/vtIFC0ionKKN/KfJvlNfLppDMidFQAVlFo9BIVOhhnslJV0FHBRgihwUIfg9HExCc92D1+ne+q6N0AIxCv+8nmGJwf+Vm2z4mpSX12PjfFD58HZaPaQkMwYPno0Pa3NlXQMSZ4noBOfC4OSEmRRRd/YR3hUzGEu4YdXV0KnmD8vb/Ta8+Facd7f/594p/j7/C2ebdY8TwP7hfFTU33EE9QvTbYhpwnKi66iqg47oV7zgCbEhuf/m1USkR1CEUkc522SO5p/Fk6l/BppsgGOKAA47DobcMdO2lUVSBCHI2PTQhs57VepEN6VHVQozji5/g+CpxWp24bayu2/nJVz4ZnCwDsZt1qbwrWYRHciWDmWaIigndxLPdaP0mDHdW+IaND9/6cSlgvCSqc+Hr32fSOJHI5er96f6d+b68KPBzgZZ1VLNorr9+TZ72pAyVhnSbew88EmLgvcrRIg4B1JbDWqfqJOlko1BoU/AJkA1FBN1WPXU7vZ4jXdn4MhgGuZxW/zl9H/HPv9+P7+FHm+/dOjyqoa7qqo977oQyS03Xpx8D389chQC3DgS1tb739po2Oo2Z2ED2VyNnVO6/Zl19/a7/667+zg/U1SyRq1ko2LNk5VQH1PjfGevys8ftnP0/o3gl/2TufU5BItOYn2Z983xodLNnN6/PqnNg/PrTnC88VnAo4B8ANgPns6VPNjUEAzk7HHj56YvtHx9ZmX6KHJoCLZ8ekg9s/SlSEzrnT6/vhjoofu+bzv8Ot5dy6YfbSjN27d9empiZtbm7WBoZH7buFx7a1u2HFfNIG0hmbHB+zyctztnucsM+/fmbJTM5m5q5bo9mRlUqjXhUAz167vbZqv/6bv7L97fUzHRXddqYLFrazREXP2A3qxFOiwn3dJPPg3vKMunXI6drv7+czKc4nfHNZ+yYBQhp1293Zlm0SAMYwhGtpwJ48eSyf8GaS9wUAzkjBNj41Y+998KEVBwZlEUHNxyGJQ7d/Fiffy8eH8tBlLCDaoMZCyc2h8/Bg17I5717zrja/Bv4OFR11ZQQH4/1gjXYbPSfT2LuxhqAOQUGPeAbVHmQpwhkOZqh3P/3oY9naYEvS+9Vba7HnxQ6zs+uek0XxKURrPJSa0cKsO2eCV3h3rVHX2lmi4sza/QPkIj8fAc/43t1/q6uCHKnwidRlxkGVui7mcZ12w2k/7365nV7vWnj+UB7rEXWhJZM2MDRo4+Pj9Hnpxxgf7NtS5Aa1ayQq4meMNRcgVLyWWAvF9dRfQ3f0aUYFP9/tqJD9pntCR8tP/WzXdtJr23h9p8QOe35TXv906yk8NHZUqPOaYZy2t+betMePnlixNGTj45P28uWaXZq9ZMtPU6SOAAAgAElEQVQrEBUeNDl/7aoNlvpUm6BKX13fkBUKZMXU1JRtbqwpIBN/fRHM6ZQtPHsiJT0CJLqQll+uS+S0vvJSGRVD/QX74L17trO+rByB8ZkpEbmEaRN0Xd4/0P5dHBzSfAW4R3X5yScPbHf7yC7NXZIKnD3y9bt35WeNSOvTzz5T58Zx2fdNlN+7O3sKMqbr7crlWQcv0llbW9u0VjthYyOjtre3LeIBsoGuhZvXrkmJznmBM0K92banC0vqjiSfxvdSLIeOLc2SYAkbGiwK8L937zXbXNsQeU3rFHv99fkbdlIrW6VyKMIFO6wnC4s2OXvJ1jZ3LJ0ll4J8OLf99VBb7Hgqbo1CfQ7JGM80svTFv97rYNm4SMHNWkKeTtI2sO8qFPz8IYvabDengrMY9p6MNd6HOg/wvXtOwK4nBEfzOQRAhbw/gFlU4L6n+tkTEKhjLT0PhawHP3QOPhBDEVzyeefnY9ZK6gZyAD1wuG05EeBFka/TowNWSrdt/vp1dX6QddQxztMJq0A25PM2PDZq47NTsrNCDFatVewEgLbTUqi61ibOiwTNBuAYsJ2FDGAccItzG0TUixcvbXlpxZ4tLOmsSmkTbZ+gWtVRobB5F/i49bCrkTW/lamFq0JG52KRxQLPCFvftTu3b9mta9fMOP8hAgpZenQXMLfYh/hMgG4LzxZtY3NLlR/rGiAwoDTP9tr16/bX/+lvRcAwx+h4RU29vbmte0DNRZYAFlSMf56NSHBZFDc9e6NNF4fbFrM+0QHDWJB1IQr66EiASI31QmHj/V1LaawMnz55ovM34KHySgDWlQ3hlkcAiADrAN0o14t9fQ4sZnEb8DWNsHrcBLA3gniMts3kpqCM5voRP6GGZ2PCPpmzBGQ8+/LY6IhNTU/b1MSUDZYGukIG9mmui7HAusyzgVCDqGA+c9Zi3kBS4GvP52NsIgKFVGG8QlTmqd+xZmq21FFxdFwRtsKzaHYgY4Z0TuTzQfrQrcSaF10UYvi65yR49l88+4PvNOonlk27G0TsIGENYK6yh/MZ+RzKM9V65vsQmA33gnMWc4zPzs+A7zgp55gDdad+n3JZ3O2C38W9cULS9x1+FozKiTnvSIl23jwbhLCQEwQdUyeBw5Ch2bU3CrZbvM/+wWEQzfZpXWJt9hwdsCnqnD79Lu4z80WdiawjkA8t1qV+kaIeTN+SRVuxSGaMnwtd9BlxJ6/v6H7yus7PKREf0r4evhd4Ib1eot9gDSUb75A9oU6QHttGvTiIFngvXsfc1jmN/A7W6XDm4fOSiyFyJNiRUZvxes/KALdC/OrdGLrJiHZYu1kPMkkbLvXb5OioyG+I843VTavUPL+GLqXh0VHlgxA+/c2jx9ZotQ3EAKIC20DZ1ipb5zTfLdaJF50LuzVx1/XBOz34vl+v207ydSro8FwtYZLB7h1XFcYtYeHqZNFaztpettduXrX9zR2r1arWTqbttddetY3tbVtcWbEWz0pdWzV1TZBJRo1RPjwWfiOHFoW8u20ZYxGnDJ5ffI6My+2dfb1Ge0sT3KKg+pmxxHXgEANWxXxi3Yw4B9eGcPon66czR4Kf/vDP4Q7cyJE9waabtTKMc39JmCaHSh0gw6RXu5WU3/jx4WHph5zoYSiwVe1vviioqFS7I8F8+NcBZPkCwc9CELC2Ec7pC6V7zgpsl/URwTh5BVUz2SkUOPBitbS8vKpgrxvXb6gQISxvfWvTjg8OxegSdgsJMTo8bCMjw2LAAYqkfFBA9InCtPkcLLQKkGrzmbE9angXBO1etFfCxMtj84U9f7GsTU3KAdRg+GGK2PAWei0sQVWOxwbFMveC9xDo4Gh8t0DXBhruo1rUdIgL4cdhcMWWewpKNgrUIvK0FJHE4dJVCwASnjNxuplFNj0eeGsQDyHMMN5vSBb3DPawO7c/OvF7Q6gWQecQOUENILZfRRhgPKSIt17LDqrZ0EKtZ95m4UcJRaHv+RQUA2YQFVg/OVHB9XAfY0cFoaP/1YmK+onUbB62V1Xh53s6m6+P8/gVN/jeP3dfGwuLYOEg8iS0IVJsRqKC+QMrzn2LRAXPn4Lr+ODADne3vc0SMon3Mi9UURReZP0UP8uPERX8/gjuxjl6Cui6DcP5azpfDPSCkPrZ80QFhWT4rKwdzPteT27evwvq9AYe99zf35WoUE4Fh1u6IVSgequ+2qc73vb//7P3ps+RnleW30VuyERi3wpALSjUQrK4iRS1dMua6ZY7Jjpiwl/8wf4XHQ7HRNjhDnfP2DOW1dMxo5FaTZESySJZC/Y9sQO5p+N37nMzX4BFavGMHXIQHWpWFYDMN9/3We5zzrnnMG8JEkUVVzusafNnLjHQq6NlhV7R3j0zMyewzosJ/B/dootnBNihDp1QfOZ6dnF2bOvPXshHVHMccDE6sZKyxlvhZYSZPu0fR1TofdNLXAeFgyBVMEaf2GA91LE5dUxlCaAswJYdw/w5QDUOAPgy31l5aEMAmPIRH5L108vnX9rZSc1mZqf680V8YiJumT6VYfaMtu3u7FhT5Fymo+KPJioGqttrYyru7A2v9rhP/Desn/z3rscjRJEe6uHsvKejQiRoKuR/X6KC+xhEBUU/NkQLSwtq562OjlhleMwevfMd++SzL+3v/uf/zfbXVr+WqMgSfd/8/t9EVLAJ9xJR4Qd6iKzx0REdZM+wzGu5LeLM1LQECajFKLSxreKU93z1pZ1fXgpoYV0Bm80lsDH7PKSIEoP59ZXSTVA1lHl6nQiySwTSH0JUaDybh21i9/T9739Ph4qlO0tWKI7YJy++sNrJrlXY/0+O5Mm+dH/ZLjsl++IlnufDtnj3gTVbnURU1AX+Aeq2Ls/tZ//7v7HttRdmPdYVz6j4fYkKgdJpHPl+H3HO0Ynk8i7t+d9AVLh+MbqT/L/MSy6FQxAHIMby9NSUQJX93V0P5cM6gBqmULRcsWjDI1V7853v2P2Hj1wBKaBmQFTwuZyoIEj13La2tkTaEuLLWsh8V0bFyZEALeqmCN9k7PO94+PTfkZFdj5KmYcfeMqsYM8bTqGYdPFAVGBfEUSF8rjaXREVqH27qIGz+3M4/rrH6NcQFYPwa611KaA8OipuroXXx10KTsmsNdcv4LpdW/Z7QarHmO/P4fBHjsVZ99ufHXWmH66/2pnkr/2HERUseuQe3JqnOy7lx/HMEcS0HRQArHsVUaE9JJH/sT+EnVUAIjczKvgdAF8XHzlRwQDV54pMiv7aETkX0VERpDLTwUOJ3TjNA1ZlMZtqa4iK9+6+Yy9fbNjYODaNhGnXbGpqRiApdenJ8Ym9+fprtr+9pYDg7//wB7a2sanOgp39fQFy2B6tLC/bvXt37OLyXAD/8+df2vLyspTI7Z7Z2vqG1NXPv/xCNnpjIyV749F9y3frNlwu2vj0lOWrVVmGMPbHRkZ1nXQIVbHRq45Y7eDAfvnLT61Z78lqBYAB0HBxaUlnI+yh3Hu+Z/sH++oE5n7hd45CemdnUz/LPJ2empH9LCA9NSzzBQ92rF/o/n6wfE92vcMFtxwam5hUtlCz01PAMfUuAc+o9iGxseycnZ6wzc0NWaTcW7ory7/PyCRaWxXIh5p0dLxib7/7rh2fXdk//epja/Z69mx1S8Kwzc1ddUZxfYDLx2eotXMi57FvUpYhvvNYBguMaqnbhHMnvxNZgoC8jMmrhttdsD64kI4zR08EBUQqU8QVt3QhNC2HXZGsYDxbInorQ30M+CddE6QJSvsran6EVd5VNDc/kwBgP9NqpnXNpqZnZOPB9XJepH7n2XHvEWIxhpz0u5IFV6/reQpzkyM2XS2oowe7Ic6SdLRNTs/Y4r27tnT/vtsqVwGvT7w4ycEuDFkOUgEAHzCR8d4lRNstcTT/UpaRwE86JFodGx3luXbss08/V7A8Z2fAR1kotxvq/OBMnjWxk21tylUDiGRN8DUISzoHpQHoGnTw7O7aaa1mU2PjNjFStdcfPrScOn7oWkD8R52Yk7XJ2vqm5uDVJcHGdJdi+VxQyPWDBw/tww8/tAY2qld16+ZysvGaSuOS9+KZMw8QQR7Wajqj8TkkvMrllb8S3vXcizi/U8NwDnBVOASFKXuAcy7jjnvH2V65Jwn4o87hy/MovD7iDAChtTA/a5OTo9Zueng4N496QJkguSFbWlrQOQKyHryB+V/MYwPtym9sobkn3FvGDKQF68JvfvMb29re1Ljlc6JInxgbs8WFJbldUDcqdNf4vYbybMidYC29uGhYuYzd2aUsqCrlojon52dntWZgKXN4eCBVP+SgLHzadFKMao3hfpxfXApsVdZCcryATHLFvJ/ZAgegFFPOB/WA5qB3kZNPR5cJ6yrz17v43DWDyQlxJcCb/TqdybjnnC3ortLYgpgS6UMnQlHPWXM7nxOeAz4FmQERxe9GLqHsCFMNJXxJtrzka/Ge7uLhLhbMYbekZszMz82m3Ayf8yfHp8KLWI8Q7fLFMyPHCJEH7wt5w7mQvCIAZFnUXV2peyY6TtSppAyRjrpzCOPm83ANjD3du7wTKm5v52QMdZDuNfcs5ZmoVqKOSfmHfaIiFRasocwFEbjkayR7Lrcy9k7KyER1gaoTJIFjyL5dYgg6jNL5NeWe8j3GqQLr6aKn00Rz0Tsu8wUI3sg1Zaz7uXBm0q2e2Eualxd2enRu42NlG6uOqWOQZ0pX70HtSPsjJO3ROZ1zXWuAvakoSxapybaJ942slHi+Uadlz7E6c6SvrBOGPl+yTvOfiUOJi6lEVKTsR+rZQq6otbSURzxNHhHjtm3vvvWGVQsFW1td0xm/iOix01VXCK4dbea2OnhcuAcZh7PL1cWlRD2QHcw95gtzgvEQHSOeIZWXOOri/MrveyK8IHgVxM7dS58R0l+ZJljBF+gqJD9l7Fui4lpB/u1f/n9xB16HmEjA6vTklCYzbZLa+BXCXOoXRGwk4XPJQifPUbUiXarw5PBAMRmWTixueLuyOYkVVR6FkxcsE+Mo3VMRyOtw7naiYTIVoSNiEQ9qh/b0s6f28W+/sJnpUWVQYNXABrK6tmZHJ7T5dqVCgJxgQUANtDB/K3miu50VYDsTGeaUVlPems3aFzEHNVlEpS6Ryr1tz589s48+/sQu6w0rDbvKzW002IjYVIPBTl56sr5xvys2i374T1LlRAC5bGrE3Lt6gbYyKlAP+7m+2HJtIXWRWicBnsqqEDjrpII2Z1k0+SYF4OBfTl+oTCJQURumAxq8v3dUeIskG6tyLZISitbayMZQK7y6T8i6QL0xovtI0cyL6ZDbw74JUoL2QdQZKEwoDNmEORi0bXRu4hpREQpsB3ndxz4O8f/FOyqmp9Sij6IAlaiUK/V6v0jNEhU3QbX+AeZGULQ2yNTdILdIwMACQbrzfp/bEBUw7DnZD/BfFc1XKGCOlVGBYio6KnopxPJwfz/5c7566fkmoiLr1Z3d4FUICShwADq+FwVqkBrZv8ef+0RFNkzbTMWfuq2SwqX/8zEaM3kaNz/JH0pUBNHHfWUNUf5IUmUCprlyrqlimEMWoADF/97eQfLbBlgr2th4VRk0kKJqs+74AYX5KABDQXBtWeKlKeUHW6xHui1be/7SLk/PElGRgrkAZZJyRippWai8Okw7W2wxT7+uo0LP5w8gKrIZFczT8Me/+Uyyzz37rPnsDx49srHpmdRNAahKh0fXXjz7ws7P8Nh01ZrGTwI1IZm9Qw6QoGv7e3sCgf6zdFTcwIRvEi5ZIPTmuL0Wpp0JYMuOQw+gvm61Aoj5+xIV10Do1K0GIc//3njyhqwQOPgD2lQr4/b6d963Dz/+xP71//K3drC+ZjbUsG6OYMJsOHNaR2500cR1Z4kLL8QHlNRAmTxk+V7qeMn11PXnSignK7QVR0i5BoRZMTKVaAVHXQgJ7b5b5ruMg8FBVNw8NDgZdJ2puDbWv9JRMXgS/TBtbRDXA8xvjteb7+GX39H+OD09aSsPVlyxuLRouXzFjlEkjhZtbLho28+eySZudmnRSqOzdtXOW3F4xOaX7lmj1bW1ly+tpUDIsoCJ0lDP/tPf/8w++fifrNfm8MBY4flkacDrK9uAFHbFeH+MKM9o0GXl3ZQRMMy99Y6Km19al2Us4skWen8OoYwP7cE8J9Yv37NRQ0voEPWA9qiCFSsVu7fywF5/8rZVx8f0/AkOBHjzwz4qTCe+eJaXl2e2s7vrgcUTk6oBmPoc1E+ODwXQREcFB3p+R987ORGJHB0VMS8FJDWbei91VJC5xdxAiXh0bLWjmixrSpWSOmcVcGhD9quf/0JrinX/vyUqvvJcboRpX19Xrnc0ZokKzcQMUeFtNB4E7GBhPIObHUrXbaFiv87Oh2xHBSMFooKOAKyfZE2SvL0h2oOooG6J2ovPEPZ8IeKIrq7s2uLKQCx7BjlWfN87Kq4TFdhbSSSg8eudFBL8pM7X63WHh2mjDFYDJ+SowBxX3guQTkTFxx996kGdk7NWO6jZ3bvLIlVPCa3s9mzp1pzVL87s/PTUFpcWZQ+D1Rm2J9TOx7Wafeftt60yUpKFytzcjL348pnAIDqRyHGhC2N+bt6effHUFudmbKxSsqX5aREVU7NTVh6t2t7hvi3evmOlSsVefvFcdjoTM9Oywjk6PRZ4/OLlru3tngrwkif/2ZkU1UwawPNf/PJDe/vtJ7a/v+/AXKHU76j47W8/sSdvPta/lYdH7LPPniqPgDm5ubWhvYUMi/2dHeUtsFJMT4xLEbu+tW3rBHVjGyVRDl0IZdvd2ZIfN3v29z94Tx7yL54/t8P9A7u9dNfe+877ej7/+t/8a1nA9YY6ut6lpbs2PXfLSpWq/Z8/+/fWJV9nqKAOdNaJsdFRI163UPJAWwhOCBNqKYB+VMbqRji/kKqXWpSOPolLEqkLiIvdCmBN+HtzTnDwzAFc6mXOfsf4gUtX4ECdSLTU6QsYHt1/jGsB3oKPHYwtFHMigx4+WpEdMfOF6wS8JECbM4IrsNtas/gf4CD7DKpqLICYT5VK0cZGq7KXQaA1PlKwy9N9dUMs3b4jpff8wqIyGfi8PbIjikXb3IVAIoiX6+rqXIgVDuvD8EhZKmeUvhACUkMnm9lLZXVgFVa0crkqUm24VBHgNTk1pS5iQEFqYfJKRLawQ6Y1RkR0nBSTjY66XVN2ZHjSI4ijtm9cXtre5pY9efyaba9t2MzUpN2/e9euyCOgA4D9kjwWupCa2CBdSsGv8O/NLdXCM7Oztn9waDt7e8rHojanvqgdnegeY5syOT7hin46//N5gddUHcx7f17JEaLb1XOT4Kvh4K832DvJwRfkBDalqOA5g4FVsEfxLPmi+4h5x2s46OwgpsDjbldiDrqZOMOWAZkJQD89t+OjY53hZ2enbKRaluc+QhQ6Uln7NjcRVk5qlDH+9g8PNQekeLchqx0fi6hhzWUe8iTU/ZxM8yPQm856rhsHiH/53/xLu7i6sP/j3/7UbZmKLnBU+LlyNnsKYb99e9FmZ+ZUo3M/9vd2bX//QKpvhfFyRiKbZHRMa+TGxpbt7e9p36fri+4K5pA6qwlqV3i1Cy/JiGB8cFYlFJl8HzJuuFeQMLwezyEAfAgsWbSVS6pZOPtynza3tnQmg4iDVHIbZDoi/HelEhe57fUO91odVSkr0CEkn+PMU8cy2upwUEeFsjLYTz1/FIJnYhyyflbdbVEjASYLXyEgvUyAMTZP5O/sCVw+OjqxAvaVZbKMWKu8nmF8MbdUH2PJFpZNKR8Roh5QmjEfLiRgUNzDIFRkN5XEGlL+pw5WnpnXet4REEJXDdgkeo0Mh7ATF74GgYRRb8KAokMjXCgkNJWtundVOyFibuWZOmL4L8+M/4JVxVzodzz2hkQe8RoQ4XQfAubPTE7aW2+8Zie1A3XeP3u6aqPVgtVbZvle1x48vC+SHUISAnV7f89++/S5yNgO958OE1JkIZh0pvR6IntmDaus7FmL7+se9QWjXjfFvwVJEzkyXm868SYCTbULGCWdlNhY8Xlww4UookZt2vLinE2NVvXcGQO101Pr5vK2tVezYglSzfNZ6A5hLjOuwUPonNLYosah86k62r/3dEJF2LucS8ojdn52maysS+q6cDs+cM6w14fIKEkEglUg6zr40fTM9LdExVePS9/+y5/6Hfjze/elkHFQzn3+1EaXADa1BqJmoFigMFCQtjPmrup373Y6FVjM2MRYtL1Nt22HB7s2XM7Zm28+0a3yEK+2Wv1QpTC5KDrYGNmctEkR8VDIq7hZW92wZ8++UFsrHqlcGwX99vaOHdbwREaBMSJCZJTWKIgQshxKJVu5vywVRng5yYrAhuz04kybs7wNOagJzGzr31hI+DNKkGfPntvu3q6XbylYF0addjAONaFgYXNUdwhkSwilAe7xjU7gPotTbGCuLBvSpizVAEx4qWDYJbmiYIBMhFIAz9o47PmCDHjjvr4ReBQbtzaSFIbUJy2SDRSbJcUs9z5Yeh2E06apeyJlhZMeKhiSXyGfx62lPCCPz8/P8n1AOIpLDozePUGnx5CAXP5MsU6BAHMt66fUkshhlQOqM/VyU/xKRkX/wJw2IcaL7kFSfGjPDkBMJ5SuNge1LhYJ0656QY9SRqoi993muWNtQgg49y6ICp5J/z1f0VEx2AgHFixZtbOe742MCtRitLk6e9/R4ZkxQbHGxsn7E2yOSvT89NhtkwDJ8fQmrPTiwna3twU4fd3XTaIifk6FjguNvCBJXU9SJMkr3dVPg68oCq6rQ+N3dbALcA3VV7JK0+tia3XpYWahWggFwM3r8fJy8P/djsMBsSygngVdHDML346hftukt6+ziQOc+bjkvuqauh0VVBxqORCx1pyenGl+chgDKBifHBfA4YFxEcLo3Rma83inV0b6QYx+TXxwXqNju1vbdrh30Ccq+gtB35YjWVok0G/wsf3B3CQqBECGvVN65H0cy3+h/yz7xatbuKZCLf03KdN9XXVyUvf2FeBnf2T5QFGxjJLojTef2BDjkPZ+gfgA21178eKZnZ+eSMHpYACqJQKbGf8OxuaMYpNgxBMd/N0jL1Tg8pAbiFsyi2e2ML1JRCRY1jt6kq1Y9uP458uOILdW0YEz7NBU/LtdWf8r751d/Lq60zLrsNKHkq+91pvs76Uzg79SIqrTHJEIoOAHXsbS60/ecMKykNeeOjU9b/cevmb/8ee/sH/46c/saHdHAcHdoY5DnunyRDSnvUHX1U+vD7XnQCEk0CFz7RwcY5Y5+QH47cQ1h5mYTjrw6GU8X8rFCF7oC0yPAPO0fgRJIQI8ZS/4mTFmdeq6+spgi0HqN+46yZB5Hr6oO5eSPv9gjKZW8/Tw9O8ZQsSvDeu8vNb1u/fuSqSAZ/pQoWr1TsvKqIKHi3Z5cmyXZ+cKEu8UyjZUqNjs3IIC5MFD19fXdGBjLSZgr1LI25effWL/8NN/a636hTIqJLdV+PnXrM+pgywAobglPKdsR8VgHXbluG6BD+cM+ZTW8ET7+S33ekz3UkIQD1D0fclzasLLV3NBe3bJ5m4t2sPHb9jM/Lw83jXvtbd2pagMwCY+FtYmdNhwSB8bHVftxbgE9CCjAmUX4KTbZLmK0ImKY/0dACBUb3xuDovUEwqu1fV2lQMCKMKaoY4Kcrsq2H04SFDM5e2jDz+y7fV1632d9ZM2qeio8LU0u/9kdx59XmVUDKyfAuTyYXXjmYavXprvg5VW2tnMPvo1f+yv3f5MuTbWpQFRgYuCr/EOlnmnQfwvs7JrBIS/tI8DX8Nif4o9hFqDWohPMjFFqPy8dTrepasw7aSYZI9wRaxnVMRnj24Qt35y8Mo7FhGX+PynPk1Lb39vElFxdiZbkgBGWCo8MDwRFbFeJZJ7YNcw2MtyuZ4d4ZefOioccHHAMoiKHzz8rp0cnSuDjJBoQDWmJb79KBsZq3NTkwrIRhUNKbOzd6hsgP2Do34Y8rtvv6WxjCDn4cMV5d1hP0PdeHh8ats7e7JJWX3+zKYnqjY5NmKvrdy1Th3f+p7de7hil3QnY/HR6ggkJqOFTIEK3ZgFFKVH9tOf/ko2Pffu3bW9/QM9bsKFsVNFvbu2vm5LS0sCOpkzrGN7O3u2dHtBe+/j1x7pM9I9srW1q/MAz5Xng0joYH/XyoWC3VlasOPDQ/n+M08RXT1bXZcv/XBlxI5PjmyYDKUh8+yOqXE7Pjq0R48f2IOVZXv+5Qv75LefqTvlrSdv2ejEqK2tvbTNrXXvPC+V7eTs3O4/fGhHp+e2t18TiMkz7rQ8iBoFMV3LCAUAeBFEQdYcHhFw6zkSgLCsGxAWCgWVQrggpa3bi3gINM+UjmRZSqH8T3l5nGHppke1imIfwQnjVfYZlZGUj8Fazfhjr+smAM7nluaCLIebNjs37aHWCIoEMGKzUbXZmVk7Pj7S696+vaRrdbDRswYgEAC0qIM5R+Z6ZEn0bGqybA9XlgRYPnz02KZnb6nz4cuXL21ielaqXDIaHr3+mjUJ7gZQtY7RBV+uVqyFdWenJc906iu6Nfo2M9jM6l6RvXFklfKIslkAi1GUx97MfaY7aHx8VHUwIDQKZt9fYyP1fUdnWd9UdT6TSEtrBVairE8de/Hsmd2ev2VTo+P2/PMv7K03nli5WNQ94AwGoE7HAs+W8w+gL/UFXYpn52fqsvv1x7/RHnN0cizwmHM/ACUODzs7O74OotgfG/PuBc6tKauB8cGewOfgmXH/6TLR+TSf74PfbnHlOZdRG1Hn83OMXycm3CbZu/sAit1pQeHj1LzJ/oWsitOTY7u7tGTtllsxY2/FmXFictyGhwsiKlg7wCM4CxEmfXbekniSGoT1CtLt4vJKawNd3scoz6/OFewMLkBtqM9ClwTBxBDWUgO6Wv8v/+on1h7q2r/7d0EtUg0AACAASURBVP9WYeOspXQXVSC4ekMSYqXlWFZDeOIvLszrjIN9Gfs4QCtnG7AO7stwmfBtH8f7hzXDEksBySIvuxlrNt9MeUZ0xwhAlYCTLoOy5oMwnhHOS3jnUwcMiaTUMysQ8F232dkZXTNzLDoh+CzCNBCK0mWV8zMcz1fWXIzZpt+fAPkdt2IfcmcHfl+ZqdhGYanNvcPeqo2g0kOnl5YWNQ/o9OZnlTWRLMM8cN7JCizseH7CiJruDMIX5BtriudJdCR0Yb3RmSfnmTncS/6snFGcPCBTsbbE/QKSFewkBbOLgEuTkHsWczaLB2k/jjN8qjSFHSjkmhyekrpSuF8Q27ymn3G9HgjS1vMqvGtIwhi9rh/ivQstiW/7ls2OzYAF8RouDvQ8Vn3GIbd3rFacDLu7MKd9o91o2PnxkbA4SMvt7S07OTlXJxlZpaz1iCaoM9e2DyxfylmzS9d7NzkScMzxnNXAV6ImCbIkW5v5mWdAaEQ3GM8rOjL4c4gbNW5ShoW6SXoIkJ2oYF6Xi/7MIGFYi7vthj15vGLzk+Mi149PzqxUGVH9sHd46JbIEL9FXzvBFcArsaRXPd72zClE1uzbZ6enWifA4yYmJ1T7glvJTr7rxDnj8uT0xCYnpvrdN8oOOj1VUDd5Mlj2CvMQqZj/lqj43RX4tz/xp3YHXlOrMBNl0u7cvq02RFrZvO2YgT8klQ6bCkA0C0S96e2YsitCzULrnUJtvAOjUXeVGyHF7faV3bl7y77/vQ/EKqooTdkVvil6F4Ev4IQcF+ywdmLPnr+wrc0tHUxps2bCoywilFXB2hxS8gWbwMplblpKBnwjBZzTOljIWwUyQpYw7r3JhsTGJzAvhVNT0LL4u/ovJ7XU8+cv7eDg0IGs2DzUeQCo3hHbSlEtICct6vIrVXA2y5UDNLKjyYQZxmGP+8aBUKCACmQsksiPAGD1Q6AXVH4A9J9xb1YOIVJGKnTRrWk4rEH8hLqtv5irFQ/QwvM4KB4oYtQSKXLF21/FMLPRJ3ZZi386AJA9wS2Ia3cfTw4esM1dP4DIW5KQbShziloPxWYDw/aJbgrej82Jv4/Pe1tlbIr8WZ6gCahQUZyxWPENZdCkzPXe/Dd/Vj1T6C1ExfmlNu18qSi/wADu+OxqoydMu1RUAQdpIKUH5Fm7rc0iCoJuSi4WSJ+Kg3ju/JtvDg64BJAvooLckYxdA+8LUSElcqcjtUmumFeLKWOEFmcyNfB/lVotHQpcIYuS9VLKth7IWZwpMvYh+nx9MOyr4aHyI/8KWBOQxw2YN1kyBGh2DbBNYzaICoglKR4SWAlJKKJCinQHx7Kg83WwaECc/L7rZsJR9ZpZ9SVzQMFzAiiaWnsopXg+hBo6oOL2UHypawj1LkVUZcSqY+M+l7U2ocpxyw3UO7IJSJZsofrtX+8Q88gtoY7SmqG7GTk3mQ82uI+DYsq/7Sr3eBoJfr92SwZPyEHmCLLTa6bgSYXqohpKYbvxPV1OmuuhTlHbdoY0ELCbBDs+rLzom5metcXbi9aUvU1CTLVed6Ro9kKu2M/X0adJdgFaEztNzUd8mb2t3hU8Xnim90mdA64md6ZgQKYMxk/2hniHkCshB//31VEUAGWsXxxqff4OVO3xW12KVL9ZYaCnb/nz9O6D5FySbPYG76cug/SzIvE1PhNAmgdMJJi1aLNzc/L255CHOmtsak57L/va9saG5j9hlTpspzZr3RO1owVBxZWgnudG+oFh8CgTOZBBZvtrZ5A3fZLDr8tHYDzbCHuOMcpbp+wbZVQNQNDsgpJpyLr+EHTJQZwkUiW7bvku2wf4Q/2UHkPaf9PvXUNUujYk8jsprPugqq/S2uPl9Y+6dcRuLSzKrkiPcbis/V/doWp6aosAVm2Dsr9n9v4HH9jyygP9eWNzwy4usVjAk7pkpVxOdm//67/6n9T9xvthe+Gfw/f/xHcN7kXqVPF9Jc10PQ+tnD629GGut6XHQuJrx6BDUl0/ygPw5+cA9WDfzILM+l7c0DjoDtPRM2nvvPtdm5mZ1+GKzwdQl0qZVBs4CRlfWMkcHByoHuN+hgKPuQ2AA1FRLo+kMG3yLQAoLgWGQmjK0kV1lB8GuU78tvG3jgMzzwGiArWYwrTzhJVWPDA0BXm+fLFmX372mbWbF6/iXHW5X9d5NljdgkhzX2x/bn4/pUiMcfr19JPXBBKFuCf1dXr0xnp0w+4w6gWB/v139t9xIUogiKz3LoRR4HTqmArFs3baPnF6kyjzdUvWLQqoNLu1tCggo9ceCBGippJlY7JZyHZLDDoq6oY9ZygVvf7xNdprgkHtobo1ZVSEaEDXkkJYA2yI++C/m/WV1pNwEtxMYbX9DmX2b7qGAanTZ/vR6z+UYntubsGurhoCgjmL7OztioSj/n/twYpNjFfVKcZ77e7X9L8eljkN7Gcu7cHKfeU7ABpCTH780cf25MnrAlQAqNY3t21ubt5qvG4pL6Liwb1F61ydqHtwamHeRifGZVcGWHR1cWXjk1Oy7BH4SbD30Yl9+tlLK5bGpPSmWwRgA/U7YNjFFSKtNVed7+/LMoMaHYEFHWKbm6t2585tgf10L2xt7gqUm5mesc3NdRufGFVHRLtxZQ/vr9j2xpo9ef0N3UMyKsgYurV0x07OzqRcv7w4s9GRsshBVOfjYyO2D9ExXLW333pdIbwvX67LxgLVJraF9x8sCzBfX93wjI87d+z4hA6Vkr18vmpj1XGNCT4znv3qKiwSLFyS5QxzhY52uie8i7Frq+vr2htVUyeFMdk01GtxXuDsw8/KBg6AXl7pvE/TxkfH9NqMJQc86Trw/S2EXJyD+N0A8AQatto6LzDP+C/3RJZQyk5MocLliqwQcRzguXKWRcgnAlv2KDmB0fixj5SHFbgKIcYYmp2dsNffWJGgD+FUvgRA27CdvQOdPx68/sSer67KPmSSXChEbri158xakIZeYKfuR9M5QIHL2E7ROZdsWFl/CZNnawAEp1uDX93Z2hSgeXFxpvWWMVQolW10AmshMgQcfGQssvRojU7rXuzf2oGGPMi7Wq5Y/eLSVl+8sHfefNMa55f24osv7c+//0Nrkg9ITt3VlUBe6hNEb1q3hpxAQlTkpEVLQNwnn35ijx8/sk8/faouC9VHEDDJRgdBI/armk/MS4J7OQemHZc9hteCyJGnP+MDx4IUJMxSKh9+hVr31AlI5wXXwrMDi0C57B1jAwEUK5DO+pAj+ZwtLs7b3u6OTYxNuF1RvSXLJVbZqalxBYhXKiV1gPABGcMECPP+3jnYFUnHHCc3amNzU+OhR87AUE9jq3Z4qDEoQLlLV6uTQ51Wx0aGR0QmEoAtYLfVlF0RBARg8P7+nm2sb0hlXa+jsiaYnhqnJbso1pi52VnZ33L2hRRBOAfewfmda+T8y+s1WoRHNxXqzV6ceCuJbOQkgUVb2Tse3O7IBTSMIYjKcwiITk/PHoLRSQjHO8BRsB/EggkxKPcyspbifCDnComeXNSpLgqEqLKjdlKAMeK2vlH/eL5F/IyspxCRYscGIVFEIDRsK/fv635sbKyLEBsfm7DTM6yfplWrcE85r7OfYN3EXIKMhQzgPtQb5LCQd1jWeZHf9e4cn5dcE9ZwfBb2FMRxjF2+vGtsULNxvXTasD45loB4yIWVUUcGvhG1Xr8rTPbcSeCBVTE4RLJpZwzxJUIzdQ15cZP21ZT1o+/3/Lyu32dNTR1LqolE4Pre7nWAY39aJ9ibCznNDQioaqVsi/Mz6qTg3Mc6hc0yRGO5hJAN8RvzuG6n51faY0GoDo/PVXs3KGkhimS77ELfOOcHJhQiiah5o8oKoiJIDScqvM7nezftoKMkFg7Zw97J81q97AM/rAjbYlg3lb9i9uZrD+zW9IT2yS++XLUydQXkWburudJOZzTWGeW0pXEPjsA9haCErKbDCqEE4gvuLTgm3+d+sJexTnAdEn6fnWkNYY3jM6l77+xc6wciEK5ZdXuIkgoLP7hZBd6oRL/967d34E/rDsxIdeTAd6PJIucFpAA+NsikLvW1DZA7LzULiy0gOBtAALbMLCYnm4p7xmPHMmS35ift+z/4ngOITbwZyyoYsBfQkpCCzihAfvvbT21v/1B+6O++87YmISHCGxsbzqaLqS6pC4T2MXVyVAqWL/RURLJ5VmjblJ0FxdqwbW9tJkA4J0D/nMAvmnBzORsdo8WYluKm/ezf/4PVjk6lHFCoU1KS8nNsMlw3G76TEyzo3DNvW3ZCwluRvcMhFNSu5qXwYnFngY57Q2EVrLpCiVBCsjkTcicPX2/npBjRhiCsqqMMD9RhFAtct4gWfBnZ4MIbX62ZWK94+Lk2tgQOxCakBb/jwWo8My146RCgzUEe2V5MxgapelmAniu02YBR/wNMi9nXpgDxQj4HqqK6iArPqWAz7Cqjwp+7s/d8/ZckKnjmcRj2osmVDkEeQBrwfDnwMm688Ekq99RREWBNgEHcwzi8x4Gc8dk/sKd7FJurvP5nZ/W6FANqix0u6mCqzw/DfnRsZ0dH1mhf+QatboCedVOLOZtjt+ltytmvPpD0xxIVWblp8sf21x+Ec2eLAT7vK4kKHQYpdK+SImzQKZAFu/r3NkCz7Pv/juWzb2GWVKBZciivw4t7m3Iduh0iDt3Hm4BcqVXC3iZDdkQRxtsLfAnFvUD1pBxNh52sigOrMqxfmEfqXpJ9XMIP9YcsCZT9cNE55YSA273ozgzG3tfdC4gKQNZMV4V7sHowWH+u9oFpJw89r8MJgiCHYzw7kQEJqlumL37GvaLz1jEvYHV9CcjXz8sHFf/iAejFuuHFJYcrbNSchMySjXEd/ddUQZwA92vjItTQg9LL8Ts+fwLYg1ZJP5LNs43P6updKFu/BzF3s7fYIb0w03lFtkIi5MQPpP0lDhPRbTA4aKSuI0gyyCy1plNkcjAelqUh/6tOzujgCOhLoXx8VLOd7S3b2dqSVZYTvOm4klF2Q/oORpa3FEcXTvAa8dlivPbXpj5RMVCLxzySJ3Cyk+h3q6Q36iYiKZ5ldh4kuPzVI/bGFOgTaTGW+iT09R8UCJEJCk78f39wDmErlvmVOKA4MB+gJwF2JbVO6x4zvgvsaw4pcyu0busQlrMLFLjdnn3n/fft0YNH8pzd3t2zS3KbaPsvDdswYHypaP/qf/wf7LR2qA4GcSiJJHSiLV1mssXTPU1AeHQ2SImuNTZLLmXvgRr+k0rdiYqYLzwnrLv4fnZtjXsQ+2msddn1Wx0VwwVbvv/Q3nv/B9ZuY2FH7QZRkbynk0qRQ2hm2MlrF+CUAzpgtzIqul2pIkVU4CediIoI4lZHxemxFYvebSEQTMA6h17227o1Gxd9BT+fB6KCjtrDgz15HwPuoNzmGQAIHB7W7Nf/+CtrNc6/gajw2eljO5FBET0eczkzgL6OqPgdW5Jq2cjrurY3+Eo8+PVXxFfEnMwKCbKEk14v7WH+s9RMbr0BQC3hwzWi4vqKRg3GlzyTE6BP3Yy1TBAVIgIEQHjtw3/jUB97SYwjdVQMBVHha3qWcIl73f9cfzBRMRAgZIkSiAVA9liTJBhIRIU6eotF+8Gj71qnDSlTskLeM/b29w916D+/OpeN2J//4HtWHca7HYDsQGceetd2tvc9uLnXsaVbCxLVnJ4e2+T4uK2vrdrtO7d1VmAtgLSkdtzBYqlcslszkzY7XrVha9j4xJhNzM8KTEUJj9AqXx6xtc+/sLlbCwK8pLC+rNv/9bNfWO3owp48cXsnrvfh48cCqQlr3dzaFmCGbRqvUyoAaF1pnqKIxs6Fda1+1ZTVD4pNCBSIhsOjA+9m7HRsfm5GsemclTjrYEvx6efPZP0ke43ckI2PVay2v+sK4VbD3nv/XTs/P7HtrS3Zwrz15juWLwzbJ588dQA1B6Bft8ePH1p1eMTWNjYUgkw3C8pjAD2U4Dwvzm61k2O7tXTLjk5Pbbg8mhTR7okfpCr2MWQQoDo/PjqxUWyTkv0MNcVodVTEAEuHRHJJ7S2P+iQm4byDwp3xx1mLcxfnF2ozt6J0r3MXbmFL6/a5gEYKwy04eTx3a1bjTWcwQM42QC+++AV1A1DvOEAIedXQqgLIVC7xWl0r5YdsuJiTVdBbT96w5eXbNpTzLgOU9LWTE7uzvCLii/xDiLJHT96wX/7TP9n07Jw6fFtt5CFtWTQxvq+adZ0zhxkHFxcS3dG1ztqjLgyIe+UIXemZ8VnPTs5sffWlViHW55lpbJX5WV6V5p6iQERyXeiuUW4FwhH81qlpWT/ZE9I6yXuy4ADOYrWMHW1tb8/efesde/H5lzZaHrEK1kDKKaPjiX5aXo57izijCA3g3Zk5OkBO1Dn09POntrJy3x4+fGgvXqzKGgwlMuA8Z2J+VpZDwil8/mkNY99Wpx7qfeas2+zIxrhScRFeqj35L89YuwIdL6nrGxCeDinAPxTODoR6RROdMhKaFOmAn1TXu+piy9vlRcOV8j3yUsqyPSan6fbCot4LoP7i4tztZLGPGndLM+YdwCO5OW+88UQdjsfndHYdWKGUF76BahuCpnZ4pPmEuhyiqHHVFP7S6eFMwXm2pBwuMjtRWoN3sC9jO3N0VNM93tzc1Fjliz2e12csLdxaUF7J66+9rp9hTKP0Zu5ccZ0dupTGRbhA8DGGWL8QazqWM6zxV7+su9WQ8nEuVTNAWLL2ugg02RzJUtvt15jnxRI2TZ5RxVeIX0XKK6vUhU08W+9Ecbwj9hkwJg/TLntOJngG8znNdzAmCVU5u9EVVcYqr2T37y9bqVCwvb1d+/TpF/Zw5b5cOsjM2NvfEQlM99RR7VhkEusv89YFbAhfsXIF5/Fr9nW54mRowe3Qqe9ZW9UNEvkUyu3w4GrGMAI3kaYpD8L33cgq9YIhSNsoxPx85XWFOtpSJofmGfNWNmngN16H8prxOlrvwJfUQUn97O/BWgMh7GC6g+p8FkS/PHudh3s8S37X6w4Jc5VX6sH1Swu37LvvvWW/+ehDG6uQRXRpw1iT54taMyHn290hm54sqztwaem2latVW11dt998/lxrb5Nyh3NGslgv9K3VU0d8IqpukhdR9YQ1e3xeiUaTlW8QMD4W3bmDvSqICgWqi6jwWlul99CQjVbKdnV1bqPVYbs1PW5Lc9Pai45OTu347MJOzy7s8OhYa3ih5NZ4jFuIKtaVcGRgnMqW7wQLMfIniiLFGAcTOD0M+/6uzs3DWhIOkU+DvZNbP/F5mO8Q6CLwmi11VrBuMc68Y/xbouJ31ezffv9P7A5MBqgodbiDo3ypyEjFmFRLEZjcxRcSyyQH/BS4o9Ao3wyYLALqE1oyOVa1hVtzKmgppDlUsKng58nP45XIpGbDJg8CkOA1fLwXFuzzp0+lcmCCxiKJXyjesnR5UHjzet1e08bGvZsC4KFKwNElgV4eaENB4Ep6D50qsDEkW4Ljk1P78svn6uCgMBNTn7yfs+dMlnxX9aQ2eeyRxD4H5+0e7WwAyljQXwc2O1GMO7HD4u+gZl/Bx48LyPIcDJeKdJWrgf2G9oUum8yQCgupjvI5kUYUu3Q4sHFKQUBorNQjFGUOaure8LdEDrFxcnhFyc/PueLX7xeLM+8L6tmmg0R2UE4SAfSjyHHvQw/WFriB+rxR1+vA7sq7nx4R8knS//gMrVbDJhZmUsH0/z5RIeuI5LEpomp01PB3jc3cN38HZR1c8mIkDuMBIjCeQoUYh/wIwwovlWxHBcAOfrxeFLQV3IydxfjkpOYaANDuxqa1aAHNeZeCxgf/SzZsFKFthf4NvuIAIXAuYSJ90DEDwnxjR8V/JqKCa0aBwCFdHQWZ67m5LGavOwu0/a7lU4WruqnCu9sLLRVQHERRRV/hIQwVyZxBlUOnU0dBfbL4SDY1IVfRvNCB/bplThTDPB8Rkz3WgNY1KxCBkxwAwuczqWD7AHYGp7r+OaOjQKMrERWJCFCV9fV3ImJqQn3qigq/H/gDO5jj64+v54moSPYiPoad9IywcZRrTrZ49wnrsJvA+FcWXNaalUXDMwfZ62oWDqlhAeY3gvsY7+9rZ3xx8E9+qX1EOoHJryB7vCXaiQqBCQK9HRfsZG4j/xYdDro2MP2UA6TrSApq3/NSH8mrciD6RJKD2wFy6/f6AbG+3msfTSoeBdjnnNROV6tDC+sQFg3VyWmt53hr86MAEIQfooxDZYtVnh/i/F7EvYtDp/8j45b9NzvYrhM7/Q6c6PLIfO7B+pbl1bKWM04guUeujwXGimcn+Vf61qsHbYYY8fs88LDX62XiQBwUH1w7Fljx9ZX5Q6t2f7x7R9mg08j3Mp9I/lwK+Mey95KDlCaohlZYanm/otSRdLlgqcK6eXFxlfYEVxLyiqjx1smuqF+pWmDDB99JzfnXPgNv4fo4n+vpQfqewpqEj3JS2IlwSuSMq0XZz+N++aHLxwIqfJzfB0Cxr1P+TOK/IQTge7G+MSbL41V7/4Mf2IOVx3Zw6J7ulZHh/p6m14LUTT7G8QyyRAV7ZxAVqAaxd7pGVBQ5gLv10+npkUCJICq8Y9efCzVB/YoMASc+eW9el9/D+kkga6WciAq/RoCUX/z8P1n9HPD61V/f1FER3QqxV958hWxHxde8vP6Z6w3LU8CJrCXczdf2sTH4uvZMEtAa3406Q0QF3R6JLeIQ7VYangPA+PkmooL6jDGumgfV43DJbt+948Bjx0UicYBnzARoFERXfD/EGBy2sToDIM2Sz1Evube226VEaDx1S+SVeEeFfy8rGPC5ne3MiLXOxz6AhyxKYr1JYyXbUfHjN//caofHsleojozbwT7WsAWp/RlEvMWdxUUbJe+Ejuty1Xb3Du3g6EQWTKzHtdqBPX74UN0Ei4TjAlLQISqwNK/uC0JACaw93N+zcjFnY+WivfPksXUvT7Rezy7OKaeiWyrawfaWTQICj1Tt/PhMQHB1asp2tnfso4+/sMmpBZ1PqK0BJpfu3HHLoHxeACMfWB0V426XyjlJliV72zY3O6N9hIyKTcKxGy1bWXlgT59+avPzM65wbjdkU7O/u2uPHz1SqDG2WB//9qlNzc7aCV3u5aJVATzzZj/+8Z/b1dWF/PjJPOA1AEpPTy9tcmpWJBnB5CizL68uPCsBqwqASfIL2h2bGJu0i/NzAdrYr3LOoKvl5fpLG8WLvjOUrJuGZWtFtz4WkwB7sSfv7+3bs+fPpVCF+OSM43Y9ZPnlVD/TGc0aVcInHqEFSu5hOmHITHQLTxdv5CWqYm8QkAmwl/ztY83kXMZ4bLZcSIa9lgDber1P8ADYMrZYk6iTAIgmxkf1jJRtgfJ6uGitBucjs5Xle/b2W29Zt9206uioHZ8e2W9//ZE9f/FSnTI//hd/bdVy2Q6Oju3pF8/srXfftatm21Y31u3+gxVrdOpWbzdtqOh5Qlg/CXhvuVhNNSfAfcstbgNgZKxyfttc37CzoxMPtu52bWpyXOAhtQnuA1xvp9ESCDZ365ZdAICXR6yHEpksQtaDbluh1wgGdC+xRm5wHRAOnim5t71jo5URu3/nnn38jx/a45UHNjk2ZjxDzp1XDUR+Fd17niPgL+TR3v6+gHWAbbp0Hj1+KIu2j379G7u8YGxxhicj08VHdB6wz1xcXQln0JkaVXgi4MIqhT2PdQzlNnOLPwMGs59AYtABTF4dBDNjAQyB9z2qHencLPJMWZoAswCDRQVdj1VHbHSsIgKF3BX0CRcXdWtBdna4T3S4XIooBKg9OKzJYij2B2UVlLCTqdv09IzGG1khgI3Ly8siSsojJds/2LN6y+cN4wZ7saPjU3VvNFuIKlCvu+WOW+y6k8PkxLjdvXvXbt++revm/nEP+KKTZn1jTd0DrGfCahBzmQdd37191+bmZm1+dk7XB7bBfd7e2xNZJIutdkedGgCnPA/uA0pxvsd+WYdAKtPF4vWgF9sJFOaMlsey7Ep2T4gbZT/Ybop0DRKKz8P9iFqFMwHf43kjOsVKTNkaI2QFeq3AnODfIJW8viRjAEwDIt3dMsjRQF7Jz8zPztg0vv6IdK1rX37xpS3fX7H1jQ1bWFyw7a113cPZuVk7PDxSJxkdZNhAQcqwntCtwphCBAlxxvuHvZPwkEQABKHAvhlW43yfa9PeFXgLIeFJkBjNuWFXrXouCSv6h+pMboNqhOjgTp0l7nDhgmG+704nDRuRJad3T6mDI5/TGs3aEvbZXJM6rFIXvhO8bgvvdarbRUG6Q3CAs/Ea73/nTWXVnB4d2shw2cPVi0V768mbtr21bavrq1qbj0/caht7umJpyKrsZ/unOkfRUSE5azrLqVZIzhVxboia5FV1md8KryPC+knn2ZR/xrODQOzXWeoeA4/DrsydWtijcXbBJlenLp3vIbTNlm8vWLXoJPX+4ZH2M8LozxFHtv2ifd0o9DsqmCsQgyK8W04Esm7R6c2c8DHrJw/mmGfxYK/un4GxU62OJRLVcTf+TUHuIumwTvQwdgigb4mKb6rYv/3en+QdgKhQ4JCjIO5bl4LFpMBPylgWPXVYcEDR2QnwJfm9sZB0ZEChyRWADyo41DwEXM/OzLjHYaOpAgXFBMoAte/mCwJq2DzYWGsnR7a1uSlfeR3y5Tc5rk2SAoffmZma1kaiRSvHwoDVFIx5WaAvCzKLqwpTMhmUp0CrYllAxCltqy/XRFCopQp2PFkSJE10Ooj60QgQKavwcuIh2TSFkl3X4gc4715woE8gaSJ2uDkO5id1ZAS6JoYe5QkLDgQCz4GFvqtgKdQU+BDmBWzR2XJ+eS5bI4WVXdat3iSEraJAMvk3JsJIOVKhuoswQjpmCs6qe3cLXrpl73AAOK97wU5rtgN8fh9kcUB+gjYDV7w6adHTwSWADQp+7Em6PYBdQucoCij+VdZNqAAAIABJREFU2jY2N9XfSOI+xMF4AGT6oT57YNeG3PcYdNC4v+EIsOq5kgfPyAtagZt966fY5BTGSXGaLLsY39jBxBcbXHS5iIDo+nOKdtL4Pn+PzTDUB0FGaQxIYTsAJqRwUYu7e5+eXZxbCcZ9ygPsL05ObWN1zboUj+yj/Kr3wKZd23MqmpfebZEF+vsX/1+4oyILFApk0OfzjoUwMaFgiUNEFGnftDB+HVD0db8T0LIOGGmTF2iD4kp+td4azEGONYqCGIJPba2O3XuhlSVSuPoI/k7j2sHAhGb2JcWpvTLB25QxXRTzIj98fsh6LLXteulxPVh08Hm9/dnXV8HtwU06CJ7ztcvVQGHRE7kV/jnULp1eXxZxkKgZ2E5wZuqwkvqFwj0DlgXQ3Mf1E4HB373bzcF/L6KcuI7CmgNdogeshwoxck+SAig+J3Mg8iGcmNWsdj9YdWnormkEsYf4V3SXpI6cQKdi7UqdK7wOB2V/UinDAUVRqPAz19S/PgWj+TPxLt0MeCgnnfS8pEZyKxgV6QKQ05zEc7nvaY39AJ1s6XVc7qV7FmoeI8clZRFQALuVgpMLOanEsYvgyfWs1XTLBEDPZgtPWz8w9zX6kdeQrKi8M8DDlyPInP3GO0kGREwokX3eRvaDPw/5YSdittvFTin2PAcUfR1kHfKn4xy6E1v9NRrVUv+Q4N00PoI0mkSKaUyk39ef4of6XIR7DMdBCEZAREXskdqHB8QbL9Gfd+lZ95VWGvtOLDhR5/OeedIeYt9IHTMZkoLPojmbAYU5OMgnNz4+4LBsglzpzugrpBwJrBv6+5Gs5vpPzS3KYqwzn1Kbtvyv2bPC+il91gBuO8ZeG5lAQVJ4h4DP5oHH3DVwW9No0HUVXbP+/M2W7t+1H/34L6xYrNj+/pEeLYrQONgGgEdtEOQBL4n9J5Zv1AoQFd6l0hWAFEQFXu7ss95RwaGL7x1RXolscJUrNWTKZ+i0rFm/6NdJvA+vzwGP8E/ZeKIoJ3ugBFGBUMbsw1/9yg53N35vosLrh7SGZgMhQoiQSCTdx4z10zftX1GPqFZK4Fm2lvDHkAjMG0TFtddVkTYA6qPW0fzSeucEbxBvEpoAGis3aGD7Feuc/yz/G1g5YDVJvThHjoGmpdf6zPF47m5P4jVf/I9rCFLBMyoA0v09+zVPBhxwAn1AclO3+H3yro24H9mf6e+DfQupQbcXv0tHRYTl8rMOUnpGhX43n7O/fPefCcyrVseljgVABNiiMwcL0OOTY3v7yes2NlJWFxQWfIdHJ3Z0QkD8gY1Wx0RUfPDd90UUo1JmV0ahjDIyXxwW6QFoCJCFBUxpqGuToxX5cl+dHtrMzKRNzE7J1jNXKogYAizmbDIzv6g1FLul88u6ffTxCzusHdvKgweya2HOPHj4SDZJkBQv19bs/vJ929nZttGxcX1mbF9Gx6vqUiBrgzGD9//21q7mBBZ3Z6fHUqcCrtB1tnLvroAkzlCAoa2u2dbOvoI/sauApMjj3V4Ysr/6q79AeqzzBaCreHaBVoD4nKXcNo/9P1dIAcypwzBH17iCb3PWvEQARdcOwGNDndafP/vSLpVHwxrr84LzmNcuqMirUkzzfuq+bzRkxbu+se02I4z1FG5NVzykBDZPnO/wBueMJ7IDMV3BOxgF9mkdBCh1tgqVOveCOQAppHOcYbdBHp//F19/OircxpasIxwCUME6CM7vAdLxWiVCVIcgV8si1N588thee/RAwCr7+tnxsa29WNVZE/EB3WvMtwePHts/+8lPWOHt2ZfP7bLRsnsrK8oH6OWHrDRasmKlZFfp/ilbOdmpkJlC+DNnamYC9w/An7UZ27OLs1PtTwVq3XZb2R2NywudJacmJuzi/Mwe3Llr85PTut+Mx4mpGTs4PrXNvT2rjI7acHXEupBdEp65xRteiH52cgAZsBe7paeffGaPVh7aUKtrhzt79s6bb9nqi5f2648+FHgmAA9xA1kk2KkUi1LqeydCRbldq6urWnsgMjiTQ1aMjo4JWGeMkBnAPaC+R+zF33ldzw3wc7cDkt71z3Xy9wApA7BlfKCml+Ci650wjJHIEOD3Q80fGY8IAXnGM9MTui6AcoSXF+d1azapb7o2NTVhZxcnuo75GbcNmpgYs2plRLkp4BeA1OypfE4IAQg6rodcJs4qdIJTSyJCmJ2f0Tmx0x2y86u61OiFYQ/aZR/uKnPDLUYFyqvLzHMNZ2am1cHPPaCjg+tl7SYngnEtsLSLAt/lSN6JULS33npDJAznW+Eu01N2dFjT/d7a2vazCfMbHIaA5XxOhBTz4qJ+qb0Iyz1ZvaWMCLqI1YXlxaKfZzodxzGGC/08GheB+V4TXa58Hl7HnTTIrQBLcLvqELS4laSLeXjGcS7sYy7M/SRgm0bkSV7kzLTWGMSVEKHsE+yN3CvEoOyJAPqs+c+ePdP3ICp4fbI86Hhj7+S+QmIhvNX4TIKQOF/GHsrawTWyF+GG4WQGXV9XfeGkMpVkPex1tbI4Ef8lO6fAYNw6y2tNdZKlOjuIDa/PyQlN7h6EYisYvKj7Ri4nz5c9iT0xbPUgKyJbUMLNNI/6ApeE/zBv6NpgXeSZYPf8+NF9e+3hitYXyCcqC0js20u37T/8w38QzkEdoJw4bPWu6iKr6VK5ajRs5wDwnsycZGGdyG/V2MlCMmqpLGHx1dosBA8DvC7bVdWvxfpnKs/W8nrGuzTb1OMiuEpWwBYLsngIkmvI5qcnrVJADNm0k/MrG61WZKUInqhujh7dJX6GomYlLB4ijlyeW/NzdnVZt9Oz89T5mUudwiUnz9vY4CG0oFvJLaJY91jXwUUjY4fxznuwv0BiikhKZwplmn7bUfG7SvZvv/+ndgfm5XVJOz4LC22MtMvS1l/R5hPp9FLIsBHkzMqVEU1AiiIKL1pH6XRQh4NakwpqrUV9Xy5iw+QteexyFDVMYhZfijzfiBxsontifWNdoEazSXglocdDCi2jiKV4UGjVxISIDzZSD0KiOwCvQvdLR1lEkBV+cNo4ZENV1GGcQv35i+e2trFtR7QXj3l+AdejPTQpFn1TTaBTbLB9FMIByMiPcGbfN0q1lgoIdXUaC3qAPVEw9VsaZS3lILisA2jLpjuC18m7IgiQlYM6/6OtuFwp2qRaJjmgoqg0qx2fWL3eliKGLgjlbnSdRZfvXlr7PZyKewVD7h0W6pJIVlkKnEutg2wqBJtxcGCT5j56LoeDWtFGDRmgDSQHUeSZEKhL6KRAZUQ7cqNFqBM/RyHZlvUTGyJs8kA5EfYwobj+ZqKCa+D+9h9JImMAilEc4Z/KtRWGS1I9xOYW1k98zgBqg6bog6vpMK2xXPCAsSg4QkUYoWMCGZPSK4gsxvlNz2k2GrHdqSA+oeWzUjaCLXnt8+MT21xblxdzqewEkoi2pO5hcEoddIk1CUrir9oyeehqAhlvdAf8P+mocPzmelaA3ysh804mJvBTWRu05fczCL55RfxjiAodzlNXTPw+xQgHfezTqDLoqmKMdztN70oZcpuKsDrz33dli7NKyU5J4KYfYPqAky8M6a9eJPa/n4C/6DpTCHG0mqvq9tZ8WcMl8FKHTZ28PTSNz6BDnIL9IFcgGQfho9x9BdpHoKr8ymmFd79UrXFSZyfENAMyxXgQgHVN553advWaHMIcludLxLUfSfygh28/BJoISQe2KWQ19lFT9f31A7xyolRFfQVg0hXAPofce1MkkuyLPKjZ393B9gATs4oYJ1pYD+nsanrGj7r+3HOWg57IaO491lipwyTGre5xRrEdhCwLlwMZhOLRdp3C4aMjIriJdKgV4AtwxmGzhR2Erw+iXRIhrXWFcZXa3QWEYNkwTLiaA7UOmuetNFL1TjYO4G0sCFHoOdmHwtZts/zJ6f8nm8YQBQWXKQhzaBCExzXIzg6wX8G8fgAE3FQwdgLRKY49OBwVFRkUA9JW9xwbEvyBUWwCSmBBIMDEn6WuLd1bYeZJLd2/jwlcUYt4misxZ/XfXgAMCWSQH66PM54nBwgnFxNBkcaoH9Bz/WfG2JS1YAJtUYL6mhTWSsnCCAuAHgeP1C8U3TFpdpMVpefIvwuwgJhgHnjweFfzqCu/eVe5u3mT5kQKJhepEURF6oyTulyAlxPfTtT5b/eJkfQvrD/xXAneDfUd5GG2o0LdXFlyJEjFdIjN3mfdK/knOwDx5nvv2NvvvCcV2P7+sd6ZIEwHAHxNARDg57OgNUApCm9qBvY06kPGAWMNMoLuT4gKhYHK+oWa7VIHMAKRB0QDF+t7GIfqZuNSB7XYQ1nLAVawZhiGqJAS0G3TOEAy7z/57W9t4+UXfyBRkYiDqO8y21OslfrW70lUxDhkzGbtkvp7RxDYmY7HV+2IvuwNbI+u/Yz2iwFRofkquz1XA+PnHF9BHDiQwfx0a58I0ya8cmZm1tfsrj/rUFDyO7IlSft3gCEBvgSw8nVEhe9Pg30qiN4BUeHqzpjPWQAiiIqoB2MMxucq5fMeXJx8vPtERcoDY0x//8H7dnJ8YbNzt6R4Bcw7BdRDQZzPKXjyg/fese2NdZudmbLHj1+zFy/XbXf/0PYOahrLAC2PHj40QnOxguCM8/SzZ/bBd9+2Vrtrl42m1WrHGoeX56dWyplNjFZseWnezg521JW0uLxkc7cXBWCROcT9Bni4OL2w4UpVeVhb23v264+/NKzDq6NjIibYRyAkqM+bAi3Io5i2p599Zo8eP9a8A+SFUDw83LWFxUXtQ3TZbG/v6eywvHxfZAtEBV1fhaGOjVWrdn56Jmudo9qJWb5km1u76j6FcCgMDdnYaNly3ZZ98P57Nj5asVyOMxvd0HTIYjnEtU16lgfkLZ76SawgcgLATN7abZEV8PYj7HcoeZsN7Y941pPHAOl/eFATyLe/f2DVUTopBjl4TkC4xS7P5PnLNTu/qGv/gYjgHinHoDJiRbq2RGC4DUaDjLQLfLt9nvfXLuqGekNruzoBUqZMqOpRnzNOfLr27O7yHTuicyKd0bTnF8nl4Vkdy950emZWVjL1OiHBbREBiwtz9s9//F8J0D4/ObFnnz+11ecvbGOzZiOjrIluS8SeytnkL37yE7v/4KGsoLZ395UZQe7I6uaGzSzN2EWzrryTk4tTWYLIL17CBBcHRS7d0cmJyKvjo2Op9RE7CIDm/EYGA+s/Ac+Vit1ZWhJxkUNw0YU8HiajWcHy+9hmFYqe1ZQzGyavZGrSclIR+/mRNQX3gcmpyaT8zdv5ybkd12r25sPXbXdz2/K9IXu08sB++ctf6vmDD0AoYJ/FyoQqn2u9al7pNbmnkIBjdCKRryF7aM+UY01gXeJ5kgXAfkkXPCQN44Z7yjk7VOesiRBLIjmuvKMiAHyeLmC0SIuiiwIZY+AL5CGFYE4WPxKzDEQEgPqzs9MaF1Vlw3DdWBaaxh0ZFVjcsH+PV8eEZ7CPce6jCwcrJs7IXC/76szMlMBihb0jKux27PbSgl1enFrt6MD29k9tZq6qsPV2b8i29mp21era2NS0MkJODg7t7IRuMLdS0vrdcuspxjFkGpklHgbvXVredVJUHSICUeSOWWXYSeSV+8s2OlrVvPUdpCebG14fsJnuKvbl45MTH2szM7J8Rmh6cn6m8YhwEqeKk9Nz3T/IGGoJnpGEpDhcFAuqH84vzzSeOKOztgdYH0JCCWCTKAhSEwwiQuTjHEb9MTij+37GOuS5DJ6bAWEIWXHv9m07OzlWBg21jMRt5Gsk+0bwG8dGUsdJviALPicacEPwAGw+I2MEpTz2WHTGxJk8uh5E5LVaul/cU66XDhQ6sbD34zqj04LX9m5FPwty3aG259yisw51cRIgXasPXH/RP/sHuRG4WtwHyCHGOXsK41BBz8fHIt5EcaUjLnPOxUl+JnWHkCSuQRCo8wpCGdbEvM6G95fv2MrdO3aQOv2a9bpcTbAU++jXv1a9Qqf47t6xzc14lw/rP1aF+7Uje7G2JQ1GkxdFOKu8V/Jmo0t9EKj9u4iKIKj4HOGUEXtBWID6z6QudJ3T3fiXe+BQJedrCHzmTFM4Qnm4YGMjw9ZJ9vOs05wGCaVnPXKhiXeUsgZwf9mv6g1swCAKwSrLtr6+kUijksTYCIrJjIH4psMMMod1jstiPDJ39TqpK0dEIR1Gw8MStPE+sc9JHPctUfHNoNO33/3TuwP/4slbCkfEd3B+dravlGMhYmFhQ3758oUOCXjbUlzhlcnBlJCXUJ+zKMhDVIos939DASUwhwJLXn6eU0Dx57kJfkhXF3piybV5nZ/Y2PioQrRZ4MslD4Fi4SYEi9+F5JiampJOGkCDVl82ASxMFCAmBQbhyB0r0qLW6tjTzz+33/zmt3ZJu3KpqEWbgpgC1fMnMj7s/eOvr95aNMXcJ7/7pAJS0auFPXVPdLBrosAH9PK2TP++L/zuueiAoAIiI7sC2ySUFXlv45JFEx0ggIEKaeOz09I+LEYaYgZbJgCQg8MjO6idWh1v1OERFSvcYxQP5Ii4mojApLZwwAgMRlXCIkgLH5sZgC7qFnksqmj3bgN5L6I2Sgpu2jfDh57n7UBKyuhILWjtdl3BYij6Wu261MFO6HRsdG7yjyYquHcO9LkVV3wJpE+K9t+PqPCiTc8zAyY4cOIsPs/s1vzt5Jd90Qdfwx7BWW0/fDAf+qoRKe2vGz1ArqE+5QurtOioILSM94Ko2Hi5ZuPVEZucGbfTk1MVE4xzMir4vL+LqMiq9wNAGdyfbwjTTp9fP/uKjIoAKvh2FvgW4JAb9B+p/RflTz/T5Hevh384UeEqkix5xP1zBS9KhLqURKNVFHE1hbSCBjjB5FYxFA3ehuvkRYAnAnSSEnTwLN2CLVQsXhz77+i+0AKv0MbUTopiTOFyHakIackPwD3AF71vj4LX1aUADSwJDsB39FpF3VcHJmMsMsf0WoC3qdNMhEd6Lq6k8Xsea0w8gQDjs08kGkV4jgKyIClFMDgQzWtFO3K768ABr6uW4Rxe9EkdnQl4j5/nZ4OAVZdeat8NAsMvOhWHSXfv2K53G3g3gl+tg4CQH96Wz9oaX1Ja4/+Lyi61jF9DLnWW90A1v+8O+Acgy5rkz8AZibhvcc/7pDMAdiJf/JDXlNpmcmKyT+j64cjXlABcWTd1SJan/6gND9PumwIlIULLFXnmcu8p7jnE0YLMusphXhkVQVQkFT6HA7JRUPkEcM24cf96D8Hkfmi9UMdcQSQNBDlgL4cyH0sF3TO63Hgd5oRCdlPLN5+F12Dv18FRns3up5sFMfVMkwWi37fINUjdRenno3uOZxeHIXVYMGcE3jT6tnGyJaw3rDxS6RN9XwE2FRLo5BRfXIcAeUgwS50haW4NxrSv7RxclavCNpvUYxoLKAw1v7C58BZ3dX6ncdMW4elEsR90nMTVPdN9vK5uj+8BWoogUseGk2GxrronbpA/AwKIFYCMjLPzS/c5TnWNn0vJ2QiiwvtUnNzwtSnWhFhf4/DOOJyambYf/vjPbHxyxjqdIdvdrblSueqe3vH76soEsEivy2sGUcF6y1iJPQ27P/JVICquZ1SkjgpU3qmjAnBQ5EwiKhBjoN4WcJLmINfJwQzwaJhAdK012HeiUqabrmjra2v26cf/+J+FqNCzCEvANCav5aN8zVYW+0UQQdl1V2RAluC/EaadfUlVCxmiIkua0METaxNjJUhyulXC8jNI7L6laCIqqLeCpGYvwmKF5y/F6g2ign+TuCYI20xHa5CHCgRNGRV9EDgJO64RFYkA5jMSEBtzPoQusR+FHMDH6aBj7+YeBlGByCj2uyxRAQAHUP7O7bfs4w9/Y3/2ox/b0tJd+/WvP1JXBfeV7BnyD7733ru2s7VuleFhBcYen55bvdFWOC1qV0CsJ2+8bjs7WwL0qI031lbt3t27dsn5Yihvh7UjB8MYr626zUyM2ttvPLaTfUK2p2x2Yc72avs2v3hLINnW5pbdml/Ua12ixDy9UFDts2dbdlg79wDXo2MbGx+zhcUlqa9ZLz799DNbXFxU5gIEk4Q5UrLn7MXLTfvggzdFQiMs2Nnek08/w2hjY83m5qal5iYj6sH9ZYF03vnbtdrxme3s1YxML/ayVv1SQae9dsMe3LtjD5bvqkN9eKRopXLR6pfndn5O533PpmbnBORw9uD+YWfTaZkd1A6UNQB4onw9gGACgycmlTWBIOfguGaTszO2u7lje3t7sj8CwGbd56zGmgJwyJ7ZrNN5v6cZhDCO3ITVtTV7+XLN9g/oABsyMi30TCxnTc6PhDTTJSLrUe8ACMWxzkIJ8AN0JMCZ99b+2sEWaTJZDHNewUJrWT9DLetq1qb2b34HRwCeP8p0VLI8j163aSPlgi0uzNuffe8De/rpb+zLp09tb/vIhks9m5qasauWd02dX15IXME8Y9z+t//dfy/SZXNry7Z3du31J2/axtamHTdO7f6jBwLBh4p5jQmeL+KIVr2RvCoJns3bz//Tz5PobFh7P2NzYf6WNS8vLAcQa2YPlu/Z3aU7ArebV3WBhDaUl4Uh2YytTs8mpmZFJjE2zi4vtK+zTI+MjdjM7LRdXJ7L3gfBFxabrOOQWJxXjw+O1EnznTfftb//dz+1leX72iv/5m/+Rms22SicR2Ud3elJdc/8LxVyer2p6UnvUriA2D6z8eqo4wQSjBU03gC0WZePTo41n9wSqCybI53LOr4Ps0PKMqpR7+/xEBhgFLwW6nfOKhKVdXupe8YFIVobU7cnezb1DOfksXFyH6pWq9VsbHTcGvWmZ9y0e3ofuhhOzo51Np+ZnBHJyZyT5VHdMwx4WUgubJZkm1Ys2vTUlLWwohrq2sTYqL3+eAWFiM7On376qT1/uW/NXsdKoyN2cFK3VgirIPcQf5KLorqYtYFzMWfknHJ4qP/ARTxzzzsVfK9KYb0FgHGAfO9ovnd3UWQRc4eAX+q/hYUFZSlQp0UeBjcO3AhlPOuq1pFux/ZEPI6KRKUThGe5ur7ha0JuyJbvLdv25pYdHx9JcFqqlNTlkT3PSxwSNaPqEceOeE/ZjBexoXKRorprWm5FxmdzoSggf0Ge/+AOcqDqdiX2nJ6Y1NxYWV4WPsWcg9XkOdDpxhqEYIj7hQC3ftXQfPCzpSvuGS9gLIwBcKSz8wsBxmH5FDUAayF1N3UNIlCuGSKGa3SSzXc/78akmybyT+mmdwcQvqJ24zNFd2vUwi5OG5z3Qsw0Kls6CPEtP0tRH/PepaLNQHy13ZmEoGvhKDm3DwvhadTnXncgzPIuqugwYggiVr68OJfd3cMV1pYFazXqVsgN2d72ttZLPasWHYKnqhUh6HZ39mxvD1IQ8iVnI6NVOzg+8243cC86asBQ5Nbhot/A5mJcRN11sywTZpVyh0I8EmfPqImjtlAOimzYeaZtP4/qdnIG5TyfkxjJCU1yfyo2MVZVluj5ZUN73QiYDlaEZxCULihU18yI53CAlUE6QE6NjU1o3m1v7+q+QIK49bcLFtmLyNGi04jXi1wl7oO6frRelPSRWY94fhCxrIPkr4CDgpd+S1R8TbH+7T//6d6BWyj+06bM4sSGxGwFwCC0DYU0inrPomhZG+4VAC6pp5wBbmsxChachTPYXGU2JGCPoiUUEuH1Hi18YYsACLO4cEuKDw7CgIpSIQokoTvD/d84EHOdKBikGsg5MEYtKsad80mO4q5tm1s79nx11U5OzlKbvPvKc+1sgEx+CimUX2xYX/3yxVIthskX0YPG/dCYBW68BdXBNNqIQ7nTtxNKobfe7YBnZ8MBbqkosV+qWOPKO0MgEioocHMUc0MK8wHUqlZpufQuEDG6F1fqEOmRp5DzNmiKDgV4ASpGIBPuf7pvDsgB8LH4sUjy97jXEC0ADxSPFOhSMiRbA23kFJiJ4XdCZnAvZYMjD0YIDGxLCAxPwdptig2Iij/O+ikAqQAZr4HJCdS82VGRHy6pQAwWns+kttakMNVrJgBJdgqJdKLwYSzcurWkDUPteql44DMLkE2BbRxoUbVAtkUXjgDREOEPmTJV2ET4d4rrC+5veVjFEHPp9OjENlZX1S1DQXxUq+nggbdmeKjjg4n1UwBl2Y1XQNcNtXF2M/+mjoprryOiQjB4mgaDgOOs2tGBBbkAeDeCVMIdFeHhm5rlP75uhfxDiQqJyHRwKQqQ9PfOaY3i8Ed4OwcG1gmKKFnnEFpPMQt4rg4Y1pEESgcYXoxA2+S2peD38LlJViCyAOr6c04KFlqDWWfUGUER26Zw5vDbsQKBaZVyv6D2t0pdByIZU26M2s8pNLrqpBoeLlpP7abmIXpSwyelKm2qyZKI5+EHj2QFgwJGwJiHramY9arMW6pT50sMS11N6tLgXsqnVFYHyZpJino/uEE68j3GrtYKSNZhDwikvlNIJQfRtBZEwGx0jDiQm1HmqAOES3NS20mKQQCy3/zw38fWgfnmbfysmVh8Ma9FVKB+A0jPkgSRw6EOhKROSgo5XlkgdQIGg0B2P3e/bwHMBWjfYh2TOjmndZk1mgNdebiiQwtKKz5fkFj+Wn7IxeOZ58g1Yv1E0CsFu4KBGSPpkMVe1Go0rNmoa13mgMnB3UkyP1gO+HM6XFxJBoCdoGkHsFOmCtfiYX1l3T9AU0AFCnQ/LPleF+s514biRwGmKGNRuNHVkUDUIf2uK4Z4jywxkytw35xUkr0SZFKy9xDlxr4cBHM6kLkFn+uuJT7AK5eCWwA5ivqGSBXtz0VXAUZ7O59NIX+JWBTICnmU2qAbrYvkhe9kgh/m/I9BaLgyzAmsJKTVnsVE4VBIcKVaK7rJXmGoJ89wuhSZ8/KJlh+/d4D4ePX3CbLW2/dNCmmNf1k0pHHCjs0YyEMG+PcAHVFWeVdRzuqtjjU7HTs/vXCTvdQnjiBeAAAgAElEQVTF8WqiYmDXE/VUf31NXUOAOiuPHtl73/+edQC9O0N2eHise0AOBCCLc3b+fAH4/O9+aM4SFRw88Q3n3kEqHB0dfpWoEMF+JcVhEBWuThxk4LAG0FEhUt4Zw+T33ExEBRYxCFUK6vYV0VYkUPvQfvUf/yGpiwPyHuw01zIq0poZe1087+gji8/XJwj6dnvfXNsHYBD1xM2fvkZWfANRoboyY/2UJSq0E4eNWyIqfF33/QSiXPYFyYLT8djQwybLFn40N2Szc3M2NT3tB/+egyWx3mXndNYuRb+qrjcy5b5q/RT3NMgSnxMDn26ICua4LBgSOBOvlyUq3KrN51rsk3E/qffPT1NwelJb9q2f0pr07u137MXzVXv46LFVKqipG/LTX9/aVJcxdSwgfLfVsKnJCc3R47NzdVTUjrBcKNrVxbn9xV/8c63tWC588fSpFNT379/XOvpyY0sd2xKnXF4oA4Iw7YXZKbs6ObDJyTG7ff+OVcZGrNlryW8b65f9rR0bGRmzSnVMXUx7tZr9/c8+tE6ra288ecM+f/qlTc9M2cTUlNu1XF1JeYmPO4AgXQfRAU19cHR0YAsLtwREzkzP2fNnL61QdPKQc5vyp9rsJ1e2cGve6hcX6gAg6Pmi3rSt7X1ldnm2YMfGRkrWbV7ZUKtpd2/fEiA7NTNqlapbE7Io7mHJc35p49PTmn+FEop3QEMHrOm6B5Q5PqxZBcKhTsi0E8FTc7O2tHxPeQp0PyIow/qDcQCwyTiAmGZNERhZcrsY1oTjszMJprCKQ6m9vrFp65u76rLAQohnS7cLABPXJYuoTls1YQTWBiHOGARg4nwjleqVe8sHAVYdDfDbg27discDamVV1O1JBQshIs98FK3Y8J4dWaVctJHyiP3oz75jz55+pvtQSh7w3aGi9YojIl7omvQue++We+PNt+z9D75r5eqoffLJp5Yvlmz5wYr94te/sNHJCatOjAkEhpSUEI/ZwfkrCcnW1tdsd39P49frYZPlE2RRvtezB/eWbXZyyoYR+CBmcDROIcFbewdWr2OPOmRHp2d2eEDHTd5u3bql+mpyetIaTXIQGxK6jc+M2/BI2SrVqroL1cGfukOpXV98/swe3ltR9sX+zq4Ivn/8x3+01dWw6PN9jS+eFefJNuMUm16CmM8djMPaGfEkz4U6xM/IZJtcSryAwJAaA3tp1i0+rz5/2rt47oDDgODRea8zLx0+DeoM5rCTOsreSN3VImLDYlR1KfWjh2tTakxOjWuNoOMjny/Z2dmVCAvq0cXbS3ZwsKez/MTYhB3sHwisZG+B0CMwlxoFIgwhFbUVOMudu7et3byy6YmqlYt5W769aL1m3caSaPDismEbu/u2dXhsjV7eRsandPYHEGZcsmdTg0gEin1OvaHzBNaqnN/jrEbeIjUo18NeShB3rwNwzn3r2Uh52G7dmk+iCM+TGy5hu9TUvQwbLZ4f9kUSvaQ8EED/egsroVPv3KDLpNlStxjgLPePmpk5RXcJjhdT01N2cRUgP3aQntvpdXkKe+53R/h5TFk41MspYJ3rdiso71h3YUVkVxBcfy7HDertcrFgE2R2dLDhIR+j47ZTSYRDTSdshLr57EyCNzIq9g/oIHWbORdykMfpThPcW4WHp9xEXSOftQE5wdnPXSt4f7+PFRe99kVhyUJNAgEX3bi4xddUzikC3JOVlrJTOh0B4llRhOMOLvpRF8to1f76r//a/u7v/k7vL0ys7R1pXIvseHumjgp+F+KZFTTERPGs43XV3RRCXdkjUX/zObDIytmbbzxW6PRxbV/ZPFi3cy6cnZ23g1rNWvWWugXAt8D3qLupLyGBarUT29rb17pz1aL+9owcdztINXNk4vY7879a73kdMrCcjBomRI19AjKtEZoXiJF0OPYWahdAQOpju8Q9A5MrWqN+aZOTVRvDWrCdxjPnDfapbs8OaofuAJMyALnXnPkgX+mW5NyMsJpxjSWcP2uTEJzrYH9X1+UFZFnZ6hCX7GUpjJ0uZWpsfz6sR9h6lTR+2YfieX1LVHxzvf7td/9E78D0JUp+P2AntCMTOlZw8AcQKXnoYqtB268Cj2CuYYZlSeC+3PJVT5Y+HASczXVbFS2ISQ0LUCKyIgFOFN0cJFhgxynKyQWgdY5WP/m94XfsEJvb9vhizfUJDACAaLFwAloxwfP27NlL+/z5Sw/upl1PCviKQp/wIYyWNpEtdF4kq6TsowxwEVQtgEGWSB1Qw3M9WT34oc83O1fjpXBYABwRFK7s5Yv3k/otWUPISzjXExEBQDOJeoTF0kwhXljOjowMW6lI+FVeCysH9qtGyy7qLfvs8+dWHK6a1vkhQNyeADAPYnbwrQVhkNZx7hsLIgUim28Hr9dUODIeKOBZCGX3BKCSfDW51ygERBYkOyh9pByKcNQLHkzUaQMywYp7RwWMNW3kgDlj85PpOSYFcEalfk1xnVH0eQHgYEmWqNAmI2W/jy8yKgCLCaWVQoECpexgMWORZ4yyUMBCyhjhEMzrsMhTWLq9BGBeUQAJCjdILkBDihD507YaannkUOjMdkPjzwkRLyK06SVAe37hlg5VfEnlgrVZpaKNivuIDygKUTqDOIiiEBLYCUFXLOn58G90XgRREYVKgFE3w0ODWNAY0+kmC1EPRnkWFMn8ayIwuTdujxM/F38WQJ46KvgMjCm11/c7Xa4XE9n3efV7vnoRFZGWFic+U3TUSHFC4Uoo+tiYDoxXjXMrlz3czb29PWOARUx2ScOQnIMir3/vwuxIbSIJ6BEg0neC7+cVeCePq154Nn7YH1gNDICbFH6bFC8xJrSOCHhCge9qEcYs/8J66orhAG04RA3IhyAW+ncq1PuvCIAOEE2Ff3QNabL4tQqs1whDIeQkhRe6Ps6j0ItOCootviLLxuejV8gBWut1UTOV/DME+CVlY1on49kHOBgqL/93B6o8O8LnEtfBfkNxB0jE3zmcUfR7t8rg8CtLhD4h4ci0FLfpSh2Uc8V/kJdOOAPOA0pQeDsgzu+GwhjbKdmspIMHHtEESPIcIcNpBedZai+RGs7vC8CLckZSXkisK9xDfpb/xr4S6jAONE5UYAPVSv7Dg6Bhn/d+OIu1MJTwcW8jDNJfCzK+aKVSxcPHyTtKHQUieBLBEusFlimy9Uhkrp75cFlDJcDIUF/Hmuz2X06QRRcBvxevyc+FSis6crJjnM+kQNm61yNxz0LVz7zgcC2Fo0JPGQ/uE+wqN59HCt9MqlwpVpOYIIAoH/5O8qvrJ3VWxZzNrkCxn8eqKeg35T/Fdd1cx4LoiuuJOci1hTVZEIe+prkXsr8X1+Vkn7p3sF6DBGgw73LqrIBc8NwNz6jwusyvOt6T+c6eFrWGdP0CgXMK//vhn/3IJufmfd/vdBU6zFoK+YjlQxsTq0RUZA/+vMdNogJglC8AntMT7J28u02dhsljF7BI1gj5IScaZEHhtZI6lnh2dNQkVazIwARU7u3tWCnnIbkAkASnsodziCQ/6+f//u+tTd3B/dOa6j7drzrGftP+43NqUATHuOKzXQMEXr1F9ffHmA/Xasi0Nt8cK/39WwrCjLAhdcjFWLr5lv0aKTpnkh+725V4gLx3EHUFLgYRwd9R72Obqq7arheDsaeqNpH/fsvzjDgXJEcIQFG+ACx7dFRoDfV5FwCA1wP+v/wQBCpEH4KBM41VLElQxodV4M37EeRwfG5fg5OgAEuRiytrY5mD/QzzJOe2rgIa83l7Z/Fte/HipT158123ZrrEOuxQ3uJYPzEHH95fFng/NUEn65Asn84uLu34+NRrw7zZ/eV7AhL52t7cUN7Fo8ePNO82tnYElrFHnxOEWz+3B3eX7N7tW3a8v23jE1V7+Poje7n2wl575y07PTuxy/MLKXkhBeneIOfh8OTEnn62Zp12TucXZR0MD0tlTJ0ICXeJSKxSsd29XRGC0TVIFsLLtQ174/UHLrZqdmxvr6Z6HeD2sHZg5UpJClC6cVfu33OhUbur7oTTsytb39q1cqVqBZ5jB3uggl2eH1s5N2TjI8NWqRRsenZCZw0AO8j2nsZXXoHcnONm5+ek4i6Vqv06lz10d3vHrs4vbIjaJtnuoPq/fe+ezo7sm6jJqaMBNkNVWx3xYGqvM7yOkHKaDsZ2S/7eWGwAqpOp8HJ1UypoiJ+KfhfCoq3PSK0AIMz9E1grgtqFcvyZ95AveAtA1z3Xub8utDCbmHQbH/Ya7VfqEB3W36lxWac5L6jOYRwOsfcMqTPln//oh0bWU213x3a3tnQ/zq/a1uwhakne+ljzJJCY9fkv/+uf2L0HKwqdPTw6sonJSatMjNiXqy9sbmFBqxr3TmdG9jUUzaVhe/78ua2ur8nmqNmCRDTl3I2PjtmDZQiKST64lXIFK6dQ4b3tXdVrOweHdt7o6BkwT7BKZs5yfpYCvVSSYBCbnPlbc9xe6+QJvG1pvRqbmBQ5QGcLAghCl1v1pq09X7Uf/eCHdkKn/8Ghvf/+d+3v/vZvFSBPbdnr+lyEdNDaVMgJtJ+enhJJxdkVu0WJCCVUAMTuScHN8xXxmTp2qRfYw9k7Yj1lT/OMClfxh1Jdey11hDqLwCb8jMe/ASayZjIuOHdJUJnIC/4dmyvmSqvdUNerK/bLdn6KxTA2piaQf28f+zcENBWp1XEoYD/E2gqCjHMI45I6hfqXmmdsdETiB4D8995+aBXmytysVUt+Lkd4WDu5sMOzS7vqml0027JXHKmWRZ4JB0EohLCEboBEFLuFttuTSkCYQ1iU7RpGkBFOEAhN/YzH+Z5zKJ0HnBvCEz8reiLbgfvjdtK+54ORNFCzF0uyhmK+MaaoPUKYgPAVG0jOO+xFFwgUCOQm6yCd15Q5krAkJyyT/ZD2G6Eqwk/62XeJbPduBepcVOc9iZia5CXkTR0sl2dnCq+nesJeh2cICQyOUqo4+SV3DUjYQkHd0pvb21LAc1anjta9JYxdNj4lw9pWbgrKRvRuVn6XcekAstdzED3n52eyweL+Mm94Zjx/aiXWQmWlyvbUn0PUIIEz8ayCzAhBbZAy2fO5n2vM7t27qy5EsAVEqJCzslBP2UCMdQgZCWK0ryeXgESOqBpKhZRscUVweSe2am11hbXs/vJtu3t70Y4OdtVRAVGxtvpS+WQLC4t2fHImDI5nvra2bdjW+v2dttHxUTmC7NWOVNuRs0rXIiSo2/QNqjnHGP0avx4/SDmSfEaNA3cqcBInsvjCGcU7XlX5Ofvrnef6jE7Oy64VvLNxZXOzjltdnbNu5YVXYg9FxgbrFgIjr6mZSzkbkdsGGCbZsdiVup07z5pueYg8hG68N7kwEF7qdIEAR0CcxIn8G+OHcSaxh5wOkljiqq5nC74m+95vrZ++pkL/9p//pO/A6AlBS1gjRWdFYqNhYJNdSlZdquA+TCAcgfWjnazYIxiRNqYEggkk4NCTWHux5f4LbE5Tk+NSXBAyBThCKy0T/PXXHmnRYEGVnUUKTA0PcF5Dikf5zLsqmMIRlSETenNz2371qw+VQeGt8b5gEXTTByHTU9Pil0CO+DxZWxgRDADZCizzTd1BBQ5cTnD4RusgNIsFBVYAFBQIstNIm6uyKGhNTmQFi6ACraWU5meHrVDKub9sPm+F7pCNFCEqcgq9K5UxqG8buy2HPoLxjs6vbHVtyzpDFM181ryUZCx+bIp4i8r/LxE13gVBeBYWT7SklhW2R7sgBVS0/6njI4VYCRrDRopCvVFPn9cP9oJyZauCF7sXmJASFD4AB+02hT2KUsDQjo3fmtLn9w3BN40ARdmIszBDHwjL2LK8iqgIKSssfrfV1kFJKoREVMThVyCH7HM8nI12ewd1vNiK7IO4vkp11FuRj0+kqKBo0CGIMKl2Q22B/J5aN2kNTT7tsaFmiQqFEgIGdFBgt7wLILWk1w4ObXtrS4FtDjC5BFiFAX66AHPNlp3Wat4SmiEW+2B7AqxeRSrc7Ki4CaS8ahFTMSBma6CO9DEeoZ/XiQrGMQeGaFm9CRf9sURFvGc8E55Vmoj6T6U0LI/UYilvzZYHd+rQmdRnWj9YM4oDO6H4DP17d6P40fMLADQF7MZBKABB/s7zQ6UW1xigjReaTgTEWIg1wcFsD2MMoCeA3BiD8XoBDN8sRLPPK1u4RTF38/PFve+DQJnQ0lBjiDDpd79dt5AJhT3F+f/N3ns/SX5l1503bXnvq6sN0A7AwAwwmBlAMySHmpG4CpIKhRSK2Ng/UKEIcoPUrugkrSLoYiSOAwa2AbQ35X1lZVZWmo3Pue9mvk40xoj8ZRRdJKa7qyozv9/3febec849N4i/WLP56wL0inUUNiKxzgPciuuP6w0wLb5P4MVewdyTsrLR9Ga1bUrdsShym5oeMB97eFYtET8LsJz3zv/e/6yoBEnNBVOVSdyz9qCif64UbCUHWyCCVXVAQnbuloYCjpICkHHieQaJIKI0JUFBUPBzkaZp7GV7IXLBPbPDX9lBFCeQ3D6FvcEBOhc2OnAYa8PJEve7hUTlZzRddRtCP6u5rthLc9CRz+WzAAbUS4HXJkA/Jz/z556v0RxgzZ9P7PfhNx3PPK4h7l02R6EkS3ZOca28B3/n2XA2BfFDEB/9lmJe9ImKfqVLzAEpyrPqmfy+Yizy8czXXw7OPmvfjGfA70WVqfbvlLR6DKH/daJCY9u3sBLoIPsdbDeKye6gYvsHnGnS7nnz+VSqns/j6GHiNgRpm4zG4qWS3bj5sr36+hvWLXlfLOaVExVt2ZqQWKGu03nfxjYs2TSlKkxAup3UowISLogK5iv9yrj3mPfMbcbNiYqDRFQMKdFFlYjFQ6gA282mEjHmO69RxWm3Y1sbG1YWUeGWZQgHsH9ST5Ju137+05/Y/vaOFSASfefXtWedVnqP6BedPzkZISA9Vd886/kOfm9wbnzVzweT619EVOT7/+DrnCgPMt1FRk5gs7b7ZIXmUceBq9h/AcLn5uZ8pLr9cyv261Abq6m8yH5P7iEHVDlz1lBvtIiJ47zwteRVcki6y0ZsXtI41mvHTsJXIei9KjkfsxivQaIi7lGxd7lkjeNT2Spy3ipmJ1YSUeHx3Osrr9qTJxs2P79kFy5eFgD74P4DO67VBBzu7+3bN77xdXucrJ9ef/3rdvv2XduBrDipud/4+Zm9+tor+hxArSdPHtvtu7fttTfetInJKfv008/dWqVUUU+CxumRTU2M2JW1FauUiAvrtnbpgk3PTFm32JFymDj0wcNHtrxyQbnI4f6xKjh++t5ntr6+a19/8+v2+e17Njc7bdevXbNa/dT29vft9u07dll9JfbdkiSRpBA+x8eHdmFt1aqVIQHn9Jkh93GRDc+buKOlPgTYE/FcAFC3d/akoKd5eLmMbSL5yKlNTdKced8mR0ZsWGBL3UZHqjY8BEBfkA0v46Nm1eqz5j00vI9QRb3paNIuW12q049qaiIO+KrGq6zPCt7jHZuemJCd0sTMjO3SF4CeYmPjqtaRj7/6T7lymn3lTM2tJ726r9O2jY2NJIZAeXpun3zyud198MiKFaq/iiJ3ATEBPDn/+B38xNGOEcsTPlK5D5BVrZR0zjLv2f90thYLtrS0IGsYqZFTtSb7nVeUUj3qMbz33zI7PTm2keGSLc9P2+//q+9buYDAjuq5c9ncfP7FY9vaPrFa7cw2tg7swtqygG56S3DeX7xy0X7wg+/rXH/w8J5y4RuvvWaPNrfs5OzMVi9fsV16AFWKathdOz6083rDPvnwY9lKca1t9V5q2ys3btqFxSUbAUQ7rtnczJwd7O3b1uamgP7N7W2BkvcfbtjRyZnVav7MoorRexhCXI+KrFFfQZ4X/W2WZ212ft4JBzP1GFlZWfZeDOOTGtPHqVfGN956S022l+YXdV796Z/+P5oHqNPZp6QYl4WyWzEyvvQkAuBFMLa5udmzV+SzeA4Ar5BP5Kjet8grq90OCAzDf8/jLm8yy/7HM2YuQGrw+wCB7L/8LueO27Kd9r34M9EMhzVCSqqwHj95rOcOQYB4DRAUooK8kjHaP9jX9SOsxM6Nec1ZjJUv60/gdONM4KJIYZrZj42KLKyfNOzqCxfshPc9ObUf/O539HN6y7z/4Uf28We3bX5pwYrqTVfQPsE5CKk1PzsrMN2rP1y0oVg82QU1m04gUJnEGqKqIXoqkM+ztrSWiV9bKLtrCadp9IRAqvgVoYcrAAS4nztYIk1Pjqmigr0hRE4c7sSPYxNeSaLcud2SspzngTUR/wbEhgxz6y6qhN0KdWd3L/Wv8f6YnBn83Ekej3WZh41mU2QJ9ww5EQ4RzMX6Wd2mpyZUVUZ+enpyYuVyQXMV3IMG4dPT08KKUMejbD+h91AV0nhGpOz6kw2tVe4HUJqfqecHZ676VZxpPvpc7AhPg/jKRUjeEJweFN7jIeJYrHvYU4mR2AcgnYSzCGvyal9PLvuW1F7d0xcden7pDeQjVgAziDhaMR3EDoLfEHdJrOPkiHAGEUKIwMB8qPjypu8eh7g4jTnBffDlFePKbu2db71t87PT9uN/+KF6Q77z7W/ZX/zFX9n5edeuX3/RrdUODm3twpodgPGVyyJkOXPpvYIICgL6PFWNq2pamJ5Xnvjn+fUPxkIRw/didjWI92tkfnGNsrdFRJkIa9Y/64L9RxXUSWSt3ECVqS70YI1CKCBEBOVi/SKijqpvbM8mp6Y0F9mv5WBCZTKN16nIWVjQvMdCkOfBHsG98jtUi3EusmYl7BZZ1FR/wl7VfIa1uAVxqpjuN1XNSBvmnYsrnls//SpR+/Pf+Y0agbkm6nBXyuIjiMrDG2Z1UhDhSUHaK5UABsva2zRS34Zg9KScVWm/e9irj4SsTLzZKwc5qiU8NOk5IX9u+fHTO6Isr2TZdahhYFKHyXfzXMGukmcRDwDDDgxFg7WPPvzINja29H0O5kSVpsDKwV/vi+HKLtk5ZX0nxN+mpqt8jkqJUWVIvZmUyOWyLG44PLlXkurwxguVKO+p0lKNXUGBoStzimrmBcjlB2pHinDKEcdGhm1svGrdwrlNT4+rEXm32baqVa1SwGqiKKKiVO1ap4harmytbtH2j2t29+G6tbuMF59ZkLIFixJVsBS7VhnyJm4kpG5B4WWwjDlJXIA8Uq8kawquPdQfkTSqDJGxADAqFTUOalZVqSiJVUkj1RPJ5onqCgBZkib+zp85UREAWw565gsoEuGcSf8qooJAyK2fnKjQgUTQODKit1TgptJwDzDwzsV/0/sA+kGQq8j5HIARDiQOIgIJ9Vdpo16BtCBYcVBF5EVGVPSS7KyigqRaSlWSHMqWpWDFE7Ml1QOJBGX4ATJpHoYfqUixlp3sHyTFtitL8mbBgxUVcc8K8J5dTJECka+utHCwva/yCFC8D0z4OmddAcahDAzlwj8VUREBioP2riCWT3eynKIc0xXqJJCAsiSIdL/1YLaSrDGEmmQgSQ7m5wRDDqazVqQuTUBdzE1VdAHKAZolMkKBc1JtOAAfPZU9wIr5pcBLChxvOh6Apqu7+tUUEYT5dfZXRTSBz9dJHsTpGaUeFrEfxV4d7xnALOs+rmGQqMjfM8rnA3jnsyOIBkyIuRYBuKuaXKHLV05URNCpMyXdWFxnJFmMjff4YX/HZ9ctgVD8QRhQdYTKOvajfN16wkqSlppGpwA3APceQJhsf+K+KRHP+5RENYXvG2Wps3jWJNRY8lHfTsNrElX+U+JN4pIAdNZ3TowEqM6fkcR4RYj7qsa987lBVAQoGT8TSK4qwrD3coDQCVInXGMehgUMSSV7GOCalD0KxvtBf4CUbqXmlXGy/ZFfr/eACqIiP99iT3ZSJC/Y6jcFzonouLb8+cd8ifnEfYdiPAgJfhZ2fbFGeA8SMYJz3oPEMK/UkFo22V3lYzcYnMX8G7R87CUFKSEeTJLimQ2+X+jy83kd1Ubh8StCP8U1YevGwAdIz3vqNZSHywfcoy+qdvDGhaxQEstu5iGVvrTnyXoRAcDTRIVUg0ND9jvf++c2MTlt7dSImbN+d2dXnxUVFdicKWpTlWmy0/CLEBG9vbMjdWj0qGCseG6DFRXR5E8kBiBbmbNyOFW0eWWINwF15TWxBM9MsUkCI7Y3N0ipvR9OpeoWUMnuhTF+cPeO3f3sc6OPQ+rO8o8gKpz9V6WL/t/vOSp5B5917F/53hpr4Vl782CS/YuIijhnY83k7xd7nY5dLXLUpex1VAg58elVnR3F83y5QhiLgfEvERU6IyX6cZsKgbEJGEEFyaiomikqKgxv/SDg3ZIu4gHCBYGF2IxAVADuiKjoKLZv/xoVFbq/6AVVKdvpcc1aiILSveGRD4Gh/4pFe+vSm/b40YaqK6dn5uz09Ewg9/FRTaAaPYAuXVqzvf1dzacLF9bsMZapXeLYhtUbAJUte+31ryXLTV+nnP17hwfyXN/Z2ZdVG3tp7fjI2k2slahSmbLD/S27dGnFXrz6oqxcKmPDdrS7K4CXL1fkVlTJgIL9Rz/52EqlEalKaZSNKp4L1RlbKQtAFlm3uaVYVVVcmvtmDx7cs5sv3RBAPTY2YY8erdtQdcTm5+fUy2F+fsas40r6hblZzYPR8VE1AocswYpnaGhM74d6ut3GDqdhE1ROEJ826zakM4Y+eQXlJsvLi/LPZg5hjcHZR7UXStDq6LDsOgDdmHvEXI1aw06OT+yYqgm8uwHFVM1w5pXEVlClxvILl61xfKx8CW9uAF+WHjYx9BSQ3ctQVU1faQxNnMl8e/J43eqNpk1Oz9oXd+7Z53ceePUZlQOdtsBF1Pk8t5GRcVWoAFrJcol10e2IAIXWlOK4Xtc5A8gMSQ9BJHK9XJIFMoAfzwZ7K1VdTE5KRa6zm7MGVWvn3H7wvW/a6iL2tmXCuGYAACAASURBVFQemVWGh+3kuGGbGwe2sbEtK+IjLI6q7GkjVjvFvrhkb3/zbfvaqy/b8dGhQPqjxpmtvXjVPrh1y1YuX7aRiXFVTRAXDZdK9rMf/8haZy1r1t3SZXZmzL72ynVZa1mra0Plqp0cHKnRNRY2AGHYO9G4m8bHh0eAlDS4HhFQGI1rOe85KzwPpPIeYPbc6njtjw3LDgoi4crlK8rbqXAAnGUu6UwYG7Nbt27ZxbWLNjs9bZ9+9LFdeeFFkXU//+ADm5iY7uXgjC+g5+H+QbI28WpHrkmxMBY3Ah+dVMXrnmevuDJZ3ciiGIFUsmf2HJ/qsTl5uCMi0zmb+uZ4BQ1NtMdUgQC4PT09I5JEsWNWpenxvJ8H9I9YW7tgtdOGTgadecfHWqeI3thTDg4AqIdsdISG97sSC3IeY/3EnCeWBdSempx2BX+tZpMTE6pe4FpXl+bVhBh7qW+99XW7/+Ch8u1Lly/a/tGRVzAkp4NhYp9iSQSfzuPxce/boTw1GQGnqmDAdOY/PQui2jBiM1WDE0PKvtWtl7B8CvcAt/FOlruyGnUyIuIYwG4XFrjLA8+HvEnVmSmuDbKcMZMAtt22CxdWrQYR1qJZMP11HI8hDlBFwig2SfKEleKf+dWCIEmgrapEMgskqd9TdTvVA0PYapaLqo7jue3t7ajCbHx0RHsM192zWyo44SOl+zn7wJBNz8yKpNCeiYBTPSocKyCe1j5drdhp3QlNt8X2PhkhABWGcu79IPi7k0cu0OSzeeYiaeunT7lsuNjFAzuB9Sl/5PtBQvGzwC0iFuHPiK/BKPgKTIdrZ52yV3jO4/09IP+Y4HyOi4nchou56jGKA+SsF+IAyEv2TdlvWceuXX3BXrl5w06PvaE4DiCff/G59saV1TUB9B9+8JHs5D786CObnJjyXj0np4phqRQWJpfWeIiC2Qfi/I8YJr+/wIZiHDwe8mpHr3imMsatdYlj5RbQ8SqjyO0k5Og9j8hV3S2k19cvYVvYMMpSse2928CReN6ccaxLVYGnxeVkUlFnJARGiAHz+4jrD0FVnit+OX4MosLxV82MXq9Af0a9XP95M+1nherPv/ebPALLOqSc5VWinw5zFtbR4aESRk8YUo+GTGmWExWhaHeQMgGKyqexhGHDbNv01KQ2q8uXLmozUUkinnuo+1Wh4Iut2XUfdOKD6AWhZDGaBgHIJL9qQOODwwO7c/euPXr4xEE3eURzaLrFjzOnXbdJSPYNkQT1yuv0Wc7kxuEQCapAiQ5K2nLPG5BDjrKtfjKFBzclYl4SKHZcTKzbuRBAcHhCDMBYE9RInZsUiO2zhpj/ielRGx2rqIS4SR+DQtlGS5QrYnlhVqp0rFDh8O5as1W0lpVEVNy5/8RaEBUlwCV+XHAmWECGK/DdYz35MFK+XqkoUHKgvaWDXVYPgCayWknlfsmagjkh8Cg101VAIq9IT1QbeNy6U7+TEsZhCEHhfSrY5FFJY/0UoFpPcZoCmigvjTWVA0bxva8mKjqwV/iLqdw+Jyp6n5cUeMyFyekpzUeqGMKzPgKrsCmpDpEYtW13FyUa1SkEHg4qcmLocGd8aA4nD/1YJ33LAuYP1k8koQKrUfScexO4qKggmaOiAoUXgQXMuj4jleqyFhh3WT8lYDDGoweiOZOmb8fajMPvFxEVz9q/9J4enoqoyIE6KSlSlQLkgD4vgVgoEfvPrt/oeRCkGfz3V+2h8bn+/Ji70nr6r2NvhgoG8EoJDT6bDv6zDzlBkSqyBLywMPr2NTnAlM+zPDjS3qFP7TfQ5ucAvQqCAHCSzUbvHpK9jGdSqVdE1qC4RwhI++fPKicp+F48t/z+A9gaBMPyACd+JwCuZxEVAcqqQiGR0Lwn+1FUW/ke6M893tM9MzNlR+q3EkRHKNmZ1/EZQdzE6wS0p8/Mfxbq7ngvr6hwEMyB3q7bimEzKHLQwf7ePp41os3JEY1lnBfRkyIsUzKiwisMst4eqWk418i9QDSTYI4Ojyhgr5Yq6ifBnoD1E0RFJIC8JipjcqCR8WG+Rnk6Y5sD+RHMqkqj2VQiFWPPezIO/QoVt8fyag2u3Qn3SAh5b2+I7s1WSUYgHbkuAON4toyP+iTofVyJx2eHNUZ8blxnECv5eonEKK7ViTJvZBq/nycVPfAx2bhFxQm/Q8KXB/WRlAXxFWPH9xknEk7ulbHivyBUSHxjnQWwofmW9SrIz5jY7+Me4meDSUSsR48rvF9Nvl/4evaeMrGGgihxu7FklZOuw/dRB8jDBo5/+mtobnjmQJ3ACa+OqTda3myQfUnka9oOQ3WWCN0eGUU8Vq7YxYsX7Rtvf8tfW6RCAQudru3u7PQqKgQuYO2R9qvcYoBPAcwDVGV8IeJ6zbQz6yfWJT8L26ggKnLrJ4QkuvdUGghRQczEGpN9qOzSzHZpXGtOmjEGgI9OVDDfzU4OD+zDn70vkFA18cn66ZdVVGjfSER/fl7GfpL/OXg25WdXvEfswTmJkL8uPz/d2qFvKaWeL+lZ5iRqXFd+BniFXn8PdTED5xqHDmIW9w2nuoIv2X0mOwpiHPYuelQI8EjWT3H+KLGOprSpokJm41lFhSp0UeqX+8R7fn2KBRF+QFS4G34iKryJLtcI8f/0ePhI5WeVAzX9MaIv3hniIAhXiIq8ogIbu1LJ3rjwun3x+R1bWr1ga2uXpJLFH5u5BvDHXLvywiVbX38iwObixUt2dFRTjxaU/xJAdFtqpEyTWq5e4pDGqWwp6NHz2We3rVoZUdxGjIb1U7nUtYW5aauUyXWa9sorN611fmazi7OqWKidHHk1myqJinZwdGz10zP78XufW60GeXJJTZSZ8yurFwSqIIx5sr4hUgkf8bGJca/Uk7XRkG1urdu1a1clDKHR5pPHNOgcklp5B4B0YkTknZ2fK9/i/OL+aGhMpcnjR1siFNg/3bsc8sXUUwErNfe/x0Mfr3xylTM1556cmpBlC1Y4Oktoulyv6XwBDAU8pbID0Rs5C3OAvWx/f09+5AKhOgWd5RBXrFMAdEBWemi49ZJXZQE+j9PTQz2BihrvsdER9QZhnyJvpIl4gcpGbrVtAsPXt/YcIKo6eWLGuYuFa93BzjYkMPY7bhuGqIrYOuIq/sSGCFWsnxn9mNGVxSdu5ZvWHAracypJil2rFs/tzddu2tQ4ivodzSUaZsueuFiyg/1D2Zusb27b5taO3b+/7qKvSknA+ne++11bWl627c1Nu33/gV188aqdts7toy++sFdee1XrmeqD93/yI60FQsirL1yzxflFGx+r2OgQFl6n1ml17ejw2A4PjqxRx2rkxJ5sbusZlIeG7fD4RNYlTkR6Hhc9uNy+xG1TFaulOAmRA1UbgPuMCQA7anTIMQkv1BAWMZz3VQPAe+O11+xv//pvVNEyN79gP3vvfYG8in14blRPFgouOJCK2mMcEVsnNc0xlNABZAO2c208R4nOyFMEcPq1sn8hvOPLLSDd0ks5blJoK+dMZyXnDYAxeTnv57ZjiaBOlqnK2VqIB72hfadb0LpknLAF5jrp2UDUg3pavZQqZa1hxSfFoh0f0VAXspFm4TX/O3Y/dSxlFqzeqGler60sa94dHZ7Y9asXJSI4Pqnb6oVFtw5mjBN5zrWCz4B/8Ay5V8W+3RSzJ2eLUGNHhMpzJIdVn1GRdqnXVy93dAWEekYotvT50MsVkhgrqo3YkyTCQbCZqveIxXo5aHJNiLUdez/WaYwr57bOdyqgWm7lzZ6H2px4ozLsc4AvWeQSk0NYJjtN2bPpGhBPArKnOE/X3LLJyXFbXJjX68A7aDIOOaWKZayGhIG5iJD30JlpZjMzs7a/f5TI3YoIb+yOyPsApt3uqqDqHASdyhMkPPOeaxACYD3ML6o3uK4g3ORcgYL+nIqaMRFZ0V/CRQopx5bY12PNwDB4Pxcb9e0X+7mENx6XaDNqdoOkw9a2UlHMxmcQb7HmWY9hkUZs4dfoOILndA6Oh92X7tM6QgbAK6hW0flXKqrSnLyEeUisRhxCZRsEHvfA+Qy5x/VRiY6lIZ/fSjEKz4D9HqiOuDfPNxVzD9jU5jGCctVOEmBhlZ6EYspr1XyaPKeivUMWbwiz9DnkVo4bhLhY+1LmoML9Y4GIOwiCBvVurQ7bxKRX2blg10Ut0YsEOyjHNz1P0/yNCpkUHAbxFDlQnts/jZFE7w1wpYRMxoMhdio7Ya619ZyoGAzZn//7N30E1lBZJiUvwZ0CQLzAaYy0f+AARlpcUj+IqfeF8lTC5ll4z09di1LBDg0ZK3blyiW7fu2qgymFgnpReJNQf50YeQ4WSrFQXnUIMNzOCWseL5ljg/TkhYNia3vbHj7CQ3Zdap0C/prazLxsOGxDkiCxv7GnBlpxcPL5UV0htUAA0CV8sT0J4nrUeCk1SHVNI1Ubbv/hzau9ITcHmPyZUwDIxuuBU1JLp8CXigfUJ/g30/Sa0u9ihQPh2GZnJmwM1rrZskITWwP6dNBfAfifxmP4sZZwKre9E4iKx3bepgR+SM0/ISp6PTQ4d0qmChmeX6g1Sdaipwjfk2oxBRVSWifwJJhiNnQvb6SSwJUwnlh7403K5qOEkOAfggRiogVJwfPsAvC3vtSjIsCwHMyKdfXrEBUKUBJRUcdnHa/RVFERh7yS+IoD2BAVeFdCrUSSLKuVpIzmNWps3KXEedtOTupexh52CAIe3c+S4ITkkwAwDnkFHPJgLcnPV/ZLwtc7XkKKLVV1SN+DWHny+JEark1NTSqxU0PW1MOEaiIOzyAqcgC5l/QPNOvMgXiv0/31diu9b4+oeFafCm41NaI1mqU1VPXUf3b/OKJiEMxQgqE55GXNkKtSXqnJPWoKJ8f44mcQFXqPZLNCcBWVCYPvHQBTDlRqjJN3OLZxAaJHEqQ5BRGRbjiA4h5wk1lmBbAqQkCkHGmDJwhhBwShSQLM19PglP871kIe7MS8zn8eQWtOdrgfvAeejKOUTSoPjz4SDo5HoJTv7XGN+WdwLdyHe7EOJ4s4rOdKUiPm8zPuRySRGoE56RN/BoCvfTT1vfC92T1pfW/xccOKjH0H0JPkNZ/jEchGFUKs6Zy0GQSilYSKgE3VFGru7KqkCIr5DIhqkZvjE55UFYrGHsM1Y/sEiByVakE6xbjFeoj7zImcPPgOIiIAKc7j/Jnzc09u8Ccl8PX9WGR4CoRdEeVziKSYv2PTgTqVIJ5zlqA2Eh2tlXT+x1iwb5LEDCZC7HF5ghTXxlgFkRE9TnjfwXGP5x2v4zUxJhHE697TGsnVeLkiLQBwXiOwLPXZcJ9pjyWURKbKhPgziLFBYoHvc60xhvkuGSRD3Eusqfh3/szyNRuEkapTRbj1VfpBQkgFxbqUSs5jhLhn/u6e2Q2poWmUC8h5fk4T2jM90zaxSrbnx304yOvJrq5TNplVe/vtt2U/wxHZLbkNmFdU9ImKYUQWEhVEDx5XSEbcRXLv6u9xjbHUz0lderC/p89Tk/tEVPAzwIbDo30dQd6jgrnbVwySkaJ0VO8mrIWyJul7uztWLjhZ6ESFExZqmAtBfN60n/3Dj+SNXCDx/BWtnzQHBioSB/tSDO4VMS8G497Yb/kzPKkH97/B1+bvIaIiVcbE3Hzq55lNX28Pjspfeb4H4e0Ehc89J5UhFSKeQRQzMTWVGrxq13BBUOoHx3XkRIXuPwEe7NvExhAVUiHSNC3N1/68h4fwCq9ilwoMoGqz+umJYkbAWIgK8gePt/uNL3mvEArl51Y8J8bnvN60Zr2uOJbrkm8/IHCKq7/70ndtY3NbMTo2TfQuePj4sWKtkeqwLMv++e9+T/Go1JCtth0fnUohjb/+k/V1edD/7vd+x62QDg7t5z9/X8TK1RvXRRBSuTA87LkLFlJT4yNqtrm0MGMHOzs2Mlq1ay9etpdevamGmIc7WzY3OyOC4fi4ZlPTM1aqjtiTR+t264vHdnTSsIXFBVnoMMf9ur2iSY6DxaLduXvHVi9ckELbCduOHRzs2sLCggRQVDdsbuxIKYonONVL9KgALKWZ8srSgh3Xjn28tdeY7e0DFqXefGWIMnK1c7t4Ydn2dna8cSpVn+dN2RrJ/mOINViUTcvc3KwahWIXSxNkqgawokHdTSXC6vKKFVreX409fXRi0k7PGra7vWOtBnGGK7KxokGhy5/Mo7m5eVteWdEZzN6keCT12wGgv3XrE1tdXrbFlRWrHWGnM6qzd2t3z2g6DJh7dt6xJ+s79tkXd1SFVigSo3szXAGaVJUDtstKhp97w29XHvtaunT5srH3ACKS05EXqdpidES9FkaGsB2qqkcG16o5ed6woXLXvv8779hotWC3P79lX3/zdbv/4L698urLVhoppz46ZqfYde3siVjZ2T3QHDw+bNpLr9ywf/bd31Yc/ejJE2sXS3bl2jX76PZt7WyLywv28Ucf2uHetl1YWrbXX31DvfPKhYp6+dQO93U2bGxuWfO8Y7t7B7a9e2i7e4dWqkAseZ+Mw+OaCA9TZYmf6wC/3AsxBvOK8XG3BYc8tWa6busLGRCCAnIggN+La2u2uroi8J33xM6Z3J+1ynmxu38g8g21OeQaew1xOqJDeeUjkCPGabVkhzQzPS0QU574qbKTa4MUi7hJWF0CVAEZ/Tl6dX/EBlw/e4usa8ol7wmQ+q0R67CO+ByPkbxJcLhG+L7kIzAyOizrFtbq0vKSroP9vnZaV7+Sufk5x1LKFdvc3LDjY7d7Ig4DyFQPjsaZsAos+Nh/Do6wjptQRQvXcnFtxY4ODkUsXVpdEqkIFoPVqapc2E+bTTUbp4qC91ND5GSzxL7BvPRzxIU+6ocnwZVXW/LcRBTSD49YqTqkqhhEEADqfBY9GFQtTNUqlnKyN+bfTlJBVPJ8AZ15H0SO6v2ZqmqiipQclvHWNaTG5OHeANFFvwpcNZgf87PzikWYdxubWICN6JqpcpAdUCKOIDAVNw57pU/EdbJ7SyQnlT78HUyFtU7vTwiLLz77XETyyvKKPYLUXF/Xs5+cnBZArtik0Na+wr66v39gpzWqO+gRxH7lwh9vZlwRScYa4RnFeeb3jp3dqPdyLYIjQLa4VSnXq95oiB65tuFhERWcW553+B7kOZvbP+ne0hjw/nmsGnFK5HiKSSUm9dcrXyIvG3bLTPImron5K+EBdlqyh3I7p2horjhVfSJS3pDyCr6PgAail7nAeSfLos65cm4wH0hKKgSHhkdFjnONzCm329pQxZustMnneD9Vy3M+uRBDBLIqhJ+uGokxiJwjxifGwM9Mz3+Yb54Peb9B2UlBMLEHRp9G8r7Ub8t70/QrS3le2hsRcUM8jYxoDXN9iI7DoSR660UPPdls9XJIr8zI89TIz+IeIueOe8h/t5+LCHFN1S1PExWKZNUTNwkcnxMVeQr3/O//O4zAaqGkA1p9JRJzTgMnFmEA12pYJUAAP0JvrqxF0VMDOrAjYEa9LVwVw+E9OzNtr7x0UxvhRx99qI2Cg21udi6VmiKA94Ut5rPTsga2H4nA4GT25q4dlf1xcHHAExzQnIiknc1taBi/0SEv/cX2qexVAuxIkdyFis1BydSYmc03MaEc4iodTB7JqvhIfnJcM+Pg3ryu/uJ6FdThbaomy17+FQHTae1E6pKhEUAGKisImJOdFeBOqkggsF9cnNdBurA4a8USVggN69DMqtuxEQgYmkPRgKnYsvMOiVZJREW3WFFFxRcQFR1UrMPWpSY+kTVKxklEkvdqlI2hfuKwQwHvhyDl2h7ECLCidFr9KvyeIGIgkdyOw+3BGFcpJ0pFbwLerPcS9U7XD2iA7HYH1QpkBUTU09ZPuaI4QKF8XUXinifwuQJXm3uqJFAgxHViFZNsJAatn+TRnpppQ1SgBnIiLBqJuco8lMBDFRRhXdvZ3lHZsVh+LBayhqEistodKS5cEdxXueZEhdumedNMBTZ4qQK64KF6UlNFBX1bOAy3t7e0VkiAeA09RAi+jvcPemqg/GDT4TZAVDCOvUMvlY/+OnuWxuSXEhUeTHCgqwF4Kjd1oO2flqhgPgF4AGCrkmLEbV+8aTaECaXANGIFMHcwQ2PQexxeiTQIVAbgkoNJMR/YC1rsP5mKNcB+TTvn6RxkyVT9PnYEXU4wBKgf4LeSCIDm1PwtAOYAh3PQM64rXwvPutYAnaKCIALnuC4+wxXnXXmiRlVMDgzH5waonIPt8T4x72QHUKfpl6t7+C8qBri+XIWVXwNjEdcaa01VaCl59FJjL7knViURCBuj1jkVTU23CEyenIMqFZ97EOJUyHn1QADH+e8qeUukiVtu6ZV+1ijZ6JMVVNRAwExPTSkRxWKONcvZBRjSVPLi+0Y80/wztf+nigo1GpZdYJ98is/qEVopMQ8wIPZGxkjncdV7TfSAcwC7ogP/vh95I0MfV0j2U+3h/BywKQfcgyjj7uPeoyrlacDVvXAHQdh4lv1kod/fpBc89xoKMy/6Y8V1MB5xDsS48/l5EppbM3EPMd/iMyV06HQUy/BFYsh/MdfysyW/zpgrvXjmGXtoJBJRMRRzOdZXrAPNubQO+B2NdfKI1rwTaOB7ovqZJLWcQBdIf1VgdQWyxP4BqKp7UKyFgMMr91BZngPWDhAVQc75uHviQvINUPid73xXID/vZZXkE/4MouKs5dV8/DdYRcV5j0AkJyq4VuYkRAV/j2qLqILpExVYSvR7VPSYc9ZhqhaKKq84twALUSrnRIV6VKjZIeFF297/yU/t+GAPh8tfuaIiAPDcOvGpszF7VoNnZlxbfD/WuZ8j0ZC3X4nW278zYuSps1kiAuwZ/aCK+fnM8yid6X79JOMJ2HBZqJMDIt3cmkAVzexLxObVqhT3kEgeG7sCNPb4eI4Sa0TFRzpDo0+cExV4afvemu/lmrMl98qmoqLQ9cb3WD9RVQtIaEUnmDxeedpWK19X8Xftz5rMTxMV6onGWGRExTvX3xHgOzExpTkO2Pfg0SOrAiqXKra5sWHf/c67trO7LXU0FQVUVBwd1qR+BpCj2uza9Rft4b17toh1zOmp7R0duL/06Lg9Wd+UlZAAyuNjmxzHnqRpU1PjNjMxJvux2dlJa9RP7Fvvvi3b073Nda9kmV+ynScbGoOj4xP7+NYDO28VbERipSM9F6pdiBkfPHxg2zu7try0ZOsbG3b5Mj03Dl393jm3k9qxgGH2GBrrvvfeB7a0tCoFL6DRyEjVG9KendnN61dtfXPDbr50XVUFjx9v2J27j+zSxUupB1Hbpqcn7PBg1y6trcoWiSpiqoRdIOPN6lV50Gro/BgfHxGZMzs/K4AWggrgkHlM1UCHJr7Do7Jn5L5QwhMzA+wd7B7a/t6BgNkKtkIAZAlQ4pxiv0JARB8AV2jTY6CmOJ0cAoBsZ2tL3vf8DPsnevnUz5o2OztvR7WGNc669tOfvq9GrQcnNQFigGasT/ZZ5rHyn3P3tx8ZGRLwypmKFQvkET13+Fyt77Svo6SHqKUHIKQQNnqsAVFu5w1rnh7Zm6/esIXZcfvw/ffsla+9ZH/6p//d/t2//741zo5sambKRqenrADIp4r1gj18+MQePd6wjfUd9dN4+xvftuuvvmYfv/ee3Xv0yEYnp+1bv/Vb9l/+23+T9dP42Ih97eWXbHJsTPF5uYitScF2Hj+x2tGhHRyf2Ob2jnUKJdvY3rFiBQ94mrSOKRZg6QMCt85pRE3lzLnslqnAYO0yV8ljVMWSbLZEVKr/IPZ8Tm6o8mWoajViSVUfuZ3S9Rs3bHbG+xB2WufypWcebO/uyqtePUjM1yd5vgiwEpjArPch63bt4OjQrYiwcBkaEckAsE0+zReEgeMMbgXrvRQhxeh1BJCNDR4VFd7vxJsXuyCNOUN8ybxkf9na2vKm06lXp5+dvn/r/s1sdmZK8xyAnwbL83Pztre3lxwFCmqSzNnGnOY6qXpS35B2W/0NIScg9RCy8R6I0QC8D4+ORMhQpQIxsLK8ZEcHB6raATuhEoMvCEx2vEazZdXhqvYzgmIXNrn1IqGFeiY0Uo8B8twCOIHjFDVIn3IpNVQu2tHJkdY/YgP1eohqleEhF8B0unai6iV6bgw7OAvwrhiX3japf0vCamQHJJGBjx1j7ZiI9xSTSIaeIDhFVKpOdpxCmJV1fasrq/pcrv8EEuToSJVk+Pnr/SCBcNxonGmv4b3oKwK4TKzH+5LzYbcloYUcQiBLyzY+7sTXZ598Yi+/fLNnBfbo0WN9ztAIa8NdMCBOITOIMe7cuSvLJ4QRnK3nqYrD3TUgNQoC7UNgwprwShSPWVxU5E4VzGGRNiIG3A6I2Ih5yJ8hIPOEOvIWP2sQsUVs4MIqr3KJGDSPGcJiNH7G77FMWIN8LmvDe6kiTnOiAkzH4wbHOxxM916ynk94Tw5+JnEmogMFtDTtXrXD/V0bHxmWAJlnBFEK3jU5OSOigkoj5gafubtHhaGPH9dE/gTBLawqCSr5g72afUdYW8oZI0+O3C3yt148pSZZTlipRyn3oaowF1qIJNLzqAirYF8glvH3S9ZQqfk2z4l78Nd4JQq9XcDBWBOsYZ13Bwdu09rxZ876YDwhkNX7N62HINR6oq60RuL7kSvFvT0dd0aFqfcHjjw9HEi4piBAnldUDEbsz//9Gz8C03UvqQtg2qsnCgLsA7RmUeSgU3giO1GR6suSBMHZPTxtS652pjkQavoWJVAoYr0eQ/65iW1mUUvBk7zgqUF2oiKlsl504Qs02QzxFxTq3kTQfcwdQIFEIIkleT5z+yd5JvpmLYDGt3z9GeBDbBJsKgRBkciyWVHeKRA0KcCCAIlx0sbCnt1uq1wRQFlK+G5HzZrVcIpqFR2uvuHowCUYVOVDWyXTBHokgcPDEAinNlIp2+rCvI3jI1spWxsbiAJNZupzbAAAIABJREFU6UrWlMd9GS8o2z+p2Rf3HomoKJU5CM1azbYHo2zWbLbW0edxre6l2NZhwSEVQBPEiYLuVC3B671hHACJ2xpx/Qruk60OQS5l5f7982RDwHh4BQUHHIGt/o0nv7n1E1/9Q4eDsg8K5osqB2fjMM7L6HoHdFICAFa0m+dfIioiIWc+cDjxTCYmJxV84vEcYxAHogNO2GdBzjWlEiOJKpeHREQBxvA8ZUMh5ZGXV+N1HIpuHSaqqCirsZJINgK5csm9uFU6WRVhRZIEUUFAjFINywspHJh5KA7OmvJNPtylmbYH6HHvPVB9AGSLe4rreBaR8Ys2MAfL+s20/XN8/vrflYo4IaFS0jMFh/H1pevLPmwQ7HnWdfTuK4E3/u+ODQ17YCoSB8BCTd5RfeDD7gCW7zOJwwrfSD3npy2cBq81/Mn9+aN2LlhTzec9EOGrr9RyxakaAqZENt7P7w/FniuTw04nDyjJMQLYD2CGPwPw7gUjsbcO/Jl/VsyHuI4A52MOeBDqIHYAwAFG86erafpkXYDqsed5kEpVg69TElLeK9Qk3GMAzgGCBzgczzrukevOP08WQan5W++Zi6iAxKYfDH7EBND0gSH4Yy/1pt4RqAawGp8RiVKAiPFngM6auSlw5jWeRLGm3FJIzfJSEiyv/iH61eA9PCo1FNVDqiAi2Whgz+NzgKSD95PaKoHVQcDkRAVzKJ51jFMEqFFRwXsHcZETFX4WRymzW+Do2Savds5eB88bKj8H2GbvInB2Mt5tmXQOJaIs9lRViCT7pXwOxVyLmCD2gGclSvGzIMBi7OP9omoi5gmVZUNqhOqgqidQXt0Tz5XfVc8D1lvZySDGyysa/GyPniBUVvD7SsCzJut5PBPzJtZHJAuxbntms+nGQ/3kvR/8WccZxs8gSPzsHCCByslnO8Uzg9UVzHvO1kheeE9AB12Pqu9cXecKZN9TWBMINE7won4qmvFEL+wd6Q/G3/nvhWvX7NVXX3eVWqFsXVkEeUXF3u6u9lDONCoqWF85USH+hOpXM6mm6VGB3zbrgTHmnpkzJHFSno7ggwxI6QINknA10y6a7AC4Zwjc7KBQ02bGT3uRSv99fPtERVVnLSQFoDFAvCwRWud266OPbZdeFtrb3eCiLxXof0x+5vxyosLtQr/qXMr33pjfvD+Al1eDPZuo0NqQ9VO/R4w3j/Q+UnE+5OdEvn/m+5vHRqjOPa720y5IWd/rARfVJLVY1DPBtsfnGnOrf5YHIcWzcmIsXUs684ia2Q8RuGDjiSCAteBEamro3SMqsPwBWHHhT6N2LDsN7U+JYPI9wu1eB8+xfA2J4OO2iPGzioqcqPCG2kV7+8Vv2p07923t0iWr1xrWlGK1LfGSKj27BXv9jVdF8iIKevDgkd2/+1AWQVtbOzYxMW5nZ3V7662v22effGqzk5NS3u7u76hHQqFUtvv3H2v9ENMBZNfrJ7a0NKe53Wk2DWHL116+bpcvAfi7ynR8alL9W7qtrk1MTdtZvWmbm9v29//zAwFkCGboXUClArY/KHuJ9/YPDvTMdnZ2bWZu1r3EpTBFkX8ikQ3PDfJ+c3PHJsanBNoBuiv2ltipaRfXLoj8BIxG1Y6i/snjLVU3OSDGecXz7NowlopUHLQBY0bs9KSuBtfbW5vqXdHpnFmxxB5MjleQjQrCmsnJCZuZm/GKp2rVDnZ27XB7T/Ettk6jUyibyUWwmBqSepu9RKB1mv/ka/QXkQVL0Rsii5ivN1RpgY979HBTPzRsqSZQ7Q7pvvYODgUYzy0s29b2od27d18CguMaFV01zQOqCvhiXgC+BjjpOYBXKCIior8Vn6FeF9jhqrrDq84BHBl3qeCpZih5ZXWp3bKxSsG+8cYr9sLFZfu7v/kbe+fdt+2P//gv7f/8v37ffv6zn9rqhSWbmZvWnJ6YnnCCsuh2TQf7x3b79gMrlar2xpvfUE+Tjz/+2EbGJ+3StWv2+Z3btkRTYIQb7aZdvnjRGvWmrMtqx6fWrJ/Z4d6B7R8d2oma0+IMVdB/LQpTiiWrlrEsw8YY+xPmRFVgOGOIPQsANGp/fle2JakJLfeOQrxeB3yPKi13OSAfZM1SpaDYVZXO9H2YtqWFeWEAAL2Az3fv3VNFH2cP1skhqiD/0V6S+pKhaGeMvKdIqQeQU5mApUrsufKKTxZGgIW9uCQJRgBiObuC1IjcFmU3TZzZf2RVVirpuYb1aexBOrYljirYCv0MsQY6d3tnfp/eH9zz5NSk7M729vdsZWWlJyLxOeYkBDHK7s6+Nycfn9D3EFxScSULqXrDXnzhBdvf25VF0eLCgkBQ4ssVKlXooUNFxdmZqim6ynscgzk9xfIK8qZvR6ncU7k8e+CZiF0Ab8UuVGvqufkezfcZP85fxVd6rucaa6pnmO+s1cg9yaEbdW9uz3OSIIOeLwho1MPz1IH8ZL3qBIaXpri9U0mEAvgC5DliM+JVMAkIEHJsVZqmKgz1K1ClPMQcfYO8dwN/Kr5Gm9nm84dEaPLLfA59KUaHh7RuuM/N9XW7fGlN/WUAz0+Oa0nMNOQNxJVzNGRTRu+fTz+9ZY0G5EzZmmfnij8gKzgLiUPYq6L5dMSQ0ew64iJia3fboB8FlRn0fYGocBswBL2yoUqW0owB9+qVFSnPzkRNEbf3sQqvBudzXeCVBFAJy4v4AbJVdm9JgMKxCrnDHPBG3557xtpywVg/1yfe4JqpzHCBGvZvY3bl0kXtISdHB7J3Zz7SPwgsbGFxWST01s6uxh9bJCqqFOuBJ8kNwWNarV1NTa/y5HmG8Cbi9bi3PL7K82QsQXUPsoLGUmxYCEbkuhFrxHNgz5L9GFhMEmPHe0flilfHkO96vEOFM31pwAT5PkQg5BoXL9cSSCqRb14d3u9Jl4ST4ayRKi0iV438L/KiPAb0CuQk/hwkKoRN9kVrz4mKZ4btz7/5mzwCU3VXIoRHpzaGpOyLhthizzkM3DSu13hJJZcq409NiNVAJryHk2oqqcSUa5A04Y2oRIlmt55bAdS7BUJYraSmtFG1kZJx50S8UZOfgL5xOHnhbC9KIHnqyvqp3/CPX5dljEAxJyuwufKElTzIK0q4V6lHUoNTDnMlB0mFwe8TUPOnSr1kFUUpnwNPbHYqPwWM5l4reMf5ITs83FcNA07LXiOBsBxSBExnTUpWKaUsWanbsqXZaZvGU3GoqqRofHLMgVNA0E7RGq0OrQ3tJ+9/aJVhNk2aosMCOwgugoFrrXpviVB4qj9GpawEzhUSFakafVg9GNNz8sxawUOQOqGUV/BCcApYLQUmr+/KGoBgjOSHwNMrKhJZ8QzrJ8YtVxTnLLlvzskiLAHkOSPdA8MToC9lfaebPB9RhFalhCbRVTUF8zt5Gk/NTIslryRPcD5LYFaoGhPwgWKI4J5xQb1GQ1ACKVQFkWZzEAJW+SHcb5LsQcqQzc8vpAZkrgI8T6oLAZt4bR8fu0psfMymZiakQmIeqY9bqqgg+Ds+2E+rwZdAHNIKRhLwMLgfCcLIDjLmdn4ICpTIXvT0AZmrHjkMk50SjTJZM6lSB0UwwQsetaEICVIjByJ6H/MM5XLv97L2pQFnSStaLNjoGLZqKJBpauVN2RhjNbXWGvXgXf8lmyFf+06oRDAQZJKDOSg93RPeQUju0fcTeYCz3gQYsq+4tY7PSa8qI+kLlXfM1Qj6AnTNA6UY30GiIn+eg3M8fyYCb7JnH3/vkRH4iibyWcqopO6JACxU+qFejvcLcDIIxLinAGAj4A6LlAgio/lygLkxJ/M1zbUFeB+q+QDyBbakCoYAs2WjlNnUhXo3lEsABmEHpAQ1wz0jwAzwLT4n9hl+HiodnktcG8lDKPkFYLPHylqlK3JsZNQJSgAvytE5awCVzwRoePNANZxLIAt/8n6UxPN5QVTIGrCKNYsrhQbJFo2bAlySIOzkvLyd/2LeevM+73fBfcmOSn6yntg0GvRscCAHwEP70/Fp8vr3ZxFfeUWFn2+NnhIuB0nj8yMhi+fP+MUcyvcersP9ev0eY17E64I44PN5nrKDSWs2SI58fEKRx/UFUcZnO5ji4HoA5CT4vG80Ag2CTntB6osVazXICu1nvbXd3xHzJCnUaKrUSVWFvCfXSdLZSwITSaUqF0CAVMYelVmqqEgJvnoppSoR/g4440SNqxPjDPQ//TwgcT+u1ez0zAlvwEfwaoG2bCxyV+IbRRsZm7A3v/FNm5qeTQA19+nqxrB+iuaiQzQizMjcILB6JFrzTNWFGmfm+/i4lp4qKo6OdM5wpsX65HU8G8ijqITLE7He3EmEUuwlMVdQrVJPGs8yer9IPUYM1T63Jw8f2cM7d6yr+MX3xoDtn56P2SYxcEjGPO+NdYoLB8/S2GvzMy32S86RRqvZJ+tJ8rODFeLoq75Q9/fsLQbWk/dJ6r82SLK45gAo4trzdRaVRgAB01PTahBKDMieQBwS9xMkduw3cX7FueNrFsFN3dotYkMHyDwRT6IAKYFS0kyPCvn4F63RBIRhDyR36O87ueghFE856RPntvy5AQnOWnaG8jQJl4jUACSokOX6Xll+xW59+rmtrl1yYKnZlt0Q57P2oWbLXn7lpo2OcnZU7fbtO3ZyXBfoUCJmTmD19373t+yD9963uYlp2XMeYFuGCrVYVnNbLLMAxFHess8SkwCGnZMXtM/tlZeu2dwM1QbTagRf29+z6blZfYbEU4WK7ewd2Cef3aOmUkIigCr2NClK1az11A4PjyWk+eKLu3b9xlW7f/++TYxPys+en9248YLvrW2zJ0+21KAX0GT/YN+Wl+etVOhYsdO1ixcvCGDGIgvQ8+ysZTvb+wLiZBtUYX05YTE1Pio9C1URw0NUipvU47UTRDgn6rcxOYU1TM3GxkdU9c26o8ny6oVVCbNQ0zPVmzQdZtxl5dex6uiIdUtUgEzJQkXgosjYZL1bcosNAWKoUdM+CCBKzE0uwZSt12pSwUtcN1SVTRMA3P2Hj1SJfOHCJStXR2StRP8omoefNpr28NETERRgYuqnMeTNeokrsY5jsTKegEyTsubxfIZNk3keoHAAYcNjiBK8KS7zsmwt6zYb9u4337AXLizbD//+7+w7v/Wu/Yf/8Gf27/7tv7CPfv6xvfzSdZucGrXbdz63S1cuympsfon+dWXr0r/gtGk7O3sSZFy9esP+xw//QaTDHjZDnY59+51v2fzcjAhcPpOqSRTJJycN21jHnrYmwrOJEI0ztVSwk1NvDkz1/BiWS6f0eWFdNmxsatyFddZV1Qv7LHbEfHEGcXaRv9A/gedCHAEgTr4McczzFQFN5SYAswBYJ70B7wCuOTPx+4eo2NjaVm8KKorIKb2qnHXhVRB8QXSpQfWQxzbsI6wbWX1SDZPseWUbldT4fP7h4YEIEIG2nJ1JVKDm6yLT3aaUdUZ+GjEJ4GnExowF+43igDRH+RxyW0he5gCxH+QfFlfYO9FPYmFhTs9nZ3vXFhfnlAsiLlhdXbLaCXvEqIB5wGqIfprEY49DpQX3xT1xj1euXFZ1F6QRFmdUE7A3zM7NaR0x5/ldxln2dwg7VDWCNfRIsnTltHBbSVf1p95z4BRqku6EjpwsCpCNY1oPAr6JoQDTQzBCfxCB654/9ePlql4Tdk56TopnqNyrWOP01PuIJittPs+FkS4K5DqoTubIoOKBeBg8RBUVZ2eyCWJf57lOY7cjvKOtKisqvLD041pm5+cUh+B24JUyXVtcWHT1fLstuz+6eUnMCgZxfm4rK8ta85yDDx8+8kqWlTUXYNBrpHsu4glweGNjS2QUAguqkegzI+KrTUXOsAh9Xzduoxg5T1iEh1AG0SfzL3I0ETJYa501tWeyx9GU23OV1JBcz8nPfcayR6omgZGEocm6UfFQwi8ixvB+sQmPU2xLxTtEbb+3HecMZz8YB2PPGnQxl6NtgO16bjQqDxt4ERreSJtKlRcuX9L+MDM1ITyL+3KCrWlLK6t6dlRYgG9BjICRaN6ee98q1p8+U2vdK6R0IqR8PI/NIl55Vr6RkDytdX8WYFAQ455nMScijoUopIKKvYF7AVthrkHoB+EpUq9QlH2ba1YQ3TRsaKQqohG8g3iXZ6e/p+oPj+1T3x/dlz+RHlYV/tPpQcUzHIwN89xLosdU/c+Z4zaZCItxkwAD9XvT835u/fSVcfbzH/yGjsB0wxXzAkaSdUWwqtqQk0pQh1gqidRGIODES8SiCafKY501cDUzGwPJDCCfV6YnlTObUWIXE4joAYkDHpQr9jzXkvpMzZ0IINRYiC3Sm6p6Ux4Utw7Qe9mhAySo9tiEvJzNwQA1Xjpv6jqc5a6p3JrqD22aKkFLiuwENmgDa9S9BGxoyNWcNP6EvOmptX0C8HqBbajPZJlVVZKj0jmxrd6kDKJCBysKZW1m7i/M9dC0jiSj1G3bwvSEzYyPWIkS/m7LqpTts8krsTcrDQ3ZzuGhffrZHRsaG7dOxxsK0UxNlRApuIxmOwKoUBtA2qRKgFB10xzWAzYHc0gOCWa8cV3fz95JDBJVL3HTgd1F5YmXKxUERWu2CGLaqhCBsaZcvaMmnV+uqIiENADUnJiIDT7f5L+KqICdUfCZERWQNUODRAWNqEolqdQgKtAvxPszz0P9TmDDtSu4APSqkuDiCVzxOZAIDsZMpbUAR6enT9mNOLhbtfm5RQcbyXsImpIPJQoQqmvwqNza2LQxSlTnpqRylQItKUtRb/+vEhUJjXiKrMi3q19KVMTBKibfFZsEcQqqkhc685s14oqoWNsePMXXUwHHLyIqCg58KChJjaoZIxKocrlg7S4Bmu8FQyhrWUtR3QVQkizpIijJg4YcnOwpN+URHs3KQPhSI2JUdDwzgdm+X2ivTAED14cfLM83wDcPFlGcuYqDeREKcj47AlUBMqmpcQSZOWAaZNLgWoi1EgFbgFL8O8CmfJxjXw3AKtZYJCIBfEfgF/cYYJiSilCtpUZ5eUVTqHoC4O+NaQrUAmjmHgMcD9ImgOEoDece4vVxnSIwRPQ6iBDPNPo8xLOI7+djHJ/H76h0OjXmjvkYRI0arCWfc1foR+8df4ZUUOD5XR3yBt5UyQAUcY3hew1ApPLgsXGRZlHxQ9B+2qi7DZBKnf1nQaJEshHPNZKdAOp9/vTv25+XAwaMqSozkhoowG4AYQA0kmIANRIs3g+vXc3ZqpNtMTe4lpxEohTeEyZXxMVc4zn0lYn9KqIANZ/aU5IaPSc3AtD1NeLxBq/lHqIxehAPg2RakE9h5xTzSclTShBjTADK+b76LGUgE39nPAOUyOdOustUFt+35Mp/1+erV1SEH3KsE64PsCVIsJjLJMPRVNyFE35GhQo9elg8vX+4spEkRNKMZ6jzef+TekNNUYkHWm1ir7JU3+zR3RKiDAKEkl268qJduXrdRkaxROAaXAmreCsqKtrt1CS+LCFErKdBizJ6BEQzbZ4F5yfXx1jvoxo388qMZG/GdXoz7QMHJZL9A9+Ptaqzd4CoiDn3i4gK1HNn7abtbm3Zo7v3rH5Cw+REVPRDzGefP/lkTbFqfEvX8wuIivylAawH4X3Waany0RmlfyKigkqjgeqOfN+PsczPiphPYb9FHDc9NSsAtlTEiqOt+CXOitifgqiI99S5gAJadhEe56DmdrvMJOxI16ZrSkRFISMq6menUm97bxy3bmHTSllCj8CM+D4ArrgGxZ7E0E8RFd6jAqDSKzVK9s6NdxVDM8+Pa6dWrQyLzDs+qVmpUJb4Y+3iqoRAVADcuvW5Ea4AqADIAGggTHr55Rs2QsyLZd4pdp51AVdUA/z0pz+zpeU1gSsPHjxUpd38/IyaTtdPTqUgX12ZtzffeNlOTw5sqAxg5kpkwPbJpWXberRuDx48sR/+w0cC41ZWV2XvxJq5cGFN9wrQ8+DhQ1teXpYP/DTgf6Eo4FLWIgh+AIYUHxZlXwU5MzE2bkvLi3ZwuGf7ezs2NuyAIGIiAERA1tN6U30RIHDItSoVCPW61LHUuNAgdWRo1BW+iDGs0KuOp6K1dnJoHA2olSdHR61Vd49+ABzO2YW5WbvEfaQ+eVRPYEWEI+3y2kUrVkaspXyuq3zIgdS29g8EVA6Keo5yftaSZdO9u/eSjeGZGh9PTmK7wTnYlGpWDZ6JOVCFy0MdW48hF2yNjElM8OjRE2PP6HKX0ty5kMAba3vvPd6PCpLFxUXF4OzX7F/M9ZmZaZ0rUpZb29oFnkPRpqanBdKOIFxqntr1F9bszTdfs5/+zx/a2sU1+5M/+S/27//tH9iHP7llKyvz9uJbr9p//eP/ZC+/8qItLk2L8JpH8Y24ruv30G4XbHtzz+7cfWBtKyrHQ3W/dvGCbJ/WnzwWeXRGL4vHG7a1e2TNZsdmFxcFINP8vTo6LIswnfOI6LCe5J7pk3B8rMqjrf09m5iaVNxCDMBruVdsiyReSw21sS0aGaaatN+ImTMM8B0BImAm4Pz83JyWN8+IcxgLo+b5meYdJNmHH9+y5jlnzahNT0+pdwN7DrZPTjYc2qia/XbsyZMnIsKxpCIH5cIAldmPonqX/QkyT82Iu5w9bqPDnOB5QWhpTnVRgo8oh+DsJk9jTCD12IcAI6PHlYQr6sWY+qJxVnUAZUd0RlLhtLa2JtsiiCH2AiybmEPsF6jKObeogKIB77bImbItLS4q7rp85QXb3tpSvw6U6Ni6PX70WHsEhIRiFKOHTkvPnDW4sDgvkJd9in2btazYMJEOfBPsQz0k9LyL2ke8abPnS+xtnM2sNcVlCBcr3l9EsUsSyDiR4xXkPBuqciM3kXAzOQGwDsh1In9hDXAuRL8Tt9H2fZ4xjSpZVUZUKrYwP2ejI1T4+HmJw8EZVt4hfDg8FLA+PjlhlSEnI+hnwX+8F1ZiXNe169dUvcNz39zcdJwlxcc8N4gQ4mHZXReLdvWFKw5K1+v2+edfaD2PjjHnTL06yDGvX7+mXP/Djz6WwAebOeJn4iePUTvqWcJY06A+YrQ852RcpMCH3BsZ6an6Fe9WhxI55LhUEEB9UVJUByXRbOozEbiYx07JhSRVQUQcrp9lzgd+4ILVpcover6kpvXqF6L+Io2n+st6o3Wv1IBA096aMKMg+sbHRrUH3bxxVf2CqEqjRw2iS0RSsxDcpw1VVBwd10Si7+xsqxpYPSRVNeMETF9o5qQ1xGDPRWWgmiTGOh/zmJ86r5LVr8fgrsJ0XLHQi1d5/mAq4FE0Wge7YexFGiYsh3XD3/1aK7a0uKR9ZHtnWwQjexbPdW9/v7cvciOyKoYNT6IrtdTKxIVPxZnpH3nOnhMX/e97Batyp5bLVkQAT8+oCrFG1ep56qP7nKgYiO6f//M3fgTGT7z0KzRoLGbA51gggOpSakaSnRJn3/rc4ilKK7UxZNLWSKbahMmUcaVkx8sH0ztoEwrm1/2r5S8vWbsrlv1XHbrUZpz8g1UeB1vunXESORGtvr0JN5sNQZE3BfPKCYJpbXKdTipzLdrG5obKiyOo88PcFQcq5ZO03ZXpEtnAmoqwcVAWxRqsOpsFh7ArBxwgIyn0ngThdepsP3YLSSLpSu4yDcU7NkaT6/OmjQ9VbHZyVP9Zl2fSlS91s9O1u/cf2PFx3cYmJ6w0PGLblHSXsJmgMgI7HC9j5nqlGiLRa/VVrQEScR38TNYO8tjz6xWxo3LPpgLoAJbY4GXVlQAib4zl1lJnDcrh+CyCkoaCef4tT9MiQCOq16ebaQfQE8qDL4NHv3pFxa9KVIA68yxQY+AnSl9IAaKQT42GAp6+WgGrrGEdYJXqiFQYbqdB2Wnfi50DjUA9mhSLlEgqBIDsuVkqKvpERYBBBGLVVHa8vbklhcL03KRUqwRbXrFkOlQhKk4AfLJdJ9aY1utXVFTE8glg8ksgxy+rqHiKqEhAHQpQ1n+6GPyLUYx45cE/FVHRlTUaB/To0IgCTgivbsHJRxTrsqQAQE/gIWsk9olQ7wT4yTPNA4IYD/eE80ZzJAiuAvfnp/Lb1Gw5wGVVcSX1tSs2UsPZ1PMgAnL+zMF1XhNVCdpTk8J28Jri+TyLpODe8qAnXhsESJB4MQb8GSBUgPBPkQBJ4cTrA0T0uaSaXwViQc7kARbXFp8Ve0MQEAGS5cRjXEMQJPlcjOqGfkWAW9AFyC3/T1mc9C1V4llobg80Og+yJQ9kpR5PYGj8flSKuG+rrzMHiL2yLMYaIhZwv1x2ZTf7KIo/3i8nKghoAW5Hh0ecQFAz5OZTRAWvD89ari/mRzzH2DeiSkDJYEbQxLVxD/ydpCHIJN7bk0bAlVM1bwXQiYbk2EQI8K84yZjPx5xEiqZ/IUaIUuz47D4h0i83jrXmo+aKWF4Xc4PvAsqrSV6vcs+FCYxVWGZFspUTFTGv+B7EbthWBVkRpF6QO1wfgIRIxvTMIxHMxy/OmvjMWCuuJfN5lc8hxQ9RMZoaN+bPLUjJuB5+nzNYIgpVu7gKXZ8rKyUnLh0X76vf+DvX6UBhEnmkPTiUvYo5Ol07OqUZcF2VlKUi9jQ8/5J6WfGcRyfG7dqNmzYzt2CVIZRhnMiAVk6uBlHBHFN1IYljIiq4/3yd8ZmNWu0pooL5x/s8i6gI6ycRFUf46zvpme9RrlyNisxOj9iNsR8kKoKg1B4D+NFp2eH+vq0/eCC7mX8MUZE/919EVOR2RczpvKICCFMKZSkSOL/6h/WvU1EhsiT2oAGiIt//Y68d3AO1/6c9XTF9u21TUzM2NQWo6p7hQVTEPhDkXsQ+OfkrIiZV2v6qRIX80wv0EDhVJQb7J9Y7Ue3iaydssACm+7YTsT9p/RK/VvpEBcemmt4GUZHsTP6Pt39P1UPzC0tWrlChVZCwR5XFrY7tbG3KFgniAeABO8+NjR379JPPJEJh3VFK37S6AAAgAElEQVTRTI+K+3fv2urSqr53UjtSPykqIlCG0kwb0mFn1yuLEE5ICKoigY6trSzYN7/5unXOT61Co2aa4Y6PS4E9PIxPfceebO7YR5/ctmKpaqPjEwJUsZ5aWl6xza0tCaIgjAFXafiKV7v2VGz+KkXb2dmxS5cuhLml3b/3yObmFjQugG1UO4yNOIk9Nz/r1pXWtZ3dXatURmxrc8ebggvUwmKnLuBtYnRY85dKa65BFiwSgRUVf/EMW7KGa1mjfmojEEWKSVpWP6sb4BUirJnJSVtbWZWKtsRY7ezap198YaOTU1Y764hAZbR4ttjtIKhyxbgTYy54QzDlTcUPDx30xconRHAAy16NR58LB13dypYKHFfR0mgbwNZ90M+sIRC4pDyJz9FZpnnoqmvPb1oCnY8OD3UNstWgcrYMqIbgqmWlKk3cy277SE521rDx0WGrdNt27coF+1f/5g+strNlpaGK/ec/+c/2vd/+Hfvsw89k2fO1r71sf/PXf22vvnrTjo737c7t+/bOu28JLFtcXrbqmFdt7m3s20effGbdQsm29w5UFU5vlXfefcc+/vn79uTJuhqIFxBODY9ZZWjMCuWqNVXxVFK/R6qH1CScWAFb4vqpGt5iCdbxUgivIm21dLZKtS1bngm354zqhHRWUF3BuQSxAdjvSnjU4G5hhB2axrRnP1lTjEK/FfIqKlxcHa8dSuNNNfbu7o7WKZUxWJ7xvtPTM3ZwsO8Kc6oXRYAgBiAe9IbXik2jl0TK4/SsVAmCLVqK5QQRONDnjZA9j4sYgjyYe5AFDlkAYjYAb11oxxbm57U+AbfXNzZtZXlRa1Aikg59abBdc/ujhYVFWTdBQmBhtbuzq/djrzg4OJGwD5A+YgLyut3dXWs1IWzmbWf/QGM6OTGlatxao26XLlzUukayrh5lNEYulUXE6qxMVYdMZYjBiFPcktl7dbJ2tF9BwJxDwmBlVBXwj5Jczes7bVVYOMDe0rnOmeuWkkXv01nwOBhMRdbSRXo1OEmRHDE9B2N9q1k9eI7nE8x/X+NUeq1ZhwpEfgfySVZvHn8fHBxprU6Mj9rUzIzEpO6YQQzbllWZ7un83HsEpMo+F4C6nVUJ5Xk59YxIz5znPDUxLuJV1c7YZxJvnXdkJS5hiLW9D0hlyG5/cUf7NZdMNZbbNLpAk/iG802VGqqycDFn4EYhwOJ6eeZ8nvKgVPVDRRHvF1ZPUdHtYwC53e+NKDs8ql3pD5oIkIijAsuJXEi5af4gkrMI34fwg5SjmoF9LAh6xiAEday9wPRC6OC4WxIu0/9BGKHZhZVF9ampFIu2u71la2sXvIJW1bVlm5tbtEKlor2Kta0qxLo3aRfpo0pS4pNUWZ6EJv2ig2dXweYYRsRKitWFEfp0Yw2oOXoSjTDPOEMCF6NiQ7UbvXvH4g0SiryK6qcTbz6f+gVi/YW1NGuGr2g+z/OFuOA58ozyPNjdVPp203mun8d4v/z7Pg48a+6JORRuLzzPqK6XAOo5UdEPup//7X+PEZiqu1WL25h40hAJv5rfAUgl3zdtiKXkU6++DCm5Vq1W6uGQ8qtINAXmC9mnutUTY95f/oKpZEkAgIBG9xnUhpMSPV2T3t9tofzAK/XK1mVtJHW6N/di4xP4nbz1YOuxv6CGWbYLOjg9QCGw9WZpJVd0JhVPqDcJZsJPmNeH4iAOIIJoERdSXHiiRbJPQKDyL9SXlNAqEKSJuBMHStgrVf1MrX8SGcLRLtKIAwEFWrdjKwsztro4rXJENnN8Rw+OT+3+ww195nm3a5Ozs3ZYq1kTL/Uq3pXuU0lAqkCzV8rqCrgAXxyo8MNXz6+AD3hVChEGgwBf5ZiUmQLioTpTqS12Ya4uJ7DzR874Mx4etFPSrO8VnR0HYMYWCJB5YsF7VATglQOIAdQ9dfh8lfVTNFpMynsBHi7FEmngagqvqCAIYT4LyIMwKpVsfnFBzwvPDCkJmzRic5IikneaomHrxbg6IO3NmjSGhYyoOD+XuuCriIqZ6blkuyHETpYV3CvlugRXJCk7W9s2PjFm0zMTKmHnGcoLs0wpbV3vT7O8QaJCQaHWydMVDPkOlYMS+SHv99ErDPInOaDejPfp96uIyoqCVZLaAWsHKZjtq4mK3vskYvFZJZEeoBDIOmjBHJYCPVmyOBGWPPZTfwit5QSCSmeZyMN8DsWeFgFB/EzzAQVS2YMcT4y9tNersrpW1Xzp+9Lz3EKFrkCrlwA50Bb2JTGX475FrqRqHAdb+/MnriueTQ6QPut59PbXtGdrDJL1j6tu+h7oAUIznwQKZH+qua+aDYaNUF9lGyDlYFDIPuG9iLynQNgjxd4Svx8gfACe/cDdvfx9GkTy6KXFMQ7s6XFW5O8T7x0EZw4yx2vz94mx016XQOv4M9Z4VIwEiZKTpYyr1Ht4cpd9DrAPYp9BECo1qM4gtwtAYTiSmtaRfLGXnCUPZ6nYKY1PFQwOxEQlj+8r0YiPsZStVOoX4UGqJwphk0IZMg3duN6oinP7BPfNlQJNVUhUBNJk1S2SALp05qa+JbGX8z2dp4lA71kspv2Fa+IrCJF8fXlPqX6j+gA78zkRn8n15uRCj6hIgBDvG+s1kqcgrZRsDQ2lqi4/Q6IahNdFFUUo+uNZsy4D1M3nU34tAu00L/tl1DFvBpOKmGsxD+OaSfx6u2kCUqQqTBYWvQRMIVESVWTWg+qLo3CqI1sPeWzryOivk94eXSzbWRurl0M7ayLYqCSioqjGzJXhol26ckUKTgCscmWI3VMJ51CqAguiIqyfqtivJFvCWLd5EgVRAUDDvGLcg6jgOaGI5r1VUSGA2G1+mHtHnFsoQbOqNH7m/Sr6RAXPJiqd+FxU8MUuJKrbeD1t/WSYrdjR/r7tbmza1vq698hKupacJIgz8qui9i8lir+goiInKkSSpyb2aqJY8F5NeG7/OhUVaoSdKgHzvc0jK50UvXOZmC1oDH43J8Zi79L9Gj7a3tyR8wyl+NT0jIAlzdMUu3Lv/XjOreZykiLGjv0tKiroTxC5QgAlvWNdMS6xp5/LEBVnZ3iWAyDSF6FPAubnns60rMdL7O3yeKY6GIXjad0Kwrm6muNqwpysn9669KYtLCwJPJpfWBaJvL65pb4QROJYBsnG9uw0VUh37bR2Zlvbu7LDUWPNUsFu3rxuG+vrNlwdkRr88HBPfcMQJRwfkS9gA+iNcWdmp1Q5vLH5xA72D6QQvnJp1V64smpDpa6NVIt2fOSWNNMzc3be7lq90bJ7D57Yzz/4XM3tUURSNSGV+cys8gVA4Hv3H9ilS5ekLL/y4gu2sb4p5W+zWRc498ILl/S7VHVubuzY0NCoFOUif4fLDpCyD0jgwUrpWouqsnOEL2c2Muze6Lym0ThRc+zpyUljD2icQaoArmExiH/7sY0ke6u1C6sSzuzv7RnwMVXUstLptnRG4kVFVdHi7LwtLSypR0e92baPb92y8vCIExVUfVlHPuVt1n+KYxxT4n/CYJK9GNsWJ2/DmgTbHJH0EvHUPbbHrhdRCRZsOue86tktboo2PDImBTpNwvl9iHtZaKgSw8FBAFDyAMRJ2JlE7sS5C5lOfoRqnhh0ctobIkf97zBzq3ZkN19cs9dee9luffqJvfrG65ongL8//vsf2vjomN184zX7y//7/7W3vvmmqjB+9A/v2bffec3+7u/+3t79zrdVVT0MobNXsw8+uqVeK1TB0XAWG9vv/tZ37eHdO1Ly0oOjMjyqqouh0XE7OsFCzK2EvOrY83l6HO7T62R22qicF0jHfpWsjBkPibXU6NeFaeohmQRBNC0mWyUH4joczMfemGbTWPlU7ejwSGSWqgvPznq2KYwXFSqP1ze1Jtmv2H8AfkWAUu1Rqeh3njx53LMM4syAqOOMpzrUz2AXJZIP8Pk6s1MfQamkee4pxoZY2NzcSv0AICfo34JimkpLFzEQQ/Hlr230GgvH2efnf1sgOj0j1LDZTI2ZHzy4nxpQd21ubkpWVjzr1ZVlqeXBGmi+DrERCnXmbaPZttXlBTs4RL1fVjUGlnElqnLGxu3B/QcC6hcX6bWyrfMYO6OjEyfmqFxXnt+rUnCvfwkLUaeHm0Ui/JgLYX3k4gEnPPld7huCSkRFEnZgU6WqHgksHZCP6ojTWl0kUACyrBsXxyD+8yOFseN7rKsA5yNf4QmyliBBr754xQpY9aZm4KcnNe8zRi+JjW1VaUV1kDdexraK2NEbPoOpsPdH/KuK2hSfs96IOxDsQHKzDqi8eXjvvr344gsi7ThHP/vijsjrlhwoKmrOXSl37eq1q6pW+uzWF/oZKSVAtc6n1BycGEdNqVMVdlTTxhnM2EaFRPw9KlQR1uHIwbhEPKteUwkLy2NxVZYlcY/6OmXWnL1YsPfMXVzjGJivFz9jPWLgHtkfgpSCnIu+IwHwu42VY0Wy0CIeR7ga6w38jAfdadnlixe0drEM5ZyUsK+L/VNTexN77hDNwhtN7fNYTRHXekVAxc7T34XNdRG2hk116vuaXN4H47d+zNG3RtV9Rj+1ZM0uRxOIFXr2NSBT50Q6QqSwV/EaRJaczxJHyQaqnuy4vPk85Kj2/ZpXLTIezFHEUFwHeZbGK83r6GXJs2UORrPuWAMRg/4qREX8bsSGvEZNxuVu4BbPXqHk1YF63s+Jiq8K859//zd1BCZO3R6h72eX6Mi0kfQ3Mff4ZzNlw0kFBlooHA6e2HjIJvAr23C9pNtB1N4GI6W/b4ShLJSVU2qqI7CNeDZKxBNVKmAngZJsGGL0Kf3WfkXpufviBvAO24iaZH9/T0kI/qkcMJSDE0zheRiJHt6Q+DGSaKopnBpneaNCbwruark4dMJaiuCOJIaNAv9DSj4JKGi2xsaNmorPIkBS2RzJeGquRVUF70cjPS9DBkSgJNvs/PRE6pyisZH6fdfOzu2jW/dVq9BtF6xECSOly2yaChDKKrnmngF5NeaMv6omvHKA+w0yRuq8UI4mAEmEBCCDgnxKO1MvjvRzNnY2Sw4a9QToNVVko/QKCgBlyAqSEVcS+ve73ZaNzdNwqd9wNtTTOUmRA4yan+k/V/bFfMuA3rCr4mBtte0UoqLbVWN0JSyAYLKlwtfUbWggKqSgatR7BEWMj/vIV6Uo8wa0rkCNWgGPBp2N53MI+iA5ohllfpDyHtgu6B5Imak4Sf6TgDoMD8SKKiomvEcFzQs1182kbkKhs7+7Z6fHR88kKny99a1avrQfpUM8vv8UGJLIimftYTHuAoh7jbWdqGDdR5cOJyogrVyloK9nVHgE0Jz3UmX+6fBPDcwpIQ3fW0pkGTWUvgLrGHNmP8EYQIzUKf2KCjVTTeodHeIZyRVAa+xD/BnkIQ3hmetS1kjt7BZovDcJqIMwiaDKlcayUvHblUIn2b/E/I3PDOUWiYkH9ipw9X0yJcv5+A8SFXlQkwNTAVTF+w7+XgStoVAPADjAWj6T68mbO/OeEVBrf0i/oymfjYEntg5exzjnwFn+GUEGuI1CCqR7JG3ewM0/w6/XyYD4jHhdXENcT/yZK7XzoDDfP2Kvidfk1RcBhgdIx78ZV5EAVVdUqoT+DNLV/VtFVoSaq1RSNRwVFZpXyWqqqZ4YTlAEOSClT6o4cMVgEN6+n3DP7CmUXXu1AgqoPtHMa9kzqJiI5xUEAsuEPXp/H3UjitPRHlHhgbMD8dybLKqw5aq6wpSvIEcCKMzB+CB3fA4/Xd0T4zy4j8d45mBwPr97ZFBKbuNzY87mVS48v/59OkjbI36ypnlxf/Gco5Iikuf8M3JyItZgzLFYa/m6it/JE/J4ZpGYal0reff/VGmpKqpUGdpLMZIAY2DzZUx4L+/744BOvKQ3ziStxaLK62kWS2MKj8CKZuWujY6P2ZtvvekNfM/bUrMTQ6Bervasn9oiAxxMGxVIGURFELL5c+NcxRIliArmHz9nrtLEldfwMwCHmCPMJ0AnwJJYb/ma1j6dkYg8q3heKHSJZ1w57X1pEB+oHxHrp2B2dHBo9cNDe3z/gUBc7UfPsH7Kn+3AcOuf/XT+q8n6Z70uSGLiCvnD43MuYKHwVEWFEPaBPTTezxul98+CmJOaf2AC2TkWe3LMyRzs7xEV4V2diCF+l4oKrOAQNMjSJZ0/fG6sIflmJ7Ar1m1+XRLhAKol66eY93FfOqITUeEWjEWB/c0mRAUCIxe9hCpezyoNQh6TxDmi++H/iFHOW9aonabKBW8+jhgIsIrff2nuZrJxatni0rItLq/aj3/yE+3VNInnoD442rMh9Qfya0NA8tLLr8pehisZGub3sHE7s/ExGsXTqPZY9wAQOTpKTxZvrDqC8rjTsg8+eF/gMsQAYP1bb7xiv/0737Hj3XU7Oz222dlp29vbV/PykbFJG5uYtp9/8Indv0/D0XEbGRu1x4+faD8mVyBGjTgT1STVtVT/YiGDDQvfg2xZXFqUkIheC/fuPlQPGtbH9vamLSzMClAHGOXZHteObWFpXtdx6fJVq9cgYIiRvQE95DXk09zUtBV0NpSsVj9WHkKvAGYLoOTk6ISqhSj0QhlLI23AQK5pfGLUTk4OrYrlTKlsp1jfzM7L3x2C4vb9+1ZrNK08NK6GyuRNNA6XkUVYzvJJ0ro4mKrYWupdV7ezJ7K/AHZBLLi1DVXf3pug2QCo9XWG+EIAHzEcBIlsvCAniHeGlWuG8tZJdleUM140RPZ98dyr81KVGeckoBdzBUU5fReGR8dVcTIyVLFS59xeffm6rSzP2Z/+yZ/Zyuqi/bPvvmNLywtqVt4+8zP9v//Xv7VvvPWWLcxO21/95V/bD37wbfvzP/8z+8G//L7dufOFCEUqXz76+HPbPzy2UtnBZOyDfvB7/9LufvGZqnsmp2do6mAtYo2OKfcMO0gqTqgQV9xRKNri/IKtb6zrTMEqR2u91VKfBZT/skgSeF/vCQchJQB9IUjI1SH+ZDE2PmE3b960z27dsp3tLZ0BL7xwRX0cfvzjn2h/mJmdsSsvvmi3b9+21Qtrtr6+6cRUu23DI24txpwCKN/a3tK1cm54rNOV+tnFkEWj2TYWRTgXYPPEe6iCARcA9V7xcxIQO8R23CM2LQhHBCZL/e8iNRfbVVVRDzAPOAl4GQ1z8zM+xAXYsKHo5wt7J8YJ0p5xe+mlG+rLQG8JjVWxYHt7u6qu4OeMD+saSy3A8NGRUTVBZye8du2KPbr/wFYvLNpLN18W+XXrs89ll3NwiDK9KEEK9jyugqdvxLi1EFWlahKeCXEq1Rnsdx6/gM3Q94XPRzCJzQ95vVuB+brxiiS3sXbxKdcWFZ2MqaogU38CwFo1HU6WPb3YRH0UEIqGKMNzdMac/Je40+ehE1zs/5Pj4zY1Mex9LcoVm5makmXW7t6+iCE1foYUmp0VkauYDZKxiJUTcWzZ6k16EJXFkLDXyW7s+FjXxzo9PTtVjLy9vWcXLnjvinl6XtCvo1yx/WQvdXJyam2srpp1auplEUiPIyqBDg+O3cVDmi5u0PET5iPXJ/FXT4DbFws6ToSFkQvbGG/WJgSQC4q8oppnwxixn/HleIvvj3H2sr9y/7wnJHUejw5iJcqTUmNsf71fE99nbUDWBVEHAagzWPid586e97io059vVJs3tS6FmbAPD1dsbXVF/X2Q0Swszml+0YOCau7F5RXb2z8Qecp+S9zJfXDWeV8rSG56QyX3Ag4VKtg0d108LavSXoTwdPSV54ExBoNxultgeVTMGIP/0bz90aNHclNx0tKxLK8ecrwnxIbMQ+Z84HsSZGF1mmIkfu6Vpr4uPV8I8bGfV94/os+4RO6T300eYz8r12BgIt9AHOnVbsmCX3tkPzd/TlQ8K0p//r3f6BGYbqDQ9IoHLZDM3gjvSQLhUChH93r5MwMYR4OXUAYmxE4gUfKKS8XdSbXS8tel3geeGPrh6JuTN8ON3hO8T89KSqs/mv/Rp8IbSam5ZWrCLcCmUpXCiA1KDGOno42dQJGDBUYXFrmoA9qb6fB7Ony1QdHwyIFs3k9KoVQixmdF6SOvwbNTB1DyQ9ThNeINrQT0p8Oc4IhyXPeXdfCZEjwlh8kvEI9bNmeSDoJpfERHK0VbW12wi2vz1u3QNK1p51ayj27ds3aX4I1qh2ERFUM0BkqKCLKAAqrvZGfCAaTDJan8ODRQUoUS1VW6Pg10z6rM8PtiBwxAUvekBNjBTbZ/Aje380glnMUElZQ8kKcqlGd6fu5BFgnP6NzEVxIVOagYh3T+vRwIje/rEP41iAqpr8plo5m2Kl7qeCh7IBDAZBAVBXy/U5MkB7cizSYC6DdolsXLKUo9VDl9/3V+mzk5FUQF5Y7VPhgEkRIVFbvbOyIqJqbGRFR4LRHNzkbVCG9zY8PqJ8f/JERFfsin6PKZ+5gvaQ98Xa4QtjE5UeEKbvcv7RMVeYVHDqrooB6o6MyDrUqZgMwb20elFomvl1Z72bcA36TY1DyRrsurd3LgMZ8jg3/nOqLaoN50Kx+er4+NW104CeJlzRFg6HsJqJV9ARVMqaFvAHD5HFC5b4+g6AcUAVw9i6gYBKOe9XDiOhz8BkT/slI1wJ8AfQXGpz0tH/PoEcDn9CszHC4ZBI3kf5sqFHKyorc2VWXRt/1hrFTiD9GLtQAq2KTOiSA51p7OjqwRWVx3BNpRhRX/VoCWbAF8v3ZiI+Z3D9SNvTH1R1DimPpmxLOUijA1ro4ELJ4bREVUAZ43AVIJQknsuw62pFJjkm6SX5Vzt1MVnghknpGTVPn9x/3GcwqgMa6Fs4D9OwimqADg/kmUmb+QnbKv6vVDcJXQ7u6ezkIANREerY72KPeR93UstVwiLHjPIEii2XMQrjqLo0l9pnoeTJICuMyBaCeAWLNfLuOO+5eyT2q/sEPy+RP/xTyL68mJv1gH3EeQS7xPVMYNzosAwQdB1lhjMXf0Z1Km+X168h9fca1BegQJFmtfayk9E4EoPXs639f7FRU5RN6vaOJ3AKc4U2K+B3HCvzucR7JIKdre/ok1Gy3Z4WD9VCgXbHl12b7xzbcFDjWaLStXhwUykTBy5mjOAd7uH7iNWCIqGueu9OO/iBHinqmowKZibHxM4ALVqryPiIqsoiIs43idiIrjIx0zz6rGGSQqYu7z+YcHh1Jt87ovV1QUrF2gouJAVibrDx/a4cGeLvV/hah4ao/9FXtUxP6otQ1RAVj6jyAqcoJMgEMSRzhc74ROJLVPxT/ZxPTv+7mtsyHFsjMzc7I04Aznd6gEi3k1SFQ8Kw5jPrpSuClQO+Z9nFV+vcke1RAMORhz3qIHBEpczlOICr8X3Ws26FprGZETZ0wQFSCxZ+xfqpjMiArlAEV7feVVO2t642ZAp0oVyz6sRshHunZhZdnu3b8rSweNjVSRkzYyPG4Li0uqjKid8rO2TULuCfSmyoNKbEBxFL1dOzg4li3LGA01T0/s/v17so4EXB4fHbJG/cimxofs+osXrVTs2t7Otg2PjtrE9JwdHZ5at1C29c0du337gaorIBzu339gS0tL8mkngsLDnobD/GyT3mUT41J/q79dqWiHR3u2urpqpRJ2IG17+OCJzc8vqkJ4Y+OJzcxM2cbmunpefOc737G/+/u/tYePHwm8f/fd35Ilx3/8j38kEB6RSbvdlH3NOA20IdYrJVVlWKFtJydYX7Wtc96yCysXrF5rWLVUVXNyPr80VJZlFvaIp7VjK5OPAaSkUBAAfW5xyfZoPFwDxGpYWwKPrgREDkh9uQ9LgFlu3dSwoWFAbBcI6Hwues8oNTJNe7PEK8m6hPxD1cIds8npqZ4PP/kN+YLHIGYjWM6kJtGuBPeeLBCgbpnrTYbp00BMSl+CspoQj2IYpVgRmy7rnFuh1bR3v/2WvXjlov3lX/yZ7Gvox/GH//r7NjE1ZBM0EG6bPbjzwMZGJ9Tc+q/+/P+z3/u979kf/dF/st//g9+1zz+/b2PjwyIC3vvgY9vY2rOtnT01ZWaJ/Jt//Yd2dHxot27dskKlaoeQd+Wq1jbCQvZzwHnOfOYUfz58+NhmpmdlFQzw+9kXt1UxMj01YdevXZWo4c6d29rT6cfy8ksv26effiobMippbty4oTH6+NNbGpP5hQV74/U37Mc//pEdHuwLzLx29aqAv431DRE+gKLXbtywhw8f2tz8ot178CDZqrbtpFbXHsC5A7g5ir1miQq8jnh2cAevDHXVv+aIbCIRnvWdDsANEAQSW/BcqA4KgFjxAOdu8toXQCxS0/cuF4I0PCYquDjHVcnuIhFVvbIPandU8XFygv/+qV2+tOYVFK2mLczN2R/+/u9rV1MFAfvKzLR9+LP37If/44ciQZmnAKQA7owVcwdLN64D4o1zi4jga6+9qvObcTk4PLa6qtSpSmT/9GoKxljEUsvV1bpmNajGvo4xTcrq1Jg5KuTOUnWUW53Rm6ehsWdM5KKQznziScgNBIt8RYzI+NFvjZxVxEesw5QLeR7iuVFYZzNuqNol/iImk2inlCpU5qzYObfj40P10akUy1pj4DKIcFzAQ2yzbysXVm19fSORo/O2u7crwSk9PMjlA8eBZOG5sl6nJ6cYSs3X09MT5T24LUxNTtjly5dEbKCGpzID5b9IyxLNkU/UP6VYqtitTz+Tzevo2ISwEMX+skCCbBt2Yk/iK8eKooIh8hmeT1SSMteYn06W+pyKM8+rRdziNvI47Y88fazHVY3vAgPvI+WkAe8dzZt7+Wmq3vVcwj8jnEE8/oocvphAeLf7Vn/XVCEfdvAeKxN/uRiAa2JtkO9j+3xpbVXWhqPYOh0dqHfL9vaOCLuxiSkb55ycnBQ5wf7BM6PHGc8WuyTOVBFpEtS6G4PShHB5oM9DwhUj7okc6VlEBZhA5Jac55LIytbcbd7HRkY138Tu7a8AACAASURBVHGnIC9i/erskqWvP6u5+XmdKdwr5GnYmwXZVEqVwhBpIjgPj7wHbXKecdzALcAkwBHx2hepPBVnpn/kRMWzfv6UyUXq1+vrzQVv/SqO59ZPzxq/59/7DR+B2TPKab0hJZsZqnep8v9/9t77Se7ryvK8mZWZleV9wVuCIkHQgRaUKEO1pJHazWy76Z9m/rjdn7Y7Nna3Z9qJlCi2mnIUHWhABw+U9y4rTdXG59x3M18lAbLdxoZiWQwGgKqszO/3fd+7775zzj032R8EoOFAiv9cnp3pUBFKBrdq6hw7/MjhVr1RTaHDegqSbSY+sfhxQHFldfrlkFola6rQInqZvHvwwoCGDYkAZQFoXn4vBrtS0YZ08uQJBWgC7NDwiDYXtzFyZQ7XGKy/PPqSGpakg0MitkWMSxAN/nNPErhMNnwCrZdL443alOqBTYXSMVRfNBnyZKvX6lhxNFs2PDwoMGN93b098fkkiJLojw3327EjUzY+OqRG1ahfBobHbG5hyVbXt21xAasFbGtKVkL1lIgGniWHCnmRohKiaqPqSRhABSAaAIgASflIOvDL6wM48gOBJ/re+NPJKb5HUIZh1s9U+kvDdJqFSyOscWC8AI1pQMvfOQxB7PO9vnFvwBkgcYBR7YN3VFCkqpyw/FKvkNRfIgdyNS/aRAUViVRUuHcnjDfl9QcqKlJVRt+gl7juJ09XNUqnbJjxhPACKJdWICxqYgdN6mcRFa5CYFxg3nnebVVjUiowViPD2Hd5NSa+tahWuR+UfowbiqHlpWX5oA6O9BukRTQ85Xpa2BjMzNjOf1BFRQ4IfBFRkYc3EYl74Snta021AbIpqXkfmKQaFYCTVXjEs20DyF2+HD7vUEeXrK+vbBKcCJjBJs0JPQEcyX5O4D8AdRCsye7Jq3dCwZCeUwx8+MNnoGMkF7vNWpr7QVAAKrvqEkouPOQFisp7O6lQ2sp6L9sNQJm/R/VP/BmJZIDkbpN174qK3J6mm8gIsDYIkDzJ8TNIPKMOmORrzBPXOIDFMyEmA7AHMNbeD1L1RFy3ktS0dvheVJAEeO6K8Q5ZECB2XGccmLqJkPx+Iv6QtMuzOv0fnx2K7Hhdfm3ceYybAw6dpsg5cRRVUwHOxeu4jrAa4v2jJNurIQDD/P1RyAGG+Wd5abQOAyK0ijY8PKLDKnFIr5HPtSv/g6zwpD8l55k4IGKHK9ogp3e1BuLaYl5JEZ3GRr0FKv7eHtNRhtVsdW1N1nL4qatKornvTSQp0cd6DMuv1NciiKogKgLojGcTn9seVy3OpPvNqmyc7HPiLie4YswjnsT7BtjJdQBu8/2cOIr30nUhKpCHNgDEnmJlfEYQWPlaCCJBeQj9h1TFCNns+1nb5ioLcrEGcsD4foBwPjZx39p7Rcx4PIi+HP5cvUJUayjZp3UfUA6s5eTxTDVmrJ2cqKCaQhYqsh/Yt6UlAEXPi0rVXnvo/Nfs/IULAjy2UTJXqrIBoyIW9E7jvL8vy44vIiryPQD7HCxf1LOp7ERFgD6rVFTs7+s58n/s7+yNUVHR/ZwCrM4rKtxD29W9iEzKBbe1g/AH9BApxwGN+95v2SbVGq2WLc7N28zd214ZwZw8cLrr3MWXHQp947mfji8fDYfctbaTrds+NiT/DqIi9uU87/aKCt9n4yufk/le3h0P+RnPATUhQDogkL9N4XNERVinuPVWqkzUB3b2k0adOALZ3NlbIs772ulUVLjwCMVpXUIVPbOi2xXENbdT/LQP3uteVKFNktTclwVmMT1XGRyqStYFBQ9NPqRqEXI3rCawKUFxrkrX7W176MEHBS7JUqTRTFYipkoIgFfiKU90YKDPfcf3C5rnVC/wTFFoA7i8/eY7Njk1aecfuWCry8tSbQMcE6enp8ftiUcftr3GllGkVmhxBinZ2vqGVYdGrG9gxLa2du3q1Zv2/oef2p6V7OixY8rt+KxDh7Csot8ZzT3rAucBdrg+1NvMM66NPhsAn1RYSNm9wJockDqcPYicG4W4lJ/p39581Xvu4VE+PjYhSx35updMAB7VEEwQBF1YhABueiU0Fe77eg1Nw2navbm+1faKRywGUcF6oB+JsfftYndbocWXDY+P2d35BZtfWrLeKpUoBcUhwB4AX82DBKCKak1nUhFqVDMkwFT2LiXyQwekUO8CJkVeEucz7jFiDfOZ5ukA+fJWNwepdW2p/5V8yjkHJsCa+6nXvLFvzFdiDyAj5x+qJonhAogYP2x7qhWr17bsqScetcGBqr36k1dEGN28M2//+b983z68csUeevicV3L3lGxwdNy2l5btV7/4pV186kn767/6G/vuS5dsYX7VioWmPfnkRfvNG2/ZXREVK1avo9zet++99KJNTIzap59dtc+u37Sl9U3rHRi2Rx+9oD6Bl995VzGZnouPP/64vf3227a0tKLvPfDgg3IR+M1vf2vjE2MS8j3x2GN26/Ztu3b1uipCAfTOnD1j777zbjrrle3cuXOah9dv3hDYSLXDI488Yr/4xet6fow/r+Hrww8/1D59/MQJWZZ99PHHdvLUafvwgyu2pcbrQzr7IsoTHiAymx4JbncpoqCnR176snLCjx0bKpELDa2POOuqeiTZW8kGLfWH5NxHTrSxDuDtbggeU93CmL8T79STARcFnd+wC3ZXAr7inKuY0NevChGab3M+P3nqhH32yWcibM+ePmV/8l/+UJbHrB3te4Wi3b5z137yyk9te5s15H09IB+pmiIGcV5E7c/PFuepSjE7e/a0ffLpdRsZHdEeivgQHAH7NwBWxxaIKb3KL3VfhR6NCevCXV99jbMXu42Pn0/5HOW8iZDx/pIIO73qwsm/oshOYooTEXvtvVwAeaqAYW1JUJmU/nFmkCCHfkLKjd0Sg8+okX/oOVLFwdot2Injx6zHWjY/O2uHDk1rfh05fER9lMhT2ftPnDhhN2/fUgUP1Q+2V7QjR46JdNV+1aiLWOPZM7+JC8wTWUpKlNXSPge5M4jF3c62SBFwC3Lk9fVNkcMQiiKEdmpax8zvgYEh++2bb6p/Ec/TYylVBr5r4b5B3kSsLNGnEyxB+JWfVaNGk3GVULRJU21EojsO0PPMANZVDZaA7YR9EPf9LOJ9YrC05NmxPqiIoAoqrInjzOdiPT+XyhYtnYM7+21RawJMLPpWMZf5fK4FOzUX//oZ13s1su6coABnCocVFiCE9INnz8i2rL/Xr4097O7MnPYtqrzYQ9nfrl2/JnICwuXmrdvK5ZgbVFREBadXeEZG4GKLuJ97kRLduX7k+Xr+qSehzo0p16aCh3XDOKonB7GEtdTv9tuME/frPVuwkHMCR2Loglc4S+SsOeAVXVwDWKLEvgnvDIss5VFBNmVpY44DHMwmO3lRfP9gPpek3Qkr8TS1IyZsWz5/Zf10r2H96nu/yyNwsge1gvv9qW+CFC7uhQ2DT1BTw6FUEuubz75b5eBFCQifkkp3xXVwkVLYnkLJQf4I2m4h1078dHC/50qNH7gNlQ5lKglOPTFUWh4KameVPUj5ohWjmvoVEDQISJTyKtDv1lQ9QUCGDWVj5XoJKiIxBv3gzefSzIseFl6y7gpWP3RvKnhz30omUOOgriGhT3YeqHw5DAA0ERxJuijdJjHm74CsBEtAWBIllQim8urBgT7bJWlqNezUqeM2MTamhI7NlDK623dmdQ2U0RNAuVcSNqmBU68JQnwwwCTvJJ+QJSg05CsaTcoTeKtkM6lsSVxEUiTVGaPqICebFYCYN+b2e21IXeR2X3sCwbzxYMFq9W0RFA7mUykjfrtNVESgDyUq95F2ps+VNuqzBcKgFvWx06FEdmPi41WGL4V7o64yXP6OAofEjKvzSopyUhe40lDJDVZQva7oVTWOSlgDTArVISfwTAEoXq5j/cTYk3iyWeckSgBpbpHhSgYpQOjb0apbtVrRuKOWWlxcsdGRMSUzc3NzXnLdS1ku4EBLFRVUf9xzzWhsPMHON/VYXrGh5Rtge+mpIsnB1Bzc83VwULERyYF/RtH4RO4XpQ9zwb0ukvpYP73X1bp9U1thneYspKMUPiX36lfj+6TG9z41vtbdx93VzTnfEeCN8xKdpCeJS9vltO17TH6WAkP3IPGcmOArgGXmgRT66h+T+vPo91xRH0pv/2w/3IRiXvMoWWTwnrze+1TEuORJRg7ZOCDe/Sw79+eH8AC9u8EpzbFEKPjnugIRNWiocqNyQKBmOvSjJorDfYxR/t6h4JBiitif2VzxPQfJvVcPn8d7SBWVSJ0Ar+NQk8/FAOYCSA6CIoB7/h3KrnzLiNd3K1byNRBgt/a1VO3ENeS9DuJnURHFz4ntsZ/4YdeVMexDHOL4DJG/ibwiJlFNIdsslMSKx27Zxz7THqMA9tUQ2atP9LzY0xg7QB7mVsubX+dgvYOBqeF7qv5g/+D7ajScSHY8xQG7OBCrsaWagPo+xxyNZxDkSVQQtudK9PtJgx1zKuZkHk9CtJDPz7yCIED8WFfx7/i9GGOuPyflALKIKdg9yCak4f1neA3jUq243YHH8I7iKxL4fA7HZzLOecWDKyj9K8ivHCSOmJiDsfF6rxrpVFnEc+LnOVHRzqmUv6TeIMnQmWuP6pN8vYcwhL2UucBzC7IixtkbO3pFBRtvrdaw1Q0HZgZGRu2J5y7ZkcNHbX5hUTkcCnPeV/Gsp1NRQdNYPkPWSqWK7Ta9osLL/H2PjC9scCDUOaSjrMTCA2CHa1tXRQWNI/uTTZPb/Lj103pbnJCPacwBSIV4LhpHRCDNhioqSql5Z15VoWfEvZjJooVD9vryst26eUP9IZQdtomKg7E1jx/3+3vkl1/6WlkV+NrWs1Dzzj35wKs6+T4fHeCCKllTWX97HvpsbOeYAuKy++meLzF3/fe7qnNsXwAXBMXI2LgIC5Ee4M5B7ifRSOSL3iTVc1m9ONm7BsDrop1OL5c8FijuIiZJVXdUM/B6gH5XM3esMdyWwe9VGqeMGI81qHWbei5xObvbOz6uEi24P30x9ag4PXLGJsfxkSfG7UklDpAFIM3mPNw/qEqJY8dPWKXaJ5saJ1KaIpeZvzdvXBfYwvzm/gHMBEals8Lq2qptbmwZtjpT01P2wqUXrFytysJmr2j2s3/4O5sYHbDB/rJdOP+A7Wyu2Ob6uhrCQlSsr+9YvYGlyLpdvXHXNrexTBqWUAU1sZ8F3PIN2xG+Nz83b2fPnrXZuVnt1Tx/csKpSaxLewWU3bx50w4fPiILHIRZx44d1dlriwpy+noUIF0G1ZvCwaiy7ERbDQBjqh1bup9qb49Uv5AiFaxN1OetV8AYzxlvd3pC4OsOMCdgkDXOmaIHu6WyQEAsOwtUTWARVavZ2PS0zS0u2gYgXZUeClQheoWll3M7iAzgByBPbh45PjOE3Im8mKoS7oW5GmS+A0odG0rF35ZbOAkEr+3ayNCQrp9x5ctBXLe3FVAneynPMbHeZVwZH86/5ITqU0Azaq0NfNghJwDz3NKv1aTJt1f8fPvbL9r46LD97NVXVI2wMLdif/rnf2SX3/vQjh8/Yrv1bTU1f/bZZ+zQyRO2vbSoap7/46/+2l649LwtL6zZ1saKvfitb9kbb7xjd+eWbHl9W/1RuIfvf/ebNjUxZtduXLd33//IdjiSl/vsmWeesvm5WREF5C4QWVRlvPvuZVXBcXsXLz6lHPutt9/SuoPsf+zRx9UX4dq167rfEydPymLq7bfeSn0dW2oAjm3YlY8/s0qlx44dOyZi5LXX/knzlfF/8cUXVc1x5aOP9D4jo6MiKq58/JEqexbmF7X+NzZZUy7yI25634eCTU9PusK9vtt+zsqb6EOVrAp5dqzt9llFVTEuvmnv68yjHs/fZGMla2LHDqjykA3Y5qZ6w/An5EFYFnFNUrcnDIT5TD+WocFhO3XqlC0uLmiPGxsbtZs3rlqj1rSvnTtlf/LHP7LtzXURVpAD1YFBe/+Dj2x2jl4Lw7a8vOr7aRWwvGbz83M2v8R5j74y/SLyOQdyTr9xc0YCP3KbrW0IyXHNU/Za5j9VHTIh5r4bWI+mnhACvSu2DSYDYQBTCiknqzjvGek5ovvtszYgCrleYoSLsfw84HmmkxGMGWss1qowk9TDgJ+poimJzFxkwt5NDtEB7umxAjHFOdH7ZexKjd9frSiOcE/c2+FDh0QIochnH2IdEmuZp9gz9RRxenDCvre/qnl9SD1BcEQwnfuD3CIuEcPIv/lcng02RRAVEMzEVvonoOyHPMJiDqyGpCL6gNy+dUuVq7pf4qas5sjrTYQO3/NqMhfPaG9WxaLv64o/deIlxENdsZXflyVX6tcCRkH8UU/KZBPq+bnHKTAUMgAsBKX0T/1C1ag5RHjO9GrPUr+S3l7vnZdsQ2WPlbABLK86PVq8Kpt+KtrDVKXhZ11ZcinOOgZCjI6epqyTck/Rnnzsgq2vLNr0xJj2MFXDbNEAftdaKRfANl1V4erXWpcFHOuR6xRmITFs6rslrC+3SXJMIq69nfvmpc0ZYB85f5zJiL+MCvktYyobP3p+QFSDC8lK2vu1MD/Infkd5UZUr+h85wbX3n8O+zEn2L3S3Ul936Mg9N2RQHsMQjLhVFkFaZDxyTkgcr7uP/OzSJ5fdeM48Xt5jv6V9dP9RvWr7//OjsAREq6kECbZiIN8HALEjEe3eQBVNRtyD1WVuqfAxoYWVjWALVIslNwPEdVbe0Fl0KWUqPc6yMk+qHM49ooJ965rsxIhT0zscX7g1yEqVQpwQOJ6OYiwmQEkRcn78sqybWzuSBVBcJmcmNDBhPEgoFF+KMUppceNWkqWemxleUWsevh7k7jQoEdlr3OzKsmcmBzTa9bW15Q0ifUHLEgKVmf03dNOfpXLS9qUx0aHtYmSiIwM9dmxo4f0uwzT3ZlZNf6j1JWS9nrd2XsSHJrARSmgV3u4uqSd2KkXiG8UCubpwBMkR5sQSkoMPJaVsHkbR7HzgPhSHezSTM1L8rAYKafeAeQobLgkRCRaddRYTdQ2AKf8HvY6TauOAay5XY1fnwOAUssnhXx3cNY1JzsxmlGrAR/zh6Q1FfNQ1aGaDnoFcCDZ97LVsogpGuh5EzBUd7IOoUE2frq9ZSV1HGhJIBx8ioM4vonh+ekkXufL1bN85dZP8b3YXHnGEBV88bnyqdxjfHtsaHhA17y+tmnXr9+WFQGzFzUJryMZYgPkf4iKpsb+3l//EUTF5zc+b2wfwO9BogK35oyoEFEURIUKRu9zpWRxru7XmBRYA31e/SIvdhI+j0WsXcURnkryfuzKUdqfIRVReh652rl9TzSWT4RbAPaR+Dh+0rG3aQNPSgSdXo0xkKo+HYxz0JN3UILUrjpw0i6+VBaeCIaYG/GecR3xWt4/B9u7geE2GZLIJV19pq7IFYZRZSAfVVkWOXER4K6/loopj4NKVLNYmyeKASDxHiIzuyyBAqztvvZIvOL9Yx7lvx+kSA7MO2CaPKdT7DxY6tpZj0EKxrMXZJcsAnOwnL+7ytiBVL4ELhKTU0UUay+qDALED/IlSBQ+T8+USrQE6nIgCfIkQHBURPG8olrAZxsiYVe+ySKIlR1EhTyVnajQPaQYGfOGR+2kQ0t7FQcc9eNB9aQmbjvav4gfQSz5PTaTvaEfAHKiQiqkfQfG8/GKZ5lfe76w3ZO+U70S19shVZxUjvUR49gGqRP5khNHPj7Y0zAOTrL5wczXofzJFUv9GcZcjnUQ8yafE3wv7iGuJ8D/mANxzfmfMf9jDudzRnlK8ofNiYr2HMnsnqKHl78+kZjpcJmvsXasTT/j88Kmon0tjCfjnogKAcCFoi2tep+Isw89YucvPqM5PD+/aNs0C04NtAFmRcom6ydIBCr2NOfLFcutn4II8nsGuN20ldVl2ZZwwOZ/iArm6draig5vrAE+l/+5Xq4dsCEARglJsp5TEpWkSpyYd4yfyI/1dWNlRPVTWIQ5UUFO0yMv8Eq5xzbX1u3W9es6cGt1KR7+60mKfG5/2d/ztSHPYE67PC/U2PfLb7M3zeN//lkiOMlUiM3kSQKH/F6CBMtff78DLM2UuS5simjUrD5zqRm1mjwk8EIVK6kZrYiKPYgKV9HzBRwdvuayOciIigNjlMgGWbnKcoKc0Im2iP3xej3DtgUa+E7nemKf6cR//1kQFYlx94oqKiqoCtzus0OHj9jExJTsbqgko1IBcAlxzmBqgE1VMYIVlLuybWVPpgFzjSbVKwK/+EIpubNbt4F+bGlcmUzeKcvJlFt/7cEHRRqg6gfsWV2Zt29+/Tmbnhi2Rm3dhgYqtr66qlx/8uhx6+8bthu379rMzKK99e4Va+2X7MyZMyIaAH8hSBinO3fv2sLCkp0794DduXNHlhoSr9DotgWwhz3JqJ4Z1iisH+YKdlBOrrQEhjYkiGkJrGdcdrZ29LN2/kAsJV/erdmRQ4es2l9RFcDc/IL7cisPKaoanBwNkoKYuyd1cJ8DPogUUBSLlPfeYcQT/qRZqvoNHDlid2dnbX1rW02fsWwJhbjiZooHqtpOAJ4U7VIiu8Ui8QnSw62AfE+E2OF+eQ+dOVNPM64bsZyUzHVseqsCjthLBF4r4WN/SaBnnzdiZh+fHJ8QQct5jXyR8eG5UwlAzlqr71o/TWLLWBW2nJS0PRHnu7Vte+7ZpwTAvvrTV2RpBBH8F3/xZ/baa7+2i089Zhtb6/bKy6/Zi998xo4ePaxrPHzqlF17/7IdO3zEPnjvfdve2rRnnnrGfq2KihVb2dhW9ctec99e+tYlO3p42j7++GN778qnVmdtVgfs+eefU0XZ5cuXla8yFy5ceET/xvuf8Xr8icc1V967/J7mMM21n7p4UdUON67f0DifP3/eDh86bL/+9a90vwiILl580ubn5uz9Kx8qzzj/yCN25vQZ+/GPX9EZl/H9ve99z+bmZu2D9z8U+Xf+/CN29PhRW1xa1LV//NEnEtZxbSiWsU4uljwGSAxYMO0T5DPMc9Yw/0ZAyXxxVbr3LQtveFWGpl6KxBtAd0iNIIBRQIfAReKiZlMElIiwlFNhhUXFFdckq6hkqRK5Y1jNsRYXFua1F43qnL6o53T6+DH7X/74h7a5tmI9yUa7OjRgVz76xI4cQ2g4qZ4s5b4BWQ8xH1792c9sZuauWx31VVUNBUhOs9+wiP7s6jW7fmNGFmxc10Ai2yIf3d3eUmWK2wsBpkLqlCXs4NqJJZwzaQpNNRBxXfmhxDatBLb6uiF+EU/c3ojKeM4A7tXve7KfAZVnUdkiMhVgGosx7xOBWBO8CNFXa4+qu9izEMq4gwBbGNXJCNWmp8atXtuxQ1PTel+qM+k/wrXTL5S1zXvz/CYnJyS8qfYO2NWr14VfgHlsbm2qFxd/8h7qaYjVTvS2K0AoYE/ZYxWqQGrb6lPAF1UqgOvYoTF3dtS3pGwFzkay5MYqtSYyguuGAJLINQHQ6pmSiAqq1hzLclKDKOgVW14BA0FBxQ5xhSoC3iOaIgPuA577Hu4kLHNf81C4BNUabvfE/KaaG6KJl4P9hL2U97lwsSb3xDPX/ksVDoC79npwm05fUvYRzwFMVk7sjfF8iZX8vlxKAmdTLxKs+Oo2PDhgJ48dthbiXyyztrft0UcftzffuWzFUkXiGcarr7/Xbt+6qX6qxHP6Vsg2F7FrwfuVyJZLB/uO8Nhz+Y6AKPKGODPeM+eR84fbl7PeRRqkvYIKHirGmFtRJbK+5ZZg09NTiuMQxpCsXlEa4gmIThe+qBpRfV6jebWfT5Wnhd28OB23AhMhK2v1Tm7j9xV22p/PMCPnyXPDOI/cL8/7iqj4skz9q5//To/A2A4Ke2cbAbFD5cSCIJGMRRi2SAI3el3NwsE4Dv/uZ5jUhbKZTKSCKMZkn5NGKoDWAAsOOtW6Uj3AyDjIRMCKwW6XuyULB20NyXtSqvoE8PB6eUYOeDkjyQ4+i5RTchCDdOCL5JsgiuKIDZJ/Ly4s2cjIkIMsBdSFbAQtbRIkqk7seINxVx5642o+m/eiVA4lFr8PUC0fU1WcOBjERhIqQRLJgf5BKZV22HyrWFat2Zkzp6QmWFhctNn5eTXQYnP0hI8g7806AXtFwCTvVQgDPwg6K8/3UQwA/LrvKgC8j3wARyj4w86D10M2yDORtEKJintPcv8c7vTeKJdIMtlgsAMooiDASxeG3PufULZIk0FICtR13qOiQ1TEwVvEVQDJGSHQBjUAqUh+UBgGUYGqThtKNId0ooLEM4iKCiQOhFwiKmiM7UAl6pKSlSolV+ZJqY8lyr2JithgOgveD0tsEl9EVLCJoW4K8BkFDVc7NjZswyMD2hSXl1btoyuolapKskgQ+T3mog5LraYtzM1Zs4664t5fX0RUfGGQyioq8k3UFWY+Jb6UqNiloqKbqLh/RYWMehPAiIINixopeZxqaqu+UX8xt7VRJ7IgB58C3I7NPScrcrCcz2I9BBCWVyz4dUANpoQjVRZFUkDCHtMxAO1QuucAbDuRT78PgZnbdeTkgCeHHfIjrj/meg5cdmKeq6BFomQNqdtxNAXNICk4dEcVgAOnxB1AX+IZzcW8QbwAJMXODpCbz5c8CQpFdoDkHVLGZ6UIx+RjqgNkqgwJ4EnKngTsRrIWoAm/n49rxKV2Iph6I8TvxZgFGB3jGWsyCINuMolwITuxMqXyauWpz+We+J/f4wAW4xN/dl9b3C/vhXcth+s2EZ2aYWtQig44xli1x0lEhQPyOnyiQOV6eE464Hgj7Xh9jK3/23sA8SyJEawdVD4cIqT62WtKWSsAD3VVeg48/53a9gFSi+cfhAV/Z69vV4ok0i0UjPm8aM/RLyEqAlSKOR/3FPM43vNzREXB528QFV7V5/NMtigCV53EjOqiWD8xT+Mz+ZPPbi+LDwAAIABJREFUjfUT1x5kW6hmI07k6ytiYvfh4sAaZe9vpSq/ZC+lihr5EPu6dfI7CEXmRCqxT3tZ+7P9ottKXidmfH4GcaVr0oHI1cgqR2e9EyOLRXv6+ResOjohIcPi4pLUihDzajKZERXcwwYeu0mY0EfjyyRm4DN0cG8zw/u2tb0hMBdCHZKCnMiJioatUVHRRVTwHuxl/MxVlxXdd4ypSIsEnERszolKcqae1Ew7yEXWo8Q1EM9G09JlqftQvt65dUNgKmpTqjQ6NMX/O4RFN1GBql7zE7BHvRHyFXPw79GjpHuf0lxN/SNYy/JkF5Dnc7+bqIg5f69PojEoc2lgaPhzREVhv9MTImKAx8BdWXl2ExV8uuI+1Y7tXLv7nnxfU9PUtA9yvWGl0L2X5P92c+rP5xq+v92fqCAnJM49dPiCzc0uKA5OTx8S0YD9EyIb4iUVFdiloUxfoSFpssqQzU/E/d5ekcVSpgrU8z+Zo7wmYilzESUuwBE5MPO4WilaY3fLnn7yUZsYHbRDk0NWNKyG6GPUsqZUxQPW0z9sl99532bmVqzc6+cSFM2AJUwX3htFMbGcnHh+fl4Kd/7E2gnSgWeElzY2FQD1s7OzIl68sndT1SL8Po2uAYvI9KWObXjD4eh1wroHCMYaCdERYiKaTrOmUSOjIqVpNuCi7HF3UHiPCqDF+kPTSzC9kzj8g3xO1RZSZ7sid3B0xO7Ozdk2Fd2tghWSQpt55LY8XpGkivdKVfNF5GSlnHoNUcXZsezRGYwq9gQS5cS68izOY5yOUNEDPDVbIlqYEwDZzBniEuc0nj/V9AK62QuLWEq53Zf3p3OgTkIarIQRsJUqsgwDsOb5jg4PyaO9r7dkly49p+r613/+czXYXphftz//r39ob7/5rj3++GO2vLpir7z8z/btl56TSvqN37xjP/zD71l9a8sOnzhhMzdvWm1zw44dOSKiYn55w1Y3EB5sqS/IN1941h44c8o+/vgTe/Py+7ZF7jE6aZdeeN5u3bxm7733nuYpRMHJkyft9ddfVyUA1ldf/8bXVV35q1/9Uvvh8RPHZNkEUTE7MyfAnH+Pj43a+++/L/KOccOSCLKA6jyeC/NrfHxCYC9zjio6nWv2HNxlXYvQsn2bnZ+xSqVPPV+wI6O/C1UMUnsnsRrCLBFNyUJ5Z7umfIp1jUghcmvfC/3MJVKh5IChzoNUdierKPICcjhAf+01sgJLOZL6A/j5l8TeG+Huap0QtwFhyVNVRdtqyeaLzzh65Kh6LWHDfPrkcVtdWSIY25FDk/ZHf/AD21pbsYLi9p5VBmiE/qEdPXpMJLHOEJzV2X/39uzjjz624ZEhdznYqbl9kxrEt4QTVFHe7zbV08KDYlFnSNY0e67HTYRVPWo+ffXqDRF8EnOoLxA9qSBj9iT28P4bLpRs58P+Fo6JYAmqXlO7qjSB3KNhvffuQIHvjhaqPIL47u8XDkB8IFZyfvN8CGLcewVSGS8kSFhFUWSFcr7ks4Ht9QCOAbu7qr4hjyUeRR6ufKhQVDxS/rlH3ueVUsQMWa6Vim7jnfUzlMiNnAhMpNW08fExzXmuhvXN3GVPYs4trawobwIbwQJqa3PDektFCU/5LPYT+vAwtoi8ylWs7NzeGjcE7pkeoS6iIXZ7s2yAbZ0v5Bbg+BLuHJwzA2fQmQwwPVU7qKFzIvRVbZTycmyoqKig6sR7hzQ1R9h7uCbWkM4mrBPlmjiA+DmR14RLQBxidV5K9mA8Qwfy3bo7cumwRPY8JAk0Uz8M3pfXT0yM2fTkhPVXStaz37TtjU1VLN64dcf6BgZta8d7qdBw++OPryh2olhFOCOSBexMlZ1BCkRWm2VtYe2c8oL2mbztD98R6Hne5P1ucciQZW7Cp4gNxCf2Ofa7yKW5aWIEYlo1CO/v88oSequw//S6NSFjSJ8pOWbAOh5odu5CLZ5BWOEzxswJkT3qI+d5TeS9kefcLztsi+2SffGXvT7eR7nkV9ZP90+6v/rJ7+YInCqjzHdlv8rtk12FDltJeYuCIvpAsFGyUbEo+TvsPYlc+J/vw5LCTSRmloDuDYNS8An7nMxzV8s8k0nTfMYPb50xjQIKLdiMBGlfl4JB2MMk+6oEIhOwxkZHXQVFg5zGrtEQh6AfjbJ5jfv/9Qn0UPIFYw7pwKFkc0MJghpa7QAid8qN2XDYzHkdZXokdBwoSG5RkgAiUdIp5YHK7lreICn56LFBU5HCxop6ZWVpSUn50EDVDh+etpWVZXnj7ZIkyKPWm9jxNr45+oHKx8ZBLJQUvrm7ok7VC1JLuNUFSTdBP8DzdpKIcqlSkWICUoH7kieuDqjeRyAAF21gOiiQNAYpsafxlX0P5IT8ZUmeUFS4b2X/hPeoCKDKS6mTVcOXEhU0Yi6ox4MSGcbR8zhVf2izwktQpa3eLFYAXonKGK+oqJQpd+V58TwZF7cecGLHyYp7VVTkmwx/Dx9nxlHl+qHKSSotJSkJXHXrJz+8M8cY2/GJEesfqGptzM8t2qefXjdIFMCNAFujCTHvBVGBku3fQlQcAAQy9X2kBhwouLZ8Q/Tfia5WPj5BbgW48oUVFUpQ7/WlGi0vs8TPvFrV83frG/8ZBJnAExQ8PJVkJ9FdTdEmH5g/qWlvPKcASvJNPOZ8HFQ6IDeARAdAy58dpbw5iJZXKETvigChY04rsRcA6b7XAbTkYHV+XQFCx+fE88pBrG6wO+4z5krcS4DKAWi5escTXE8Q3abp4DU72RdzICcYpLRPikV+HtUUfP6BCoGsosPXR6p6yta61myWZAZRwoGUZ5+TATEWjGWuxpWtSFJrRUIX75mDdk5UcGjyWBFJLn+2GwQmi6oAgqPqJWyIBEBRPp5snoIcYc+Mzyah5ZCJNYVK69NhUOX2qTIFQCYH5gXGAtCmSjdZG6R4ClEhRXmz0+8mJ7D4XT3P5Ms7RNVEUkSHWl1xMHk+x/OLZxL2Vu59689cXsUJlL5XpUw3mNo9zjGX4/v5nMyJiriGmDt5XAqlYHyPmLQn0hIFoKuZUmhVzlJFPak+Qg7uxbyP+ZLPvxiPiAk5UeH35vYeEf9youLz95ofOBxEiXvMyQwdhhrsi9GHxqsofA0kO7DUtDMnPSLXya8p5m80+dPrFZ4TGKCmy95cm6af5x9/0rZarpCbn1uQCo/8JdRmBZSsKZhiTUPul1dUhOikm6jY2FxTPjI0OKIyf8gKPoNDHn22cqKC9+Or2/qJ+woCV+vWVSgHrJ+CrAiiIoD0TkWF9wnioLuxue55T6NhM3du2cbamtYS1xL7hYem/3iyItaFYi9xMhEVAD3Ju+E+e6ATlJH7dtaB570RZzQfybklAunYLXWvt/uRFYBCfAEcjI1PJEsdn6/dREXYeyi22UGiAjFI2NmJ6ErkW8zbWDeRhWL9GfckcAXhRephFK/t3p9zoiJfhweICjWU9spb5QyqqPCxPzF61g5PHVFPhrnZeTt16rTdvH1b5KbOKwILCwIGsZ/xlJkeCC3lINxf2LGql4F6vwD+UQkZhKiTB0ylUCc7iNe0vgoAaM0uPn7ezp48ZnuNTatWCrazuSnbi4mpw+rNsL6xY59dv2OXP7hGWbqqJa5fu2bHjh+Xqpjxv3HjliGwoQIckdKZ06ftxo0bOlcAKjIGU1NT7eo9SAzOGKxJng35OmcJcnO+ZC8isM6t5jSGab9pJgAToQIiIN5fQCdK9k3IGAcG9axpUjsyrFyXNQwpIWIdwK3iIgSs11gGxT2v1qcKf2xiylbW12wLP+/9om1ubQvE0nkzxAJclxTQw7a8tGQTkxPu/y3bRxrscgaD6PTm1YcPHxZpEJUWAr4h1lO1OPml+kgQ26jCAJDEUx/yTw266wK4pY6l70oJAsftrahy31jf0LxhHH0+Alb1SeWPUI39iIol7peKrloNIqFmv/fSt0WSvvXmG/r+wvyS/eVf/pn9889/ZY89dkEN21977Rf27LMX7cSpY/aTn/7SvvPtZ+z1n//Gzl94wB544JwNjo3Z9uKcvfn2u1ZrmNVaBdva2IYNtycfPW/TE+MiKt798Ipt1/dsZPKQPXnxSbtx4zO7evWaQF8aaR8+fEj/Rv3OWoG4IOem4a2TcUUbHRnVeXZrc8vV2P0DiqeM1Qg9FKJCTT24vGIT8I5cxxtRo7Cnd5fbpwIoQ7wxD5v7NIVeld//xx9/pv0aAFzg+Na25g32lKwvgF+voChLgY51W1SIeqPb5Nmg3pRuSxYiQs2/EmA/6nUIDgD9im2sr7fFOO28GICYSiFU9Ns7ej2ALGMkG8OEh0SuS2Pygb4Bm5qatLn5WVUfUA2wMD8rkdwTjz1sP/jed2x9YQ6fAav20RPR7PIH74uoGBkZS5Wg3lOKtUXV1vDoqK5PNmX0j8KGOzVnhkALm74QLXD/4ASA8sS0a9ev28rqmj3yyAXbrTftZ6/9XPe120hn40QC8f7KRfYaIp3iDATJwBhFJZ2elxoe05B616i4y3OjOLOrjwfrR5bgnqvynFywWbFSGTyIamsnmOmLBUmF/RPPiO8Xi/uGxTWVelHZzPv29bs9JSAv1+y4APs8FmuVNokEPsE+xFjIelsE7o4qEQCb1UNLfa0QJJZV4cj7MQ+pLOR500MEIoh5gN0UlWlq6l7c8/hVLNvdu/NWLmHN5IIm7JCIFVSNVKslxasG5xbA6323mlaYbHoTa8Uk2am7aC3Ii9hrXaRUSWIcsBTcSqJabEhELbN+amrCTp06oftbWlq227dvpyqp/IwFcQEBx34P/uQWmqxJ9U1IDc35bLcudss2Afci+FyQ1+5j2D6ruahGFrLkszpbNNRf9dyZ07a+smSjg33qu4NzyfzisnpR0QfK8wDs93asTnwv9tgMFtZ1fkZVbDlbxx3L5lwcmefUkQfn5712LhRixFQxIqIm9Q4hnlFdPjw0KOEOzdL5OcTpwOCA5gkkvEgKVQt6TCAmkt8Sn/oGBhQvdpJNus4yEuVBiHkvC3IL2VanniPEJY17F9ES+c29ksPI5eI8H0LE+yaSXRUaXxEVXzRSX/3sd3IEThTLKj8kiUUtwEE4lKxRug+wQcJMYkmZJMF9dnbeAyGlob2Ard6kcl8B2xs8eTChvCvznMth1lTqJpuR9CXFhCxkQlnlP4iDpsoHw0YCwC0RJ7yFrE1oPpTU1/yeWFuA/bSRwvxryymhqKknz0Qv2yOQsZlFrw5nUmkG5apCEgcCPxZMbEokdAr65huQb5p+IJO9jxhzvPad3dahW2rCghJ9+UL3VdXczMsAUS1Rvlm02vamDk+bm+sqcaQ0mkoQlXVK8duna9C9UYqXGtIxDtyjkh/54XsZLAGWLxIQxoSNnHtFSSTyJBEEvJYk3WX0JAmQFN5IHK9HfT6+x8lnH4sonl8kJu73upsaz6II5lDL+7hvJQaQA5MO2vt7OKAZoNJ+8l2MA3AOPsn6ST7QPZp3UsiSNEEs9HgyE4cwVJWAfwLgSJ5UPeH2TiQ83A8JFGMt5Xuy40C37yCNgwKQK7ksMgfW/Jo9UWDTJ2nPm2kHiMHc4HAQQHMQFaNjw9bXjwcuDR1X7JNProlEAWRRkpYAOCkY9lo2e+euDir3Iyo0CPdQJMYY5gHqwH24G3Vb4Z+DD774Osr//P29mTbP3u1kvEdIbrfx+SsNABCf22j8KGGPnqMfRLAgagP1JIepJwXPWfBOZuESgI6aVqUS5bjGHPzrfm45iOkk3sGS0/Z9kmS2HOiIBD8HvON+2lYXWSyLHi6h+stB/e7NIlfLx5rgT55dANysLZXhpmbAce9K5ACOkpd7DprG3wV8111xFeB7vLeTPZCJXgaeJ0bM3biOmOcxFjnhkBMZmm+pcqybcMnHIICq+F5eQdFdBRGxItbUvYC5Npgue9FEWiYiwg8/HTutUO/HuIe9GuuO9ZlXm+RWE4yFxjIBLE6mlRV/mUfE1Zg7InuYD3o2TlTEdYtsYK8i9oYHfFZRoedGCX1m+RTzjvd1z2FrW+wEUJ8TFfyd6wwLw3iuaoqYemvEHGKvz8kgAXsJGI37CWAu5udBcD1XQflBKycF8pgS1xFrJ4B+YnL08pAYooUXMESFxweq4nQQU6l4wwZociju1PcSxt9JnGh05z/rjmdcV8y1IOQ81nfylJiT8fv5mo/xCDLG85PP37/2NXISAea+p4QSPZS6avqYAPR8TsfrI945SIP9ADlAM1nmONgN+CrRAN+Vpc2InTt/wQp9gwJGqAzlYEiexr3XmZdp3Ii5qOqioqJaqlhN+7TvyzGvPF4hvNhQ4+C+6oDUt6ifA9DZ2HBfaUAy1hBrLGIGABRfso7IiEqNZfo/5nqsSf4ty6iW5xtBpqkhIl747L+FHlVriKZBfT5711aXlnydtasSItomCWna6/IY7M+v8/Pu+Hyvf8e+GnEnelQoRiCCAVz7Am7kwJ6U4pX2v4yQ8Ofr7oMABfdbUzF3Ds5XAqELhaimmZw+5GIdeesD9kePCCecpV6XkrYmgrBdUUHelQRCAjcyoiLftzQO6dq1thMJiygA8M8FS/7Eo8ooBxxQgcbaasfyNA89JytYfYfGlT6uDnh5jwrW/qVHviVLmycvPi0bk/fe/0D3izIW2w6yFSqMAFXxngYwdGBpX/HULcNQGCfLVCkyPS9wcNDzPM42KrwV8O2NpgGwmrVNVVI8+MBJe+qJ89bYWRdx4daoBdva3hVZYcWKXX7/I/v0+owNjkwo18Mrn7MVZxi3CUHsNGR37txOuYfvaQDunmvt2Ynjx9M+tG+3bt2UIjhsWziv0ZB3r0mTYK+QYN0Qd6iGCLBeUaNgNqam41u2vrlpu6kvUiWRkMwd+sCg3oVnRelO42A17W62ZItVoxedQDesNsyGqASuN5IwqmDHT522heVlm19ZFgB4Z3bOjh09qs9GzEXvPOYJRIk3i93UmROSgxhK3h65NvstY0ZeL6ve5KUeAjOeCacU7ldnk0ZTBBCWO+RIO8k+VdY46YzGGYs5AAiNNQwV+JvrG27fFnaegN+9FZ1/OUMMDUAq7QgoLZeLduTQtO1sbdjTTz0hW6Bf/+pX1lvm3Ldr//2//1d7+eV/ki3Uxvqavf6L1+3iUxel7n77nQ/thz98yf63//V/1zUcPTphl77+nB07fMh++atfW2O/ZI29gtV26jY00GcvPPO01Xe27OrVq7a4umHF3kGae1h1oGr1Rk0itGgQHVUn/ImtjgsgGjp78hpybYA72dbJFjS5K9Tr6ksiALrRELBHI2mqLnAKgCSbnj5s77z9dqpGgnzaEnEM2Lu1U7MTR4/Y6TMn7frN6zY6Om5zc/NyDaDXBcprzeXUPwE7Fu59YmK8/RxoWA+Z4edxr7ZgHQMoqllwIrhYmzyTEAEgCmNejE9M2OICJD0q/JLvGQkAD0EJa5q/c172CshOBSuTk39z/pgan7SRkWFZPxEXea4rS/NW7inb97/7dXviwsO2OHvH+rD2KdE7ad9uz961w8eOWUO5YUUEQKNB1Qc9JMr6N7kZQCkxmefLOJDnq/8B1tFra968WQRiTdUFqLbVb6zZspVViJiSHT123K5c+Vj5AT1wFN+TLZ7yJVwNUp83MAAXTPpZDVwHfIC9m++Ffen2ljcJHhoaThhDzQnMtBdz7cTkaDoeexP3DwbAemVtQjKWenpFXvFcZLVcoqq5ZP38DIwiqTNYf557uUNGkClUelENRmVXNEYnH+BemCME5P7+XsUK5irVJ8xbEQWFfVUT4aJBz4/1tQ0rQEg1vTKBMRsYpC9Rv9tGNWoah0ql3xbmcdwApyhKjAReUCgwtjiOcH2MN4KjZDckUtzP6Ih1I4dS0/GiyX4qP5v4fuMN4cF/JFhN8Yzn6j3nvMeC4vT4uJ0+fVp2VsR1Kprm5ufVNyzyV7l5JGtGxeg0p9V4Pp3XZdGlvm91nV8kepK9NzhW2Xsr8HuJ9Ob65LASwHyzYePjI7I9K2IvtrVhO5s7dvaBs/bGG2/Z+NSUyDfWLvgPsafBPtlbVT5K5RP7xN6eV9RpLkqg4b0ldaaVsNPPTN25Wp47tfNvaXaS2FD9RMoi5lR53mwpJ5iAkMIGL53n2Sv83EO1DXhiUXFJ55cCFtxrNjQ84jlLT4/mGoJdYpAwwd6K8DLuh2sXfprOKF4NnvrpdBEV3FN3Hhz3mGMT+fnlfq/vPn98RVT8S7L3r17zOzUCZyruMUwSEtUDYmHlS0diWpSyheA4C0DP4l1fs9W1df1ddlGoAtUcx0t9lXAKqPBmY17scBC0zKgJbVKh7hXQsBeNzVJj7LY61xd9W+2eVKkR1OIwrcOLeih0bEjY+LkGghDXX+n3smYUQ8Q2AhcJHq8h8OjwQhkkCYOaPW26UoMSzbr3f2DjCnsTgD6UIWzaG5sbOmxwnQRo7o0xZDNhIyLRxz+VIAl4wAa5urKmQxPEC9ZJbLIQSCiiCJocrDYpgRQx48owDuaMlxrsASokEICET+BNsjaJ3hUCE1MDw1Aut1VHqSG3l8J6KaOSAhonqgl1ScG4UKBJWbXdOEhl71I2ooyiJJLEnkcaDbQZW5RLTaRWqqzoG/dnEeBjABTakLoqKr6IqFAyxrwDpCm4n3l4Fankr4cmklWNQ08ZpQcJEo3BXH2r6gWePap3TUjBBAeICini74M2REMqrpuDE4QeioduZW4QFZ6UVLyiYq9pY2ND1lvlULwvooKKit5Kn4iKHIiMjWjm7l0G875EheZEer4BAvK7/98RFZ1QGOuftUDCBEETFiChjlQPClXHJKunVKIalk9hAeUlz50qhwBbo6oo4kEOpGrD94FsJ3Q5UE8/gFCJxrW2AbOmK/0dgFJb03aljGJNF6Ab18MzdjWmN77u/joAbqZDV/6aboIjB5IDWG0nNfchKvi5DuNSkXlTYr54r7x5sSfP3nAwB59CUR3gbhBo3WMc45ADTzFvYzzjNTEn2S8E0nPoTA3PeN+43iA/Ym8IECvGKMY9QOcAtyJhj+cQSaHKqZMFU3jv87tRah6fzfrMgX/16klVDJoDifwIJZmIxNTXAUAkrl8xhhiclNOeiPv80/9e3qJ9VGMjjh+Fpu9bVKTlREU8l6j+IEkGjHEVG1Z8BwnFGH/2Lt4viAbeJ5T58bxDqRpjGmPf/ewUc1lLab7GNeVJdNxjxKB8PnFN3URFDvgGQcTvClCRZSCgM2NHg/JYhw0bqPa1c4tYYzHf7wWIx7yJ5xx/xj3GetR8SX2uYgwPrNV0iAoypvuAceB9U7NeXy8dooJ9OA6ncTDjNQdjVqfyIK6RZ8//moMBYgfUT+xHUFAo2KETJ+3omQdluwAQBVir6odE2LFfRnUcognej7nUC+mWGstyLZ+zfsqICg7/3vfCrQAgDLxhJM20+5Qn8MX6CttLr+QC9O2QQlrXaV3E2lIqwHuurhnihSApQgHKdYmcLhT1GioHIF2WFhdscW7WrScz4qk79t7zoJu9KCxHvyiZvx9RIfCGZwS48C8kKrr3Kn9vr3LjPiWuSVaB96pii3l6YL66tFOHd7zLxyenBEqRP3qzyE4Wzue5PUgSHexHj4pUuZBsOFTJJQsej1mfIyqigiz96RW+e1Jsui2dnnayGuysB8WVBK5EnM/34cj5701UuK3eZPmwnThxUg1sUYljC7O0BPAH8EDMLVhvtc/W1zetRn8lLFJEOO8LpPB9ppAaf3sjWj0XAZadynGJohIJCSjGmGHNUSntW2Nnw5568oL1lc1OHJtGcmJbK6s2PDZmpV7sXCDXynb5vY9sbnnDSpV+vT/nBCrjAM+JzfRd2a7VbXpqSv0qTp86Zbdu3dLZgWcAuH/69Cnvq7C/b7Ozc7KOkmVRvSGFsBqiFr3iWs3T5bPtZIMArLQfonalgSj5Curg7d26GkdDUPDM1te32ra5ssPA610Cpx5bXVrxyldEQL2pYn131/sH9fi/GfvhsXG7Mztju1jHbtd1n5x/sEPhbEEgZ00DdjNXeW8BflhDCfjx6misiAJkJc8mphEnNJ9lVxy9MhB9eUVl21I05ULEOURfEtpwNmCtpT50vJY+PVJaS0CASn9XNjp8LvcKQOggaUNxhqoKt8GCUW/ZSy990zbX1+z9y+/a4GC/mrT/6Z/8ib36k3+2l777Hfvoo4/s9V/+1n74g++o2vs3b7xt3/rWJXv1tdcEbi4tr9nJk0fsR//pJfvHl1+xxdUt26BB7eaOjQ4N2n/+gx/ZXmPXrl+7bnvFklUGR22zVre6Ghg3dQ6hgo65Arh++/YdnWVr2zt2/MRxPcvbd+4k+yPvIUNu2IuyGuLNDXv8XJ5sfR999FF79/IHTsy0zM6dO2snT5y0V199VbkH5+KwImLJAPxPT03a1PSELSwt2NjouF2/flOAK8D1xibkuAOhsVcPDQ2I2JI4IeXbvt+nOJWs/CSClG1iUfMI4hxglZjNXgNRL7AVQQd2bQl4ZJ2pkr7EPINsKvt6aXhlgVt9eQ6lfiuyD+Kc7eNx7Mhh79i4R/UUll537fDUuL307RdtqNpjG6srNtBbFhGxvQupsG3Hz541o2E9Dbx3atZf7be1zU2RCwDU2Hn19fd5o+J9ehVuaPz5fPZt2UBVsQouiJiTQFH+ziVVPJHOMw/584MPr9jM7FzqV2GylSI26PlybiyawFpVZLWrnwMIdrKW9QSBpd4FSXPGOAl0TSIn1ghxgXUgrCeda3lPr46AjKHSBlyH/j9l291FQR9N64lJBRsZHlKVEPFUZxFsppIVFOSf1r4IJHdiiCpUEbmJJCEHJm5KJEQPHQhnzb0p4TmQryxNb0K+Zb2MZQHsxavMVW1QKto2FUfstS36nwDIUxW0a5vrkBYIfuLzse6i1wfNzdkjyOO5fvqBeINokf5NYRAgAAAgAElEQVTlShLwJnGGqmqTA0XFiRjmKpVjrAUIKV8HVNxgQeSOHL4+wCt61O+Hf5NXjI6P+R7X0yNbcbCZmbuzwp6YxywZ3gfbMtaickvFP8/fVTHSU/Sm9UoafN63RTWpL0Vzv+VnGJ0hXbzka6uhqqJDk+M22Fu2Fg3FOVsVS3b77pxV+wdsa7sm/GxsdMSuXbtm/SND1mjtaY4yZ90G2O3VdMFtokIX1F73kRfH2sxznTw/8+nqIAJrg2tm32bc+ZPqMubRINU25bL6V4mE5mEqjvtZ9MjhQ7ZCn1iRPElGtF/QnohNFPEiRC1OortohrlDBWAQ6jqLKAd166f8/BF/785DI/fpPm90n32789L89V8RFV+UtX/1s9/JEZiqJ9WnyAL36mdNscBI6GKBsejY4NjtNra22iCXPAtTibQSvyJVBTRSgzEn8eGAAkhIoHQAwM9clBlSduaeiW0gRT0RKONMDXSTP7MvRA9eKJ7C+oJrli9iUltH0yclGKqCqLhfYWqww791SHE8Wq9xlZRbEIRCVoer5EnLeKhCQeREXRtYbJwKmrJXMvnfUZ5MsFdvAZVx7ui9Uc5QWkpwDjVulOmx0aBUIUjyOjZUNgWSTF13C5sPmlS5Oo7r5+IhCALwEtCV7CtCVRuAr6tE/HAoa52UpOSHYxEeSd0ZbDKJBgz59Ru3VAlBzBUYnt5Hz1SdGZP6Tokk/7F5O1ER/0NY9cizcs/Kw04IqRolAZNtcCuVJ3YSKe+DIvCIeQMonCoqVBaKyss/sW13JWU+z75ctl5KarEFyayflFSnZmHMgRbO3ton3UbD1Xve3M1NeA+qZTsbTqcSRNZP2HOlRInXBOgXRAVjLKsjERWolIaskhql0aPis89uWhXikOZmKCtSiXMoIiAq9r/A+sn92wMEcCAhriPfyLo3Pa+R+bdWVDhwe6+KinwTlsKk5A3X3EoHUsvJTeZn+AmLlMhUmf5E/HnmRIWS+UjAEsgVT8nto9qYSBvAzROeqFJoJwYxB3wiuA1RiwMch08SZk/wApwMwDvuMQc7Yy67v2dq6HUPFW8AtvdKvNpzPmvOnavlBRZnpMv9KioC6OaQ4fY5fh+qAEv2T5rlqTQ5v594XQwlc1sHiBTD47oD0IwxzYmDfB3rGSYbKQHLIig6vUNYQxEPghhSPE5er90AVk5W5T8L8Kwb+A2LQwAPKZV4xg380ynXTQB8UpTF2uWaw2YgKknaBFZYTWBlk4gMEnN+NyykdI169skKK+2D2qdIoBOgJ2uzZH3mzYVVj3OAqIhnGZZP7GXdlRAOiPvaj78HiRrxlrECzIjxyAmxnHAK0jNAyXyextj6dR5UB+XrLAiuPP50ExV5pUnepwLfYMAzkd8ID1ARkq8kxTol/l6w4vMqJ2JiDGKddCdncQ3x3LUGMmA7xi+f4+33CPAyzZmIs20CKgFiAj6TT7JX8zi4ouq9pBj0e898eoULO0ji+n7PeaLqVIRZEI/JSx9LhZRUGaYrzKvegSE78eBDNjY2KcAD4ApQLHK12NN4LrJxSc1qg6jQeor+CG2Ryb4qPKmcoJk2RAXKUBF1rZYAo6hIYl6yz3FdOVHBugul4YFnksg7xczkS0zMXaOXgEQTbq0Z1k8AARKiFIpSvZGDoFzfWFu12bt3Vdkaec69EvN7ExX//oqK/ZL3C1PjXg60+V50wHoqtzbtEvF0VRjzeIPW4Xnle1cnF/E9r70uI19mPLWf9tjI2JiU5dgtqNLXOtaMzOHcsq6x5wB4eK3JfhHVqIAj1KH3JirCayvy71hXUVHh497JUQ48h2QXFYBErF2PYw4a0oeku6JCPSqKBTsxfFZCkZMnT9vi8pID31gDVQHFIWBasqbY3N62za2kyk5AOnsRoitAeIAeEdXaqxy88ipiV7fyf1Tg0QAbVW8Dq5QW17Zj3/r6c3Z0esyK+3UrF7F5dZuNUrlqfSMTtr2xY+9/+Jl9dPWWFUq9Nn3okN2imfbx41ozgKvMewBdzmE0Iz5y5Ih6VBDzomoX73IplCu9trS0KFDIwaZOg9zeSk9S2A+qokA9AGQMzt7ScLC+aDY5Oa4qhi32eAWook1NTyve1uoNqVCjzwXnktXlFY0VOa+ARCmzndiQcKnesCq9IFKF0Mj4hF29ft122OMLEB1YLbl9ruKnwMO6wFVA3NiHonosrDR8Wu9rzx4dHWvvjx67vY8goDygLvcpqxlZNHl2Hz16/PX0ugMUp6LacyPmOQAnS9WbZKfKstTPi/gFAA0AqHMFZw/EePt4mnu1yne/8y3b2lyz1//5ddnd9FbM/vIv/sz+9n/+1H74ox/YlQ/et9+88Zb9/u//QPP1vQ8+tRdeeNr+4R//0av6Gw07eeqYfevF5+3HL7+iHhXbu4jltq1nv2jPP/W4nX/oAXv99V/YndkF20FIU4Cg4Zl63yqsas6cOWkPfe0h++mrr2pZcp/YQ/EsadCuHEjqZa8YrpRdka7KxERq8RqswWimTe8LKhq471MnT2r8f/vmbwX4S0ggMtMFQawRLAinD03Y9etX1cj9zu27Ll5Mnxfe7b5/gC9gPeW9JLT2k68880uqbxpha741klK76E2IeZay13FLT9k3Qaam3oHcPGQFjad1lk/iIZ4t4GNcs+yRZAed+leknL2ka9m36clJm19YsIFqxY4dO2R3bl23555+wi5desZWZ+9Yf1+vrczN2G0IxZER+dsfP37Cq0HAUujToObXXrmCxdnq6rpcFbTPF4vqLwPY6Q2WPZdjvq2tpf4EstMp2vrWlq2sb9rOzq7Vdus2PX1E8+bW7Tu+y0D8YXujSlQXK/En1RvkvBBQIdzhOXB+S2mNhAaquoVcABPS2HpvJN+a/PwQZ13WjfoltLyPi/eppNKpIJLCfzdVp2mtQwwXhG/QkJ5nSCUF94ldGap19nR6eFDV5ARNr+IT8W9oeFCgMjGb9Qxhyf1BWHDvgOhyxqD/zP6e7H4gtMghIWH3zSsK+bxqb8WOHztsiwtztrlJ9UpDlnv04FLLRQNrkpxKBKo3UgZfd5cISA6e0fDIiK2vrmvsZHtmzE3vm0Isg2AVEay5WxbhNYAglnculUTQ0lyd/kkIUhljbNc6/ZOorPe4KLGZhDxeIT4wOCi8iXFm/4BAosE963xiYsJxu+y8HILWaLId+FCp6L0KCf9cO7FRIqt0XmRf5DnofNdq2qHJMRuslq1CH5n6rg0PDmpu1xotq1T79T/xu3+gT5VNxXLFdup1ubEQ/x2ASz3TQkiYNdP2vbaTvUVe0I1ltF+RqteFJ6gCy+cN8Yu4xt8HIeE2NvxM1/KeNppMwjtLNjQ4pNeTgzPf6fMzOzdvmxtbelaMuSwDkzAbYi0EMcQcH+sk5CJPkAPGQaKiO2eLs+uXfT8/f3XntAewlq96VNwr5f/qe7/LI3Cs4Ad8t1ZIIFbJVQFxbEP1r4QxgSrrmxtKZBoAeerPAIvuPvJK+uibgGqODQhQPalVOqotJwZQEhA0iQC8TwBZO7vuFekKL4gQ96Bm86YcVd6TG5vaKCMBU0l7AjAA97lmt6TyXhvco5QxbKhsIFLqUPpHOey+yhBpeMQ1EszYPEkiYenZyFfXlm18YlJMMJUR2Cv19xOYkwIFR6KkNCIg8jsk8VIaaYPz32MXALDvEVjuDC7Bkddyzxwk+btAXDbi1Phatk/J5ilIEx2G8WlM9leMoX4nKZWl2qShbcaoC2RLE1Ze7wnUZ4y0LcPeU8WhEtmaTU1O2BKHlCIlnCRUVNH4a2PzExutswYJrz8vJyu8gbb79AOw8ByK1jvqzyUAqo6KUp4t9wcYyOUg0kLJlxrPJhpMFmMOgEK49bj1k/pQUApZbqv42oflYPHT5ujAXDpIJ+wAsuaLiIoAi3OiQuBXZuHAHAAkUjJFM6de5gPKn0E1LOee8bG9dXPGKiWIClf1kcCQeMSzmZ+dtVaDZtr3lmnuyyC7feEHbEY8eXXE1BNz91lu246k59kN4PjmGFb7YYnlpIbmDwd9EkOSgXRYdKLHdGDVJp7s07xJPWsjgLmk4JfK3wEYB2wdpGuDHun9ojdNNHgPFZ3uIvlAdu7LD02RWGuupvWjqqTsvgRKqgkcSqpOA1/NSzVr90NujE0O5jLP82vlEOB2bx37sI6awlVqMeYByGmM0/OQPYauwQHZqCbgM0NJmwPwOTDtYK0n4epTo2qBpqvfEyDDXFajQOwyZOfmBzyfx2FR48Cv4kEiCUj8g0j43H6H8hpVv5qPpmqBrE9L930E2JYDblKfJJsjVSSkpmihlI/kNAfhc6LmXkB4JHbx3MLuKMB9Hx9voK35IZ/jTqWJT0FXcvL+xDap+xNBFPFY+5cq27z/DHFcJEAohOVTkoglAQBp/ZDg67l3xjuZxCbFvJfwR3wMJT3XlSvMg7DJn4sO+qmSw6+dWNxRsUe8asfxdO+hbsyrWGK+CwSLvk/3ILsPgqT+zjmhoYbtgEPZPIv3jnkTRAWfJbsCStD5rH1Xx4pwS71M8LTW4Q2iIprCp0MC6yeU+zGvpAbL7AajB0QOiOYkS6ytfL3lYxw/j/kV88LJBCwRHaCIkvC413iPmP9BfMV45eRJzMHuuOxCDfZWqS3c9i5ZnjmZX7IhKmHPnLPNrV2rN/etiq86jX2T57hHNbPaDgpLn1PkEk09Hye6ovLIr21PfvuoPMlZOPyHgpDnsrGF2oycycloDnFENuZaVFREhUYOzXuzY5/rDo67+o+/r66s6u8iVisdK0cJVMgr912NjmCCa9/hwH/ntkQhgBQOn6W5mP4elUfdz/LA+tEue5991rns9l4bB2jtK7JoKup6FC/bREXkEfl7dkbBG476nufPJb0uiPMDd+LxozN/XCl/YL21hT2ei3BYpqkr1hFGBUzWo4Lfi9ycOIatTwPQnXih6/c9MEhHz/E6QoiceNQ1JMCS1/ja3W9XVMQ81u+LyPMx4LOioqI9nolsFYDM2O7tCzyWpVaKI6qqkZra7PDAGfVPeOyJJzRvf/GLX8qaAVJiYGBYNmWLS8uyYwBNA/SEfIi4BkCBWhdVN4Bq5IJBFgLmye98tyFgam1tRcpZB/wKVu7Zt71mzZ596jEb7C3auTPHrLDXsK31NZs+fNia1mP1naZt15p29dotW96o2fp23UbHxkQikPtjs8pcV0UFilTETxubNjk5YTdv3ZI6lUbg3O+JEyc0ByAwFpdW7ejRQ7JoIj4CEpPHb296M97JiUkBNOoHxp7S9Gum2vnc2TN27PgRe/XVn1mlf8BaEFgSuXBGGxDwhpe3npGZnTl9xu7evWNHDh2ya1evKVYQ7yCWUUlT3dTcrVsfVrnkH7Zv00eOCFxFUbu0siGA6Mixo7o3WRk2GiLPyY9RPUMwAdpvbqE+77FGzZu4Rx7G73sF+57bXQmb9RxJYGICYokhKH2xc1paWPR7SGcexc1EyHImiwqJ0eERB2t3dtuWn7KXSo23AZK5DiolAMCdMN+ziqxDzL7/e9+xI4en7aMPP7TLl9+1+dkV+2//7c/t5R+/poqKt9962z784CP7/ve/q0qAD97/zJ6/9JT9z7/9O+sHSG427YEHz9g3nn/aXvnJq7awumVbNZqk71hxz+zZi4/ZhfMP2s9+9ppdv3XX6jCZ5b7kgOA9InmPr33tQTv7wAP2yisva07RW/HpZ56y+fkFu3njpgBEr5LnHOhV+QKdUdBLPe+NxIm/2FRxLxAVfOGwgNXYG7/5rdYMX046OTnPnnvk6BGbmhq3zz772A4dOuqxXNYz+wKjRSwkYBXy0/caX3W8F+MsTEEVT95Tjb0lbF65JypisCPke9q/EvmV90eKcwS/r/wsKqALBVtYWNAcJGar8iLtOxGXHKIuCAQfHRmx5ZVFa+zWbHpi1G7dmrMXnnnIvvXCszZ/95aaatNMu76zbUtrm1ap9tn04UO2uLBoI6NjLrRoUA21Y3utgnolQEBgM9ag50F/VX0TlleWbWJy0hbmF9XYmi9Z/exsq/IFHOTdy+/J859YRo6PtRZjcefOrIhY5YdUd9TqSRDWY036QybL53B64N+MFY2lWUvkrdhvyR1gZ7cNgDPWkCihJFcVJTkl+VkSOQiUl32nqQ8LMdp7d1astkOlDIQhhDjnD8gO7weCUJMqGOynwIQA2DlH4TQhwZIEil6BMDjQbwP93tOQ66V3KH+fnpzS9XEvvBfN4+nrRBzCGWJ1bc2Gh0dtcGRM8x8x6ODQgCy8/vBHP7DhoX7b2lixa1ev2ubOjgggCP1KGXcNql0KmvvMXSqXVPnbA1lQt2qlV/EP+1fEvTyz2taOn50gTxG4qlm740tUT8gafN/HG0vevoE+CT/4It7euHXT1tfWtTaZd7L+3t4RnkYM9/m0Z7X6rq3xulQpq/HKLIBjLXG9rGnyMpFSsiRVmXKqAE8VROobUZRe07On1AdGVlBO+tD/E83puVPHrFXbsl16uxgVuVV9NtVdm9sNK/X22vDoiJ08eUJ9KSC8IaqxfhPZ1YPFlFfcevWoZw+5+YpXIXd6c8VZ6ECuln5B4sW9lnATNa2HrOqFqHB7Ruzqwjo73BdcTOjNzhHsTKrRulcFL84v2KnTZ2SthRMHuBfjT8xURUipR3tUnK0RFHvPHo+ZrA16VHh17hd/5fl9fpbtzvvvR9J8RVR8yQB/9ePf7RE4aq6kyg/jshKCgeyrWo3mdQnIYlETKNTZXkyxlwACplNp4MC4N9+FnWXhSrVLw+IEWuigagUtcBQUcZCLww7JRKVK8u+Mq4gQkqxdEiT3jGRTYFML4kQNnTMAQuW7lBJKmb6roBxqIxISgrv6TQhg9woPknh5wLPLUsrXV9WBKJQIaros/3w2aD8UquQyeXHjXegNilyNxftDdOgAWK4oCLv6yIOgFDsQKBAyvZSdklCgSMCSigBbUQLgRIWrMVXSJ7/JaA4bpWUOngUAqIbZVCyoRNMtBNp2RFENkdDnBMvrfQPwEjAgwsJVOPi3uioDlbkn+p6YJk9fvBj3IaW8D0ac8ZykINHwagcUwmx/1TFPbKWuViNCr6jRV7KmudeqCtUJFRP0QlE5awL9BFr0OLDK4ZPkCLWnkllIikJZSoH4ah9W0je6/+3fZtO8P1EheDlt9G2igk03KbO0wRa9ZLfM80TdMTIin8vdxo4NDQ9YHwogK9jMzILN3lnw/hkpKYvEOoC2xYV5a9R2voCoONi8Oj/wy+UhKRZDLXw/AO5em2P+XoxM+98qCXalSA4mC7BhnqpnipcT8yycxXIVWv7F7wqMT8ryqLDInxd/V71VVO5kYKk+Oylx21yNX2g8SulHQ/0c1x9/kjQyv6RWJs7Jesfd33sQbKWqjkia4vdEVGSWPqxdfuY2TcQW//z22srtXTLwKcYung0kX/xefFaAxwGIxnMKEsPBFe/TQw4qIH7XG2hrNgPoiFCN8mQnd/1nqWopqlkSUBcqfJV5p0N+/twC5PV1FiSJg4xxTwILUqPmGL98HPXaRJTnwHznvg7aa8X1erJ5UEmsEJI8WfO5w/tKzVSp6JDAewsgQUEatl6JdGfviLGX0jw10/Qk2Q9mcZ1x/7yfwFmR9l6x4KXqDsImvC55nnM/7jcfCvIghuKavXoDFVynqiKvpIjx1jxLpc3dzzL+He8dlXwxRiLEk+LLFb9u65ETcbxW9oCaW07m5PEjnwtBYuSESDyLWN/x7PL1p9LsNKY5UUGVnPYdKdOcMOVQpz2D6yh57oIoIuIFVYFOPDrwHYRdqAEjL8ivVYBq1ifpXvP7fgeE/LU5SRdzCmBFisFkKxHxh9+L55KPV6zt/H1jrbTnZNpzAExzoqIdF8hpmHc9ZoePnrTeviFr7Zes0jdgTXNFvKoTE2DHXOUr7L8aiYyK77VBaaovNtymAHABewIOteQZ8nveXNcao2oOn3l5/WNBQP+z9XV9RhBF+TjogBnVYcTwRKqh4AdAYSyZm+REHDxl1yLLNPYYqjw21bxSavjarioqqPooSCDxbyMq8vHv/vu98oj2GJGzpV40B4ldBvwgcXLgfQtUBn/euk3rxVPq9leQ/0EqRqzN463/PfXpYG8FdO4bsLGpSflzq8a2y/op+qoBZFBRoZxRpBGEEPPVAchQwcczzONt5OTt56vnSlWN58KacwlUjvge8Ug++anKOWJQPqeZs63artGoXIICqjv26VcBAGZ28dwlqTUvPHLeLjz+uFSb/9f//bdWLEJiVezBr52XKv323TsCzCH6NLdSDOXKyEUBYryfi1cKicBO+5egm+iRl+y5+B2yh1IP19G0P/rR9214oGzri7M2PjJgte0t7QdT00etUh20lfVt++2b79gn1+dscGTURkZG7caN60Z1hkCuWk3rBRCH66B34MT4hM3Ozqhqm1iiKt3+fq09rgdwD192nbeSPRHXpTWahBCcNRCP7GxvyfYJQAZrqIcf/po99uTj9ouf/5PdnpmzQgU72kHPIbCC2tlNPTMG2hXZWGOcO/eAXb963e2VKBtQTzsqswvWi499T8nKAEbNpo1OTNrG9pYtra1ZvYHNTF3WtsQSnVtSryavhqBRsp/NAIZK9FSRN7rb1BAHGCP+rlwr2SeqUkRBEpK7pe8jEKonwJuzbADYWlcp7vgc84bbrF2aaQPcQ0S05zGWwLJj2fO+ArLr2Td64UHMsOPU6k3rLe3ZH/zo+3b27GkBpWsrK/bRe++JMPj7v/up/ej3vy/A/8P3P7U/+IMfCDD95JNb9tyli/Y//sffCpwFzH744Qft0rNP2ss/edWW1rZtfXPHarsN5aFOVDwk26Ubd2ZUTdHi/z3sbgs6owEAP/zwQwLa/vEf/0EAPcDz17/+gt2+c9uufnbNP6vp1Ql80QPAeya5NsvPZ/Q6LKkS4623fptshFr20EMPqXfB67/4RRuM9ibUkLWeW504QXP4ftvYXLOeYsWuXPlEc1Ee+mleMFcRA8piin4lNK8teqWDnktrT3OAtcl7uhd8VG64CwS2bdqzJITw54rFUW795PmUWyrhL89+pb4VpbLWHdY/NCkmd3bnBxczqRqjXBYpx5pbWJjT+hkb7re15RV74rFz9tI3Ltn68rwVWnUr2Z5R+b62vWtPPn9JdoQL2LIdP26Ld7HOLtra+qYNjYzb8NCI7dZoyowt1Jb1D/XZjRu3bH5h3hvN15saK0QAA0NDDoJaQc90aWXZ7s7O6WccfGnuDph64/Ztxw3KZeEkNE1HzS+7P+XhNKTeFabCc2LONFRlQK8O+kX0OEHEM2Rd0w8GJX1fn/Aa2SenKguuJ2J/VJvxHizHWm1b7+nPhx4I3rcUzIT+Dn199Ozo9QoniVG9av3okSMiRdk7XRjE86q560VPUQ2cK5WSnyn7+62/t2qb6+uaK4gTmKv05lGvlXKP+sFQ5QFRgQXgyPikLPTIX+jfs76yJtuiJx89YxefuGDDE2NW29yxjc1t9bNYXlm1BtUge2abWzX1Z+E0ODA47M4YikH02dm0Q9OHRSYQg7e3duSOwdhTfQWhwb2wh8rSam9PVSMQM+BJWDYxH8C5dP6QEKGkput3Z2b8s2WFtacYdvT4McXklRQ/eS7gTWALWDrShyzORxIA9jAW6+2KI8ac//0cEvl3qqxn2nOdbBZaTe6cQYzDslwk5r7Z9HCvPXjmhI2PjVi1XJJgZI2KkFrDWsWSbWwzb6o2feSwekfttpqyhFpb33CRjYraOthgEBUexD22hzAsxyTi/OHLM5e8+HrV3oH4OtmZknswV3geEFuQ9lTw0DNHzcpT3ECgAaGtnisSiVYlFmDNkJsRMxgNrp+YxLOEZPSqNHKchveuSD0fo5rJc/QvyigP3kd+1viKqPjicfvqp/8/GQF6VISyUAqTAP/YpGiMRsgQyOPA2U5tW5UUrFjvl4CazwdLTa9SEyG3dEK5ZEqGVDottp2yUg/Yyik5vCSv2CjzpZFfXqXB60jW2Rimpqa1KbAhxPGNzU6HndTcWIdGqfTcr46/RzNjApMrqUoiLEjeogkXZYBOonhSwH2z6bGJkMgAWDFWS4ur2hBUHp4aYLtyACXtbruBNomDAJEiik8/UER1Bwmub+qpRDD5YrPhE+zK5d6ksnblAIzv1sZmByhinMveANGJCAcHAyjNAY/2gRJFEuRFApyC+e2ApEnNp1I/lP6Uv7m1F4kPhwsSJw5KUqu21SeMvjeWdubAyyK9Qa/bP0VFBcB/edhVbN3AZnqI91158iFNFkBxvxxeBeD2FBJw5U2yXZ3j1UJoYvg/AIaclIiN4HMbXnuz/NcRFaHO1vqQatB9N1F48RyGRrBeKFitvq0knoSLIbtze8aW5tf03Ms0Zkwl8VJCJOCVRm717a378/P7n++DEADKv4eoiISge9z075Yf9v0g4HCKv86sZ98t0Pg/AO8OqOJkW3zlwDVHhFRT8blEBEjAVZSdhlvdoHibRMjrRjkgqVkOzyUBJlmS4zYzkKBe7hqQEu9VRvGeV0hkhIdX2zhoEor3DmjvSvAAXQ5UDt0jyQowV0BIwcHtfMyDqAhwPOZsJKL8GxBSCT6qOkBdxWZPOF3t6yRK/E6M/8Fnl/TCaY2y3gEG8nENkCB+P0CzWJf5z3OiIuaHEzkH+2EE0Bsgcn6/3UC+x7d/GVERYBO/E/sA10EsZr0GASNSvBKxI1mb4EFa6djbxP3Fn0E0cLjgAOHe1fUUI/0QoMNvFIrJC9ZjQU5eRSyMcfNrjviZr6tOb59Y2wdAXxFsyToqrZEYa1WqJBBaB8BaOgAm0ibswOJ9Y37lFmGxZ8f9d+aPkwIiXxLxHM9Xu0NmrdV+f+alvHs79n5BaElZTuWVKvHctkyHhUby2xVhuefPC+CaMZWftGPrDF0AACAASURBVP+eLKPaxNp+Io5SxYusLTxpidfkREX3QSGPL/fbnGK/DQIr3g/AXs38EriZr+d4bvnndX9WxIR8zce4MhY+Lp0v3Q+oLWT3XtNKlT4bHpu26sCISvHrew3PQTJ7PdY31yJLtKxHBe8qcjnFKsZ3e31DPSEAV/FA5/ekYqXxNQBDE6Kir93knesnLubNtKOy5sB161lwIG66nSQ7dqEowJZ5yvro7fMqDXKRqF7gwKwmsWoCW5bQYWFuzpaXF22/hZDiIFERVSRfdgDMaho+98i/iKhQZUcSzbhSMD7/P5CoSO+ZVz1xkd3zyOOAWw/ROBvxDE0uexDpAK7uH7R+Yi1FXGjuHyQqCGABijvp16moyFWO7f5Saa9lHJX3Zs2070VU+J7nthN5XIt1xfd79grWwLIOZWvKPYEOaJbK3Dwz8ZDA5AsXLujPw0ePipB55cc/tpmZObt06Rs2ODRsl9973+bmF2TLQlUQ54ElGgqnfVwNNXvpw9bSfgGQ6payUcnmVRTErtu3bgu4Zs+tVGlGvmVPPf6InTl5xCZH+mxnc1WWZGxVld5+a+wVrdw7YG/85i0p5a1U1bzlfEHzaFSbzG3OAFi6sK+gQOUcgvp7fGxUn8eYUx3jDYZ3bG52zg4dmtZaADA5fOSwgKiVlWVViFMBxZhBHmxvresMgM0JVUc0fz558ri9887bdnd+0ZoQA619G5T3Oc3VGwLEAGyoJGccpBDG2rfmvdlYm1TAQXKNDQ/J+olqW/oeqKK4t89uzdxVo+6W5p33N2St+DnR+/GgQOWMwZcAMamuGyKj+eIMAoAUxK8qKAS4dcQMiIJAu4PQ43d5phLPpcotzbFUNSrwulbTa7gWxoj3BczyfdvJ+f7+AUUTSNBSmRzSK/EZZ6opBvp7rb67Y9/4+vNqpo0q+6lnHrcq9lOFgr3+81/ao49dsHfefteufHDN/vRP/9hmZ+7azZsL9tzzT9rf/M3f2uDwoJTbFy6ct+eeftxefuWnIiqWVjet2dq3UqFoL1561h588Iz9+Mcv2827M9bq6bVWEYumhuYa40YcPn/+vJ05c9b+/u//XmQC4r4Xv/migFoUzjyXaCjPMyaVFTBNo3L1DSF3aeiZP/bYBXvzzd+6crxet0fOn1cF0K9+9Wu9N2IwtwUle3ccASX1yMiAzc7etcnJKbt183YSQA7oWgTGltwKGRAVkJz3inNyVKy6l73bDfEcQjwpjICzFD05lNf4+pQKW70HvLKV61LvkhZ9JAfdPlnn76rEg97Y18U0UXkqVXn6IrZUKxX1gKnXa1atlGy/WbeFuQV75uKD9vXnnrL52zetv1KUOAtCcW1rx56+9IJjJ5BshYLdun5L17+ysmEnTp2x/v4hYSdcbxlxZrMpm5moCkKhznrgmXDmCTKA+Q2egAU3vyN3iz1Ejn22ubWtuKHGzI26Yobsp3t67NPProlcIsYgCNNzlj0yn92wHYDu1NvS81H6N3rciyphj81eTU/c0c+KPRpfWX6rzw+Cr7o+g3UtAnjPcSLlGj1UWnBOd7yBa5DQtadop06esrszd9U7we2lqGLzeADmU62WbWxsWLEHxTxCv75eBLXb7WoR7oVqK8gvt2JyK6Ud7IYK3tNhbWXZsMVr1jZtHwty27Wp8X7lNOPjU1boKUuBv9Fq2vL8ovq7bO3syjaq1SpYo8V8qdo+zaDBJUQQQJZ4RWmch5m7suure3UQcx3SR1VfSeB5+/ZdOzR9yNY3NpXfyIIw9VJhgF2oWxexgV0VRBJzltyS6g4ICl7H2mQ9QXyQI7EPRJWT8Jyo5E7nrrDyVd7Acy+WnJZI+jpISuWTIokL1l/ttdp2zXoRYjSa9ti5o/a1MyetXCpac3fXtmv0ZmlYrVmwxbUNK1aqsnoaGRu15ZUV29ihkXqf9ir2VpGiBSefJYpog/md8w7fjBw4coF7YzW+WLl/3kvWoOm8o8qHfn8mVEaxR06ItNgUIaMzG3aWkODlsqobabrNHru8sqYKI+aNxMKNuq1t4CjjzeqF33DuKOKgst0WqO3hNpPEd/9aoiJyuXvdZ57j5Ylp/tqvelTc75T21fd/Z0fgLD5yyadbm4YAdweSQ4HKnx2Ag/Ix7HRorgwgA4DlCQYBUoFNCABl0MAM++opoMMmdbFmNtCHutr9SaOsj42HRUjiQMILuBnJw5LKoN0Ois921UWqBEkjnwMn8r0P65HkMcvmFPYkMNFSY3IoR00gNTd2O954Sw0ixZLTvNoP8A1VBHh5KZuRvoeyKykx1bhIDboBJagC6VXjPg7o3BuvJznjPSE8SARJlKJsmdDMRoPfIAGUTT0Ojrs1EnpPyL1hUY+unw0LP0VPFEn43etRh51MPS9fahh0NjKRT6lRWupJoTK1VClBoNZBG3/PZP8lFYRsZVyFgTqDg5mPc0vqLJIPNe3DVz3ZPakFpMBfAAOIDFck94554hHgXH7Q/aKKinZzKfXicGIGBS0HaEibnrLPCYgKB77d6/R+REUOGgUYc/DA//mKinyhR9MkKfvUGHC7rc4OX1zmPKouiArWDIo5EoBafcdGRgetl3Ww27Bbt2ZsYxXPzD4947BHYYwCGICoaGBpcZ9CwoJ1FPL5ZidA9N9RURHjdGAzDFulRFKEgjjGkWEf6qsqYeSZxDrpgJcdGxq+F0C0EmHA/axqI+5FiQozDAAmI0W6iYqc9MifF7rrbuAvfo61mkBiKpAAsQHMkoVFpYDvcqfBd7yH36sDpgF6R+zkftTXAidwWYJ4dVh+rTGeMb45aIrqqH2P/kFecZK8+PlZrB9fS96rBwDBlUip6fMev+fJoEr5Sx2iojvR6X6+oQwmZsVzDeAxrjWuPYiKbnVt3G+u/uV3YpxiXnBvQfTwPf6t8moAjKRYic8KMPx+REXEfm1DqXeEYgXqvX5KuTvEUhC78XzCUonfDQA9J2Ei7sTrg1DkfYPkiOoTfz6JcBBpwPxzG5YAGWN82kSFgGaPbxz2omorv54AreN7uTI5nmGMaztOpkqJWKd8bt6ngucWBFt3XAwCQ/NeTSw7SuOYQ/F5Pu/9gJMTEO39OM3bWKP5WuLvsedFo2n6B6H09PwDv3EHMskRiJE8G0rIAd7DhkhWMw0UaA5e8bt+8MXesbdtURbzIMYzJyvivuJn9zsgtNdQUmsGUSG1bgugE79nJ/nymHy/w1YeH/z1nV5Hzlz6J2oMGggJnPAN0iOICtYManNsXCq9gyIregcGrd6qe/PQNB8iz+P3o4k86tT4jCAq4tp3N7dsY31DilUpjJMtEyCoxCTNZpuocF9ut36iMoIvrelETOXxB0BE8ZHPTiQ/ACNEBTkh903+Ru7UIytHV+BCPnPwRGWPHzZqbkDnublZa6nC8/NF9/+aA2B+jfH3L6uoyImKTiz6jycqYn7n43lwvvreJKJij0N8xSampqxcrVqTvS6rqBARhB1F6jdVb9G3p1NRwX4c+3iIMXKirb0+0jxXz7ckJORnalSbwL8gKmLfV04QAqn7EBWqd6w3rZkqKrRO+D04OQlhzB4/eVFg/LkHztmJUycF8qFMRnH9ySfXRBQQ/9zCpySyLSwzAG0AI7k2zh4AQZwPuImt7S0HMRvN1IfO90Pe68qVK/bhhx949WQPvun79v3vftN69hvWX963yfFhu3ntmlTapx540HZ3qXgs2NvvfmAffHzThien9F5UKJw8edIqquQoSO3JWpIFxdKSHTt61G7dviXfcua7Kpo4IyXfbDzAR0ZHlZPzM9YNalyNcbFHFq7qZ0HlAr0pAJv2mra1sWrf/vaLdvTIIfv1r39jt2fnbFfVawVZpnLGA6QBAAo7OClxsS3UWsU+ior2okAzvrDfatZqNowqnDNVtdfGJyfto08+tVqjYY2mVxmjHiYeyNM9VSGhhCVfZg/1s0ZBle1Yqjhh3an0ly++rMq8Ap1zAM9NYB2QIsAg1elUn6C8polxyidUvcQZKZ2TwpOcPE/e8FZQnFOPi+gLk/YTSCXsZ7YgfIoF2TzVazs2OTGqpurPPfuMffj+e/bWWx/Z0cPDdv78Obv47DOy5Cnu7dkbv3rDLl/+2H70w+/b/Nyczc6s2dPPPmZ/8zd/byOjQwIjIQaefvJRe/mVV21lY8fmltZkP9NjPfb1S0/Z2dMn1L/i1sycNTnvlPusBfinih+PuVg/nT59xl555ZU2ofXCC5fs2rXrXrEjIYQ3nuWMx5k1Gs/GVkMuSe+R8w+ft/cuv6t+fozpQw89rDF/6623U2Ud88lthSPmnTxxwoaH+215ecEq5ap9+ulVkS3sHcxhztkCuJteVcAZkefOc5RACxsluQh4jwRVlOpk4GdlFiu/p5CTqppFfqQm21yP3q9c0ryJahrOzcQuzsqqIkzCBfZFqjAix1Zen874nLEPHzpsszN31CB9dKhq2+vL9vwzT9oTj3zN7t68alM0C97dtrmZGVvfqdnTly7JihArofHRUVtZWZMV09LSih05ytiMeT6IyILm8Xv7dv36db2Oa8Bqmt4FrGv2ee8F43FH5FmJ/jN9eh2gd7nSqxgv8SUWyBXvF8qZn/v8q7/+P2W/BXEhEggMQramTiAgqCFfAaynFweiOcBnKrXUY6EFvkPO5RjR+rpXQxFjIHZZM1XlO5A/PEdvVEw1G5UjoY4XXgHEUPRqy6Ehel05qcQZJUB+qt8gJbkuxg2rspHhAWE0szPzNjE2JDcCiAAwFqx7pHIfgpRtidAiTwQbGBoeEUh+7cZNzdMTx46ph1BvsWXPPnnB7lz/yKxZs131GHDLZWJJZaDfHjh3VjFwh0bQt2ZtYXHVhoYnbGMDUapZpVq12zN3ZTlFVQT7xp27d0QKAVgTu8CHEMJ6ZQhYgFfKMG+xeAL30XpMwjZiP/k58R+8hThHvCeP5drWNzdVaUGs4H/hBClv895KZqVKr1dnIDDepnraLRNd2OtVbcRykbdxnpZLituJ7kmEtyc8gkpVRKH0axEpWy7ZD77xtPWVTHbUbtG2Z4urG7bXU7Hb88uqzFvd3EqVPGVb3wb76lMzbcg1PTNV84SUTllm2wQh8l/+zEWtkZvmuVl+lib+8HosszTn9lxw8P+w957PkabXleeF996jUN4bVFVXO7K6STZbpERSFEVppInY3Ynd/boRu//UbOyH0Y7GSBoOxWZbstmm2Ka6vPdV8C6BBJCJTGz8znkeAE1JIUrBD8ONBoNRXSgg8833fZ773Hvuuefw3HkGyM51d3fF1OSUCBtIYuIxRfOMz9HR2qp7T+xARYS40YTkHD69a2vKRxUfU42q60uNP6aVVBuixpLu67+mUbHzs/2ztcdvkB6/alT8Y1n7V9/7vb4De+pJ8DA1TgzDxMIk2OrgQKZmvRRdnV0KtnRWCSYEcbMWzEIwi2NDoAG/x6EhvWMMZdAu7er2qO/ColkPBMx6fATMqGDjk1B6XNBBj+8TbB49honhUTaBGUlCJmvlbhWQqkl9cBL91FGlu1rfqJFBOs+a6mDMFGBMLDxki6pKhgn4XDMHMwkLnwPdQILPZq2NsRnFXlgqODlWwUPDw6bQ3d2dCm4EMoJbZ0e3DnOPP5oRpOsRE2ldhT2HLgZ/6FIih9M/MKDkBKYSjBUx3FZIEjwKnVkfJB8cwGJJJYNKddClq2/WuRtBlo8SgALjVc0ij6+LqWLBAbNRU9LO9/g7iRGgOO/J7zpR2WmI7gPGYJj1KqlF3R33gcNn2tiAicDvAa4gjaMr0JrLTSIntz6yPJmR2+uy79Z1qtsvAMyJK/8tuYCdoHUyGJUOP88FOZ80smfTc68NJVgyIN+W/VDBn0DRDJzruhLIqd/bIZOTfQV0v6Tl+mWm/87v6Tp3TCnxOzlxyOzAXBwIbNiStMna0z7NlZMn0DwnibmQUkMiJSt6Juk5eprBbnfSzU8ZgCU7zEYzuJjuT5Jck5xaYlvYqD3Lfhn82XmA6r3zhI0AiTydRROwTsUNr2fA2CA+r63nkR+uM5DEtLfJoQrtdP1ZFzUz4cyY2x6b1LNK0hIZ8GN/wVLh/fP1ZqkAFcMR9sqhySa/DctYwbxgDfEzjABznfXJM8eSPvZj0LNPEhA8M8m0JUBG75diUr4/TqgYI7UMUR575nVIpljbvDbxVTGUmJiepZ53kmRyjEsp3j+YfrVmvYq2JA2Rx9h9D2xOyu+zHvJ+yD8r5lqNJfJ0fakh6XW300LGcgwpiKgYpNGttSLd8O3GkNejtef1uNNay4Rjnz8e2yU+Zokl7XX9rPf51t7PnyPtq7wenaTjEZK0VlMS6T2lVWlQV0CvjTzzJIXf0wUBRQRMLJiwOiO2PDcYYXcczmyvPKmQ7+sW0zmZJsNA9DlnTyc3AnbcxxSDMuCYwUbWPb/H77OvtwDJBF7n9cyZkn00uAZAIO5znmISoJneL08POupbgj4/G4AZ6dZmBj3+SUmeIzP38/2nAenJEdh7NSrKAARozOcGl2OnY07eB25gbDdicyyzPFYyPa1htB4WcHvyV7KxHbE6T3dsNUGSuXQG5AAwskmg9WIdT/Jz9j1LsSl57+SR8xzzuZesDYHw6dnn18kxjr2r/Z5NoNH81VSVtb3JV2BiUYzBaubfuru609pz7MznshmHqeGQgDRdb2r2CMhNfgECa5KPDc8pF7MZqAGMy7HJxI7mrYaU8ietf3sBmc3sZg/PUkCOTFc3knRmjZ4vMRA2MaCQ8zPHc35HUlopzszMzCi2WNu8Tuzg3JDy1K7zB9YC71uA0bbli2XmJYw1vljDnBHcJzUqVKzCYEPLuU3XCYi1slLUtCn3D313AeTIcpKfpnNS058J4FlYmE/nici4aV0A0DTpdchPYcm1tLfH/MyMnr8BfOuvw3ZGcgufKbEeBebSHKaZlvy/FP+Sd0I28U3a6dsNK3ehdq4rg7XbXhPZY8WBK8XS32h46XlBQEnscBXJWZ5T8T0zFrcbhzm+aJ8nMFdnYpLNc3w0U1bnW42lWk2Y8LPD78EN3LrgnsrRQEcKGuqNup853nMN/C75qeKINOyrW9ITee3mz5CBSX4me0WQbwOidXV2C2yHsIT8J+DhJxc+j8NH9stToK21LcZPndL5xrleXCtKNqWupj5a2zs0DQ1ItIguvc5x5EhgU1bleweAi0k1jS62HGcyDPSxsbGYmJgQq3Xvvr1x6+ZNTV6PjAzHxYsXrYtNDrFRinNnj8dL505FeWUhCguzMTo8qGmjjUpN9PQNR9Q2xIcf/DoeT89Ha0efQEBiFb4SNFfYW4D189L0N0BL/HcjvCGmZ2bkC8C1Ia2xvLSs7/X3DSiv4PPgFUHdUtXfYRh3qJ7gZwFulhbmRazaKK3GsaMH4+TJY3H12tV49HQy1jY4Q5qkKQ6wDPuV39dU5SZ63k06+zLTHTY+uT0qHjrfqxvR3tIa9ZIAdvNgYHgkHjx6FCtra9GQmN+SQu3o1J5SrKVpsbqqKRd8A5jSULyrYRqC3NY/Q5ygdtJ0B/VGxTFH3kXIi+B7IFAM8JRYUIqe7m5JeuX9J28L+S6ybk0kMUmtXp/Rubllzzjf2OucKz5nq9Hd3R67d4/G7Mx0nHvh+ehobYmZqWdRWJyP4yeOx9z0RNy9eycuXb4XDbVr8ad/9kN9tj1HjoKyx9XPLkZPd29cu3YjVpYr8dy5k/Ff/+bvo7e3U3Xo6dPj8dz4iXjz7XdjcXktJmbmTXSIuvjG+RfiwP698dbbb0v6aRXMvh5z2MoWwYc9eujgwdi/340K9jJA/CuvnI87d+/qXqwmz0YaIMQQGhUGi5FNseqB7mdTg6Sebt64rpyQAM7feWaXLl3RGeDz2XkV94ffpfHW0oxUEHJHBQH0nC3ce9aTDHtlZB5qIrFOWnmtJL+k3l9tvep99gX3XiQ+NU3JcVxT8rnstbEtpyi/iQSsc4aoboYI2OYzgr3EuUZc20nw4z5w9othnkhBblzUxeDAQNy9dze6Otujt7s9Ht17Fv/2z78VR/aNxcL0RMTGumb3wStWN0pxanxck358NibZbl67HqtrpTh99rlobiUWzatJgcfE1PRslKpIANmzxcoFluaBoc+1dnR2x+r6ms4aZJNI3gCxd+3e4/spljeTQvYYEZkhKTqwUQCIMWqmof/55xflg5OnNNQUbeFsbY3/4//6P+PiJ5/Grz78KB49eaoYRyxKhbviN8+XtZJJKco5kNqRL6hJiar/dZ6Zol9b43ocTABciRjGPZZxt/xtOvVcZ2fJI8xSF7DPmUZ+JMP6unjxxefjwf37YsAvzc3rNbhHPGPiI/evraM9NdYr+szEwCIeEs3UWAghVvW8ejub47uvnY/FqcfR294c83Ozsb665vUI6RNFibqaGBoejp7egegcGI7yRm08uPc4FpdoyGzouXV0d2sahtygrbXDUzJJEp3PrImGbDZfy0RJs3KbFnwp5LPF+UDNu6H8g+dJDLTckA0f8R86eOhQPHr4KHr7+6K5tSXm55fi6cRTEUFoKnP/Weee4GtWHjLQ3++9w7TN2po+H3kWjRzhSso5nQvYo9HqCJD2FAPKJcW3KtiNSA81ceLQvhjfv0sTKeRn9qiMWGfqEdmwmoaYXlyKOtYxzelyWdM+zW3tMfFsQmtYE7COWCKzZkqJ5LZzUfmPTGM7Fm/7pKYfdl2JfDpS5dVN5dusQ02agWFtcIYiG9aiNcIUF0RfJomIrKwd1v8K0mwd7XoWrAPuf3d3j+IMhBpyYq9rY5ZbfhcieUDIQKbOEszgZtuTIjuv9Mv//U8Rl/Jn+qd/M92pHeoQXzUq/rm79dW//97dgV1p9I4kkPCQx+wIrBqHRV8wjQjm8OGizcHNxZaZ9QJ/ShjO2FQI4AK9zMyyMLjjkXKSPhIcEodt8MZoisGmbZmkxYUFG54mgCcb7PCzOsCMvG6B1zuBuFx89fZgksPUQ1ssLC54OqCWA4JOM4e0GQF8cU0culyr5Z5qYp6udxt601UlVgLxE8hF159gqNFtPh8JNSCApjksn8RBioQUAZp7m9mbFHto583PzysZb2puVDCUTwRTEhQpBD0OLA5sjeahikrBX4kWmESwpNSYgUnqoibL4xC/BBjC/AaAppmQwBCbihlUUVG/g3+YSCp6XZlzJw8BGBN0pble7o/ZZ0gzeHTbhXaW1TDzA5NrDh8M/KgCbMxu0FDAkd7YIMpvfmUw/kvFNcCNXsNgK4iDAdCsf2xw08xG69XuBPUd07cZromOkxKxZJ24g7lqAC0xBJPZpYHYLB2ybfZkoMBJosDyHYa2vKsmccTacRFAgudGnUHonYzI1G+z4aRez5eon8kmndv9nHTv/RqZSSq2tSZnfL3ygEjAl4yXBQYY3OA+ZRCRAiED/1uGl8msPTc99D6S+drWk8zAy9Y18iNfApNhdrroZJ1mfUiDcW5ueV8ZpPLIc2K1Jfk0g/4GggT4pcmg3OjiPufGFwVL3mssL5IRFToJnNO+Sd477HWSRPayWDCSJmhQ41CxRw3UtBZ2JFDEBEm7YY4GQAZokcHFtF5yss06IknK4HcGPsUYVuKmSJaY0jsA+gT05YaHmgpJkkBrIa/XfF0JzMyNTT2X5GXA59c0VNKFzyBAXnsAIFwX6yHH3dzg4PrEmk9MboNLvifW9vT9ztfjRkRqHqdEMgOvGUDOez5/tpyjbq379Pm8R9Kzzc1oycE59rBmc0GwM9HV+6c1zs/lNcq15SYmryuJpBQa3PDzXsqAsQtwn01i/qcpBMsQciYwsk1jDPkBxyIXlYC5bohwLRlI5L0F/qTGHq+R1wbnWp7uwKQvywfqNXT+ZMNXA+9IUHjPuKDXvUryF2YMuvgQAA44kM7LvFcA1DNg5Pvvzz4w0B/Pnj3bmk7IzwpAkLXhiZQQ64/YMb/gwtH32MXszuedryHvdb+Vgfr8HInlPT3d0dvbp89DEUtRBevMLHI3m7UEEvhN8cA35bPR2CiGsoDwVKwzlZHXxFZRkOKWiAsCWr2J8jrgWYiRlgNv+jfYoLyGpoJSU5LPzjloSRKwuooMcAFC5mZntVcha6ALrliemuw0dgBHvdbdwMtNsfxzbrq68ch4vgz83F0UuNrb17t1L3gtT1eh092je4E8jWpdmgftJmwQf2XumHI3ziJAQzGlU3OeewogyZ+sKe6/86kNN55FnPBa598BWzF2VHyvVkRMAYzgfpEnoMcO8QNWJyw2rX2aNGlPAihq/6aiS+SUtN/1b/UNmtAzU66qZ0yBTNymYOT68nlAfsJ1sf4gnrCHAJORwjBDFUDKTTb7hsHW7IjJiWmRWgBLZ6amxDilKQELD+CTaVoK/mzky3tzJvA9im5db1pXKcPRPcuNwhyD8xp048+5a9p2zmN3xMzc8M3NTRXJqVmZ92OewMx5UCZdeMKJnM/vo732GxOJWYpVkSRNBgFCW9aV87dW2s1uHjnv8tSxgUmxD+VPwh6sCshrQvs5AVUiFlTdVCslubJ8Xfmskw+HiByecub8xWhW9x/pD33e+ujt7tXn6GA6KDVKR3ftEvgBa7laKsfRw0ccD4kp5D+N9dHR0R0XPv4kJqZn4+DhY3H77n2ttd1jY/HZJ5/Fgf0G++7eux/Pv/iipgtYE2imf/rpZ3Hs+DGBday55194Ia5dvaY1PzQ0HF988YV19yEBbW7EN14+F+0NmzHcD6N2LeZnp6OjuzN6+odjdgYj1fa4eu123Lj/NDp7+3RPl5YK0dvXtwXYz83OixgFO5j90j/QL735/r7eeCavirbo7bVBL2tyZnou+voGtK7Zh909HbG0OC+fFqJad09fNDe1xtJiIfbu2xdLCwtx48b12LdnV+weG4y6us2YnHwWxfVKFEvVKDJRItCLqWiMT/GbqJepOfU2uQAAIABJREFUNc9OOvcQLdi7eQK4djMqZaRxGmKTqS3O47oGGYSPjI3Fzbv3YrW0rokoAECeKZJBgHswwp3HsIcSqzax5AWC6sxyjJY8rmpTJJpqNZEB83hLAUC1ovXxFQ8SoQ6SWY6tnMvyvdiSIDbBgTqLtTs2NmqPRXkMWgZXgFS1ammXCu/vepX13tMFk7om7ty5FSfHT7rx2dIcjx/cjy8ufhHnz78U//Vvfho//ss/jyivi3mNFN/li5diamY59u4Zjr/72zdjYLArlgsrMX56PM6cGpeZdmFlNSamZnSfyYBe+9ar8n9444034+GTZ1Hf1BaBD19drUyMZVJb2Ygjhw7FyMhovPfuewLvyGNfOX8+7j94IB8ES8+Y1EasUh6dmtnZ7QGzdUA7/C5oyBETiKXIqwGw37p1O+WDZuiTE8lXsVLWFBDnZ1UeYDWaDOIsFxt/cUlrlak75aPpbGJaRXVzqv+zhEuWw8lNWzXEAfFFKikLLOX5Mi3R1WXAW7JPem8HV0BcyTOrRjdpBABbU4OYFePlQJ5GQzYFY36mra1FpIPOrh55yehaWxpi9tl0fOv80Xj53HjMTT2VXExhaUUG8y0drXHsxHEB6fjqtLa3x9PHj2NpuRiHjh2N1k7Mo9eisb0jJh49ianpuajQQEHGKJERMGlmrSPWjEqAmqoQQpMv4PrKqjCBkbFdasaS11HF83+Ijjm3FVgKSRCspNb3oVBYUeOVnIRnAJmC85P8AIkrYgjG3j/56c8kHQeIznoBDIewlQlhgL05j+fsoX6yfxDTL0xOGT/h/N6J2IKZqKbYrKac3dOhQ0NDMTk5LX8OTdAKDyIvRt4IM/CWOHxwn2Ii+crq8rJIn9wblDZ41qx11gW5FQQa8hGk55hCUBVcE7G+thKNNZsx1NsRf/DtV+Ljd96MMycOx8zk09hzYE/Mz0yrZiZOriyv6bzXM2hslr8IjcHGdmT4ivFsfk6SRwtzS1Ff1xTVDR18Xmspx+Bcw3tG8Q7Cb32dpKTaO8mbmTqpjwf37moiav/ePclDpE7NYnr7Cwtz2jvsV2TU8j6hVotEkpydn9dn5tkhuUTDKud4rAX2lOp81Z/EUHvN0pQ0egI2YHxABAd5NrI/6qKnqz2KhYXYWKtEW0NtHNk/FvuG+nW9UzOzsbpejhJ5RlNzsAqXWSdNTVFYKUZLW1ssIUm4YeIBUobO/zHtphnlJlSiP6aU5h9iQTnX+af/dH6jZkULeUNTarTgR+M9LnyxBj9Bmu1MEaVpbaaBmNaVNNuC6h5eiwYQ5wwkCf5tBX+bRBpiTzCFqXw7mYLTjCYO8m88L9VXWRv/n/8AKQfMGM6Xf8F54vZ92apjfoM0+lWj4re80V/92O/PHTiaOvE2L3PBrpFLFaJmQsFQESMFPUemBZo5ZKouyhOYk4ENbUwB5ZYT4nAk2VXhlJIPd8r9+p0kFWx25Il2mJp6NNlTDBTj2fBHADqsgQQQZEDS4/gORNtxwX8nKOfmg0bsFJyQ1oAtYrkmgBC+8pQHn0tsAelgwy4yI5sDh4IEEMRM523GPyPPMJb4PdgJHi9d1/ugicfYnjrYiTmXC2mYThT+TvKS9AwFeENjdLS2R0dbW8zPzccc8gkkg+DzmOKKBeROMc+O5IzkBwbuNrht8EpgNEzGNMYskFeltT+npKJ+o/WbJy0y45+foYBkPbBeSPgUkOlYA4ZJL9iAnQttS+O4iHbysv19r5M8wZCBfwM/Zl1use3dx/B0SJJ84L+32KV69GnyY4uxbGNEDpl1MWQS2ysxB/SwMziQ1mZuLJiNnRoOHN9p5DuDbAYg3axTkp+aaxnkyvq5FLKsrYxz5akhDrA8ycMaYF1krxfuWZaO8DMyy5jftalsRui2gY0MvEp3PXkweGLFLFQZp2WQGJZbgzWQ85TPFliiJM5gnZoFyTQ+gx5bE0hit+Tn4+eQmWYyMUtMSzekXADRQBM4BztOky6p+ZYmpHKzk2tmj2nkOgF0YognNr2ZGAaUc7NCAGd+mDtutpg1LS32cYFtl6ZHMuMdwzOukYYqiaK9BNB6bVTTkWugAFoqrERdg3WGtX8SQMP9AHjMoD33zIwKN/bUBBKb3M9QMS1pLxuwcvGthmFqembmXm5I8TwyIJ5le/yYXFBpQiZP2CQZFiXHWaqqznq8WgtpssrFu3WiBb4nhitFOc8a8E2TWcgDweBKzawcc1kf2SCd50sjmWdhOT8X+/rcqfXpMjjL0+xsEP7Dc1ISHC1oPVuzNj/OPNFjsMKTHbxXTtbynyTuWbPae8cNgtzYEWubCbkEgGZZLM4RAxleX4IK04SUfH1SM5Q4lU03HXYstcAaz/Jfme3PucH6gqnN+WL9ZJuy8cF8/TYszQz6tPu0ngH8c5NE75Uma7w/WRfbEz1cM+uR98sTfjqLtecc6mjIf3kyykx93pNiAoAwN1n5TDT1+vr6pBmcwW8DhiT1Bn3E3Kut0dg7b0ShlKeCuDcak85N1fy4Ux/1S7yp1GjTZ6RR0dsTu0ZHdP5qPD2dm1w/jcutJD2ht7mg4J7zTAHHAUaQSIRp7eaQz1bty8S8l7dRkjHhvhEbPWGappdSc8xrcVMxQT4JeS+nM0b7t1pRYQMoDfg2PDgQ3T3dMT01pTO5o7NDAH2WmuB2UFRynVmuUvlGMjfNTcz8Wf0sc6PZUl3sF4gOrDHOYwB6zmfJCzDFUzLDmmfDnhoZGdG6Y1/DOONnYPO5sdAhYDhPm4p1u7ame0l8BwwUwL9BI7cxAFKyX5nZnLVi6vLv3ASYtAALea9x7Waw+1wQkFKNLU1mF9I+P8TeT3HU+QcSAxtq/vT39olduLaOhEVZ+SP3ljXJ/QRsAciwPCemvZ1aq/YimLExctobgPC8Rk93pz7f08dIOHRGZ1dXPHv8RIV+Oyy7InKjyCLUx8TEtKZnt6SQykzjIk+VGxWp6ZwmR3NeZWmGTe3Tnd5TjiHEn6at5rGnCb6c56oZJOlH4rSZ4MSNPBXpSRdPSOYzIjfEtmNVnujyuSQ5VuUWZlY6hXZD1qBgyDOLxqFyaPaj8md/jpwHIROKNjl5Hgzsnv7eWF9BMomGh5ujU1MzYpICxFoiJLGgIe4Is9rU2cP6EEFgeUV7gc+je9bQrHOHv3e0ci2bkvRgall7lhixGXH65CmBi+S2SH80tbVGXV1j/OK992NqdiGOnzwdt+4CONbG2Mho3LxxLY4dPSrw+979B/HKN74Vv/7k19pTI8Mj8fnnNCpOqEkxOzcX586ei6vXrul+0AS7du267qMIEHWb8drXX4q9wz1RXkP2FZPide2TuqaW6OodivJqJd775YcxtbgaNfWNIk+xb1nDfG5iheIMTbCNivYfcjnIsRCPZ2amoqOjLbq7YVEj4bceC/OF6OqymTZru7yBPG29JiYAogAM0bxHVmagfyDOf/1r8X//+38fZ8+eDJYAjSa6SavlaswurogQVcvkSmtbLC0syQOoHjtVEc88pcz1Ab4p4AH+lVZlzt2GtC3nbqns3KK6GUOju+LGnTuxztpJU43yg2gAMPLUhAx/eX3ipyavYR57kiGb/1JbMNnF2mGdso9sLu4pTO4fZw7M2QxaSZYmNc0zUSBPUbDvskQUtRQejK+ePx+tbU2aWOlDsmduzvXNBjXvmhoVS4X56OnpiocP7uvfOtqZ9umILy5+HueeOxM3b16P3fv2xoFDB6SfX62U460334kXXnheXg+9vf1x9tzzik3UjE8eP4lfvv+RJUM2KvHiSy/GqeMn4yc/+WkU10sxM7+oe1zaiPjD774Wo8ND8dbb78b03GLU1iNNbHoY/o6QBWnCjp8alxLCB7/6QOcaDZ1vvfatuHv3bjx9+tRePzwwTbgZRBTJTooFNNtNNCNGnj5zOr64eFFnCXnOc2ef0z794tIlg5tZ1k0TKpBiQk3AjvZOgeDcMyaTMoEiTzjA7ic+ZLlM4hTrhTWQm6t8jwY3eZumUpVfeiow14+udSxJzDMlVopsk7w13ahnyp7n6OlMgbyarDVRjBrFtawn8ERekUkxUjEd0d3THwWa7cjAbBRj+slE/NHrZ+K5U0fi0b1b0dfdE8uF1bh67UYM7R6Ok6dORnFhUb5ONNenpqZjYmo6jp0+pamiudm56BsZjeW5xZibX9L5sby2FtMzs6o1qAt5qPW0KpA4hhyDlKLOSYzTAb/Lce6lF8Su57MyZdBQY4+VtSKqDQU1SWh+rJaKOteIm8hJsy/yxNri0qLi2czcrO4Hi4Im7F/9v3+dYhvEOht3i0CRpkBNNjDxK+9X4ipMdJ4tZ7PymB0guWqMlE+sy+gbyTzqEYzTLQeOjh54MHGQf6ps8owqagoODvbFApMU9fXR1twqKSJY8pwr5bKnG3l/zm5iOE0LMKRGDMHlb4Q0d21U1ouxe3ggvvONl+P9t9+I504ejRtXr8cL33w5Ht++FSMjQzE7NaVnp6kBcqmNSpQqXE9NFGg0tbbHwOhY9A6ORGFpNRbnlmJxvqB8wd6UngahSdLU3BY1NQnEZs1xjtc3RnGtHHNzczE3My0fiPFjR9O9bI4yDdWIWCkUYnnFn0nNd6Sy9BqhhijrgWkR7okk2TfKMT07G/OJ5CtiiUzQnQPvrAPI8TRFTDNYtYyVFETGURytSmpu9+hQfPjL96Ovsz0O7tkVtBip8ianZ6KhuTUKTMZB2KEhgbQfsnvgaxv4HJGDOj+amZ7Vs3VNlvsHv5tGRS4x3Kiwl0ueqNCZlXxu+DfWiDEaPGqMBw0ODWrNZZIi9901H9PGbvYtF5lqQiqvQXGNmEnMVnOVydHUaKQWs//Sv6zpsrMB8ZsV8leNit8fbP2rK/0d3oFDzWaisAkzcKmCfGMjRoaHBULw74zEk0jzNTs7pyQfhpsZnrnoNMMZYJDiTGY9sMeTybZArw0YCuggthnIp6uZJBYMUpJsGPzmtey5YLBXBXDShjP7MUvkaKAwgQtmaG6x5AMdy+YtMDEbaKHlSKd4anper4mxEgVqoVCMkeGBpI1MUmqgc2p6RgUwBQlj3ACWdGA56PmT1zAgnNjuKvbcUdc4XyrMXNh5JJPfIXHiIGWkFVktQFM+DZ+fsemezq7oJNFYXQ+8Oqq1dKvRXqxEDV4erW0qdACVOXB4TQ4FA52WYMmyEorFSgow5/L72+Tb2oUCwPIEhsxK3TAgiciJW14bMj4DUGaUl4kFFZno35oB6zFcvyavL3MtvY51Zv3+O6cotpmkOwHRXGxk0CaDlG2JQaX3Z43V1mnUP0+wULiwXsTo5Rm1WKuR66RoFEMrMRddrPD7BmK4Xie9Zt1wDynUthoViRGrZ5X0tEkss2EkP8fvSQot+bJ4zNFNCA5Onl8GzDNjmokY6UMmJjZ/Sp4iAbYCbZORGQ/GwNU28KtWU2JBuoHmoiGP5bJnAWN5CwHCmA66g6NrlSmixriZJipHM9IACQzObH9PX2SAuKr1ymtwuFPU6L4LbDKDQc2GKkVAyWBCWmMZvITZlHXLAUetO2/5OIG3YspnNjp7C6Z5k+4J15EnZ3hvEkmZ5iVGMPdARmZr67FSXNPn7gdASQxhCrcthn0y5eO+tjXbDJbkBL3niclJj8FK6q0mKmXWr8FOGdOl56MR8tSoyA0aG5q6sOBzUmhlnVd+L4PDOaTnwjuzZzOglZmAkitLLFzHD0Aem5F5zwGY53tq+TZ5D6iplqU0ADLclGlCWkqSV+xLN6j5zLwmshkCIMXYSfI7tbBRLPeivcR+SdMVWeM2dwC1TtJ6zawSGy57ekZAXGJQqqlIvITtk4wQKapgbPHZVVAl2RFio436zJ5RMgiwnyaoOAsAuPKkDbE3N0Uz+JobA+wNmS0mgAjPGIMiBklYa0zCZdkyNRY0mu/mVx6dVnM4yZ/xObgvuYGopD+dozwz4gzGa7wnv5+NCKWtDUsHZg+FOCyxlaLOoDxSzBrPbHqz3w2oY6TKvaBRQFNETNE0peRD04U316+zJUmX5QZZlg7IOreAprzn8MhIPH78WDJMnNPcY57/cqEgORTYg8R7TQUuzKc8woxOTw35LMvnuQElP3uuyM82nxMADDBs1wXwj43u0n2WWSl/pqYAn+3e3buOp3X1ahbyOrADHzx8qO8PDAzGw4ePtHYB6EWGlQEiUhT1KiKnxJjH74CJlEZPgsqo0sAq+RDvqT3JPZXfUJPY9W6+0wRuFFNVUoxMaalJWCOQYPeuEbETnz59Iram9g1yM2Kju4DleUJCyFrCkrxMa4nnKzA/TQ35AHOeYVlG2JGNAh9gKPKPAJ68Lk0H7qMJGf4sAB/cI4gRxGEkdLgfmJ1SrNGQ5N7CQpQUJObZxaKujzifPWMAeEolEzv8fHNzwew0T39sJnNLG3Wzzyj2AaHc6EtNzXx/19fTlIJjEACozrIk06izobIRe8Z2x9DAQMxOT0d5oxQrqyt6LQrMlZXlmJyaisOHDgm8hQXO9CwMRJ4L0maw5bg3anYluSLyrpYWP5O7t+/H/v17Jf309OEDPReaLcjAwQyH/Ujxr6ZTa5u+B/jB/5H1kMZ+E2aZnAt8Ruv5q0GT5KhyoyqTXMhbiClcczaBFciWZMTyuSkAKcV4gwqYZsJET5IfkH0AB2ApJz8nwHpP3ya2YTpocvxUDpblXmnWp2aR4me9vZkAiGhUmIASyjfd4HWuWVyBnEPTCUJINfp6OqOzAwYqZ5EJPgA6k0+eRn19U8BzqNMZbyYse4N75fvLmnduxvnMPdYEW0OjmnzkxIALw/2DMT07LTmTvfv2C+wVuaC4Evt274mBgT5Lu3S2K1fv6OiKN996LyZn5uPEqTNx8/YdAd57do/FnZs34tChQ9o7z55NxNde+UZcuPCxmh3DQ0Nx8eIXYpBT9/B/ZHmuXr2qiSWaW3fu3LEcCmtqsxwvjB+PoZ7W2DXUE8Xl+SgsLcSBUydivVSJ8hoM1rr49adfxPzKetQ1Q3Soqt7gtbL0K8BVzt8BVEZHRuPWzVuSIMEovr2jRfuFfUGuNj01F2NjewQGE077B3tjFgCpthIH9+9Xc+LS5csC9GCzHz16JIrLhWhpbRbAfuvGdcmJAHy3dHbH4sqypFJoVjAlifxsIwzdNInKmdXY3CjyFM+S/Q4YD3i/vLgQjcQ59PepMTAiHt4V127djLVyKUpJnonY1NTYotoGQI5r4/yXQbg8w9wwI35TexGr5DmQGpmOK5DeyHE8Abxt+uuJCvYtOS97nvjHOcS55lrHk5iKoxBR0BSvVOL06ZO6h1qby8vy92DNdXd2RnNjs/bI7MJMDAwOxicXPo7BgT4Z+wIB0pQ4d+5sfPDhr2Jqcjb27B2Jb772jejs7Ym1wqLA0v/w//xVPHu2HH/4vVd0rg3v2h2dfQMx/2wiPv/s87h+/U6cOTMeZ0+Pxxs/e0uA6NPJKRtNB42K74jhj0fFzOyC2N2wlRtbmtWgYW8uLSzGvr17JC915cplN2qLq3H+/Ne1XmWmjWReaho5H+OszDIpPnPZo5wtp06dlB8F94o64eWXX47Jial48PCRanmAbzdPmaKErBOSMtuze4/yb9Ywa5pnSAzBP8XNim2pM/8bOaVBP87G7FnAucL64Ky3KsOmrovPmqc6iRk83+wXRuxRw1skIfzJDOSK5FYibq24QZImTR1zXfORKLEOOTfJg5sa6+PAgUNx/8HDGBocjI7Wxph5dj++/sKJGD+6Px7cuRmDfQOxuFCIjy5cit2Hh+Prr30ripPT0dKAkfla3LxxM1YwSj97Orr7+uWl1NbWEbU1dTE9ORMd7V1x//HjqGFyAfnstTVNMFGv79o1FguLhVgoLEZDml48fPhQ3Lp7J8b27tFaJLcjb1tdYs0jq9SgxuvdB/fjycSzGD9zRq95585dxdiXXno5nj59Fg8ePlAj9PSZM/Hhhx8qFh0/fizOnDkTf//3P5MUmaRsOEYSqSlPatM454ESi8wqAktpVINEDa+ELJic44YY64pnQs5JzGAPwu5n7fb09MX09GwUV9x8dMoDxgAZrl7PgefY2dbhxgyM/olJTWLwvpAvkHoixpFPI3FH/kPOTYMHLGB5pRCtrU2xurAURw/uju9866V492c/i+dOHYxrl27EK9/9dnz2wUdx4vjhuHrlcrzw/LmYnZ2O3n6m2SYkHTg5MxdPn01HbW1jPHlWir37B+LgocMxODgSrT098eTe/Xj89JHWTldvT5Q2NjV1UFhew6FOaxmYf2llTYbN+IIVFhc0CdPd0SoPBSbkWAvEIRoYz54+FcGEzdXX3+dJlbLzLaTRJNfORFhLc7SRwzV6aoL8DQINsoW53iC/JR8TmUU1rDEeOoSadpSUJTluVaod/b3dsXdsOO7euBp7Rkejp6sj2pqa4vGjRzG/WNB1zi0Wo7G1OTb1WrWxmQh4lh8zqYK8TvmyZBdpDBsTzGSqLfaor+ZLUzi5Rv6n//TvEHsgNOSJdOXySeqNQoD119/Xr/yfn4XAAtGK3MLkV3w4PMHkBpV9jhRLICmvFPVzxL12YW8m9RFT2CfFdRvBEwc9XfvPX/m/5ie+mqj419y1r37n9/IO7K1rcCGZ5EqkUb25KYBiaXExJicntelITiiiKFIoCNjcfKkYrlY0hmdQ3uCUO5BOHCQhsLaubjDFAQVhZklnEN1MV1i0dWbppXFQfp9gwfv71ErBKAO0SdaD4TWb1yZGB+NryUSaJJPiXAbfyfjWxmG1CvwkPRzwBHOKcDGc+Z+MQ11kU0Tqc5EIrK5qqoIgZLkCAC3G0xl9NgCYzcCyhjRBj/FuA7B+HU+HmF0gBjHSDg32DRBYV1srRnhPZ7cSN8yTCqurUa2pjdaOtiivWdtVzAUBxEw5wIrdNhsWu0VeEe7M72QZG9g0e1T/kkB3BUBNX3gSRqx/gm+9wYo8sZHlvhh/I7EClJdviHTJLW9hmQIDF2KdcaimEcYteZz0DPPz5VDLzzkX0WppJHBTayMZGWVgJzcR3FSBjYy5mFmmrAqKZoM+mQXtpFSNkLRzLfPhszGzeXgt1q6YQNI6T+Bq8mNQIy6BxTv9A7IUkNkkfgf2DwVX1lfUs2ANIsUhZnO+lvTzAszc2DLYkEcCTUne0vlPWvBbAEjy1MiSGu3J9NQgvw0jMY8SkKopIphy1qTMOvoUCbAebfDljkn2B8kHM0XEtjyEC0WzOX2P8v1VnEgTSexv6bvr/pmJkBnSNoa1VjC6llkaykxbN3a4Zv5dQIyaAJmZQZHpZ8S6Zf/weowti6mailD2ug2VQ8Bqlj7jc7C+KX7WiqtiYZPQeGS+qAQFUAjmLD8H64QkEFBPxoAwjJubNdaavQW2mK7pGfNa2RdGn0drkmdiwFpsFxgtSh4NfEs3NGnfs3ZIfsSmarDZoJiXSDDs0Ck3QzyZzdfXq0jkvii20ChJWs+aiqKpoc9jPVgSPJpVKtoqG4rd0mlFGoD7n6QXYK96KoO1ZF15fh8Gn4u9DcXI3NTSc4ZdK6Mxs6W1ViTf52ZU5tSgIJslaFzY+PPBFDTjFj1US4Jx/ex5rT1NPmAm2mF9dQGtNuU0IOFpCuKXm9xpyiP5NLi55J8FmGctcL9krJoAQYHHYjK5ics9sE8DZsStahQonqapAZ4xzyhP7bjpvj0xZhDSe8uyJ5gX9qrw4+yAdWd2vD+jG1bWlOb6NZ0k+YlOFfA2etseEc6s79w4UNLN/RQrHu193zfOMgpHQAID1CsCayiA0QPm39IBrPMO8MfA+IL2IT5Leu/kaSSSgcb90+RcGgTjvbJ+shpPKohorLlhxv8AR2Fx8tkwBKUgsIyM7ysF2zoGlX29lv9QgeGGHHELzVmuCUNan4U2AsaQUd5FDQ3KV6amJ3fEeq93Xq+1pU3gq6QL1Pi0dIUKuDRBqMlKGpVMNPT363UKK8uJcFAb1XI5MBMdGhqI23fu6FkxPYrOuI4DaQB7bSCtJXYZez/tqXze5MLN02PpDBJLubKl1Y8sj+/lhsgMmGgaJLbWNfGMphhrkO8BIA0ODIpRazapATp+BzBLhJWksawCLJl4Ytg7MUE+WCcQV14uZTf5+UjEPpFPKNDSWYNsUgadeB3p5BeWPS2RGk1bBRexYLOSzNrJ6Fzh5YYNDdE9Y2OatEHygbi2VFjUtBtyNuRyNNAGBoe0ZgGAAF0OHDiggpj7g460gU5yrLqoBWCtItvZHkODA9J/hkHJtMjNm7clezIw2Berq8j/1Wm6DnYmgBnX3T8wGHPzC5aVQEMexqm8Nrj3Zrdn0kieiNO5lvxWiJ2spa3psyz7pElOT1RIdsMvotdjD1sLHGkG7peJL46DeeLS60Va5zRtADkTGz5PT6uhpHVteUj2IvdFuVSaOOLMaoGI4+RMlwnow/nX3NwWhaVF5c00GJGJiajE2OhgDAz1xXoyoSaf51k8efxUwA5rBnZwnqpBPgjghmkVnQ9pOgcAnmcFAJP3OFPGrE9YzY+ePI59+/fHpcu3Y6CPtbgZTbU18eLz52RurKaPjFvro6OrO37692/F3OJyHDl+Kq5ev6ncYNfISFy7eilOHT8utvTk1EycOfd8XLz4eXR3dWgS+vPPP48TJ07E1OR0zMzOxLlz5+Lq1WtqznLmY04sCcukff7D734zWus3Y7O8HD1drZqAWN8oxd5Dx2JlBdmZuvjVrz6Ju48no2dwUI0lQJNdu0Z1FnAveE3ODmnpFyFPjQhURO5pdm467b8WxbZyqRoLC0vR3YU576ZArMWl+SgszsnUemx0JF599Xxcu3pFzTzOuMW5eUludHX3xtEjh+JXv3w/Tp85G/OFQkwtLMj4uaaxQQ04GbxyRm1sRndnl/XN19eUL1oixOcqxCTkXZnAaSLXbW6ViSuAVP8dMNIQAAAgAElEQVTwcNy4fVvTAfVNNDZq1JhSs5rGlZ49sWMbFGLtZ1KG5TlNzNGklGQ53QiX5CRnp2o0y3rw7/w8/y3gGeAsST0hKcOXpaPq1GRoaqDech0kbyERjKr2XoFMkYhlMv/t6oqevt5YLBRidmYq6pQ31MhfgcmUV179elz8/LOYmHgWKyulGB7pjR/88R9pAqx7YCCmnz2La5evxJGjx+K9d38RnZ3dcf6V89ojbT29cf3ypWhqaIq2ppb48ONfR6G4GjNMTkBsKVXiT374vehob4u333k3JqbmNKmzurYhLX3uP41PQNwTx44rh/ns08/SXquo4YCHgrykIBmlvJ4GMmQskbISqMj5Tw7b19cjyTGaEuw91nxfX3+sFdcEsLoG5fn5jOb3GpttYL6wuKTc4NHDx2oEWsqxIrBZ+xP8IeX15A+qLRNJg3yGepx1QcOc/cCfxAOR/RIB0NP9JZG/do3uUl6vRmzKSXNdlglbIhmkCXyReJSTbOiMcPwxiU4EoM1NNV05I/v6IT88lln8QG9nPLxzP/70j1+OI/tG4un9uzE8OCwfjo8+uhj9u3rUFCouLUVzg2v9J48fSzrm8Injkv1Chk0T/6ulKK+Wo7BQEMi7uLwcT54+jQMHDwtPuH/3fhw8eFieInOLC7GyvmYiFaSJtdV46fzLyrXJRXg+tdVaGSAj2VZcK8UMdQ45pBoIy/GLX7wfKyur8b//b/9rfH7xi7jw6eexf8/u+N4Pvhd//df/Wc3Y819/MV566UU1zi588qkaStTlAOOcKSL1lZ1v8IXslTEaT8XlRjoNCs6q3FySqXkifNngGF8LQGFPdzsWzlCxm8gjGTCIC8SRmugj1+EcqrohIpnRlBtRjxFryJ2JHTR1mXiimbJ//4G4futmLBfXo6sLn5LNqNkox9hwX7z+yvPx0XvvxKmjB+LmtRvxwtdfiU8//iTOPDceb/70nXj99ReVTxw+cSRmpiaju7cnFpaWJAX1bGIhpibnRRbhOc4vFOL4yWMxOjYSdc2NUVhZisLKSiwur8ZykbO+NcrrlVhdYQKzXhJJ5Q2oVbWxXFjS/kXuG/lJjnI8LNrbOmKT+q6mRvGb6ThkNdVcTN6nfF72lXIbTOTXilLf0KRLIlBRpyLNSU2RoTQIU1YzSGSHJEOrCZekmtLT2aHGXHFpMZqRgersiIP79sXDh/eVDxEPy0wViBSBPNK6mtNMdojoI0KkayXODoi+LUyXRMQ8UqW19tDcnjvYOYHwL0H5nfOIkEnTtqHB6i/JOxGyNXUW65G4SG7Iv6vWls+JCWFZIYLGRW5eslblW4f5+fKyal7qPepl8iZNMK1azYTnQL2oeKIa15Pvv+uvrxoVv+s7+tXr/Q97Bw61ELRt7ipZFZIEJYAeQeXQ3jJolvZ4kj/a0hGG+eCJB5IninGAVwJGBlFUyMLW4xCF4YiptSSLDABkFl7ufDIanAttkhGSkDxunMEag+sG3vkfBa6Sz2SWnYFmsS0iBKAVlmGnYgJoYJCPkM1Ac7CB+UAQY+rDoGGdEmCzrzejvbMjGJNUSgs7MBktkozxnvwsN4PPRyAxU8CFnrqrYTa7tPdJ1Ci8YAMxLidpCsYfOXDrohbArK0tRgaH9LoTU1PSHqxwKMk4zaAtB5YN5axHjB63GcxZfikZMQJIp/uWtYbNVnczIZtx8bxoNtDaYASXgwwQR9qFFLTJo0Rk/Kx7jsQJzZLUkSZxl6aiTEJ9eKhQ3+FpYDaf30PATQImMvs6M5R9+CTT3tyISmxc7h3sWIoNsZhTgZ8bZlojSYdb48Ek5kpg3VDKbO3sw2Dwcpvhy+9z3Z42sr6zDn9Jnpkhsu3FkjT0TU1IrFnLdWTmMCPMjBLnL3nA0MyjaNvhQZEBquxp4pf88gGep010fxMwK9mbpJ+e9VmZPtF2TQUFyTlAHB9TDTOmCbIsmV7Hk06SHtDoohmheYrDJvaeXOKgZg/Z28ZsKDWLUpKvIk8ycBjbW6BJa1v+YJ6IMgjudQhooymW9L4aBxaDKgHRYro3mf2WQFsbqFmKjBdGm5NXZp0iWcefxeUVxR8bJW9IjxVGE/tQGsSJrS9At64+umDwybSzOZ48eRZ1mESriWjNZ54joLLY5bD86pggqbqRkYx2LZWVJJaySbHTbINIyRSMPynSzECy9AZf2neJ7U8MlryLRni3jU/1OiSnafIkA1b6fRnmUtxRgHlde917MkcNPVj8iZGYGwQq4GGSFYuWGkleNipg6+o0hZGnBTQRxzkhOTCuxdrkknKQtqzNhfkcW2bqSdJop0+BPy9ngWOCmhBIgKA1rmadk8Y8AWOw0TrT/HeOFVs/w5qSRBCNQGSXzKQ3iGq9f00EKj4lcCztWYPVbtbIQFOTcxTVaR8wbVK0Zj1rwZJ+ZnOS+PP0siyBwBYBMDQG3ZzJeydPleR97+fi5rjfOzWh5GnjJJ814qaDJwyy5BT3XnGLvZqeM3/nM0orVc13S0Fxb5lUBMAFnOMcY0wcxrI9EpgMYirDUx0AwjT73Gg2o5/GCA0mkn1r3tarWAaYIqaIjZrM4DW9QhOS55tM8CQvlMBVNWEAMGjo1CO9hAa+jez37tkrUFjNsFpkVDZk3itpRSZ9kvwVsZ8GhcQMU22jaSdyGdiASZ7LjWrHPcA1aWbTGCSmJfPO7YYADVdPhgrU5lxEoxuwjaZ9U6OmK1ij1vp285vGPaaDAN979u6NK1cu6V4hU6NcKp1zPDviPjJGAqH17NwstnFuk8At7TUVPGZM+jxCEseyFbDvdI8rZZnMwhgk32HdKh+JmlgtFrcmJLMWdSdmgzqbPVXH9WDKS+xlooXGoBoKNAtlyr0aE08nNMmA9AznLj8LjMm1kp9YYg9pjjShC8tTUpEuIskNuXcGG5m0SY34NFmTZYIUN4glybRTQGhNTRw5dDBGh4Z1fi0vF9yIrKuJw0ePmmOgRnlt3LlxcysXhWVJA2txcSHu3r0frcgCJa+mBkmfVKKttTFGRkfj0mcX4+jhw2qo3Lh+U55hMKaR58KMmTV29+6TGNs9qM+kQnejKp1mxLRhEmpCWE1ANxE0ZZOMm3NOKIAu+TFZcsX5qMAgmtHEJR29BmvVgNgyuya2YYDOZJnzEL7UcEwyqzpDE8N8e5ovyVBqytLnOc3KXIxLfpXzJk3g8Ry1l2X+ydnkyUhAKsDrGkx4eQ8Zz9aK5c8a7Gxvio6u1mjSNeJ1YHP6+3eZUCH/8bRJvvCV1WLyxuL8b5TWOGuTRiP3F4kTYjgAPo0DYn4boDBgem1d9Pb1xMLcQiAjMtjXH8P9fcrh8yQSDNOmlvZ44+fvRKG4HoeOnogr129Ee2t7jI4MaZrgxLGjesaY2p4990Jcv35VzSv2FpI3p06Nx/T0VMzOzMX4+Om4dv26ZJ8gPSCl49jI+Rdx7uSRGO3riLGhnlhZno9ytRwdPd2xXuKMaI66+pZ4790PorBeiY1NTL/xryPGNqu+IIYCKkmvfm1N/2fKEX8VJPE0UdHeKjNsGZiul2Nudin6evs0/cfCae9okz9FI8B+fW0cOLBX6xwoiTMKvXy8LTar9TE8PCrQ9NiJk9HU2hL3njyKyZlpAeTNbXgRlaOxvik2mESFICHiUehz2ZowS43ZKJcY34UsVmeXjEkBObt6euLOgwfyvqA2Il/RBGUJuULqFJ81mdggUpK00iFvuJ7xZKhzHxolAE6SzE0SUD77Q2cD8Vxmpqm5wX42895x1t/3tWM4XltTjQ0kIauVOHHiePT1oN1PzsBZuaqJHssBVyXBogwtEclojjLAWE8eXVwRcPyzn/xEDObmlgY13b/9B38Q77/3Tnznu69FU3unPDxY22/9/M1YX6/Evv174+qVW/H1V16WVwnx49Gdu3Hnzr2o1tSJjQ1TnHj52re+ocmNjy98EvPzhahpaFYDSM0eDZ76nD148KDOf2SlyHG5NyO7RrXWVNdUaaa6NvV9ZbKs1f5qOg/MtuD6OXdyvSSmcdG5r4lNSYKrBFGimH4f5YQ2gc6AxzxXGprKeZEP1LmteQ5JkwLwCWRXbujcPcc7fjebXruZ7/NG9Ybe37V/nijmetiXns4yyYY4mglS3AhP4nAmLCqeWB0CE2Kmi00+y3kbU9n79++W2gITXEgB1lRLUVkrxr/50Wuxe6Qvph/fj/7e/piamI6r127G/uOH4uChgzE/NRPV9fXo6u2NX390Mao15Tj/7W/qMxYWFqOluTWKhWIsLyzHxjqM7fqYXZiPJhoBNJYrEYXFJe3Rmbk5ebww7aQp3EpZBME/+O633ZCtq9PPIhUFEUOSanUN2sfLq6vKP5Ceeuutd/Rv/+7f/S9x+fKVuHzlagwO9Mf5V16Jd959V+fq8WNH4vT4uHws3nvvl6apI+24im9ns2IWuIz8PmtrRX4g99DkC8oGVaYkjHPwLMjlRERJ3pF8j3heXCkIVCbfhNTA92ZnFyT9wJHnuoF8GClgFCRaYveusXhw/4EIswDPjUnSiPdkn5KP0RQbGBgQniL1j8ZGNXrIdxtolFY3olwsxL5dA/H6qy/HxQsfxP6x4bh26XKc+9o34sKHH8f4qePx1s/fj+/94NW49OkXcfrF8bhx+XKM7hoVCD00MiyPimq1PorL64rb9+49jbZOplzbo6m1MYZ3jUSlpiaaWzujuFEThfmVePJ4MsqlSjS3dcb6xqa8SWpqTSSplCGiMVWGjw+ELk/1co+dF1NfWU2AfJs8wrHQspHEajUmOKsryBCVDLCLDNCqdX3nzu2Yn2O6YmNraimThIgR2vvk/uQb5Y3o7WqPTs6a0nrU12DO3Rv9fX0izd66c1cTi9TcIV+r+liVbK8JQZm8KOJSyc8YebTx8VPyt6FxlnObjOg5PU5YBxIgv/VX8rQkPjRBaGhIpETjdMQfZN8gGHA9ecKLRIx6g/ipiZN0DmUSZSZZg4nhD1OU/B15flO0iARpYgeENpHoEqEoqxZYpeQffmUs7rf+eL/xg181Kv61d+6r3/u9uwO7Nre1GknsMxOa4pLDg0JGZrLZGDiBm9aXrVViwuZm9I4/+T8HmWUHkLFolhmU9fWr0tGDzU0yYSDbRn9MarBxNZUh7dz6JE/TpCRGOnC5eZJASjNHYd7RqDC4Z3O0pP+eAi6BBm1XvmDKUoxnXU35UzDtIT07673DRuAzUJi3t5kBD3uEwp9xWX6fUTHrKFsaSwUfnz0VfgR7GAzyAkgApP02ADVro6u7ywUACUZtnQ4+DlxAez6CQYj1GOzrjb6uHn3+Z5OTMYnuthgJmR1dUXLZ1tqhe+kC1Umb/24TJep3nkFuOLiJ4WkJF8mJAa9mjwE+3dckqZWN0ngtAbEJeBVolj4fiQvJunP4rMGfjXST/E+ausiTGpZI4BB2gpqTSCWeaZojTyRw7W5oJOZO0rDm/mUjJJ6lpxyQdjAYyzqBbcN7ADTrtZM+P2+ZJzuyibtAv8RKF1MuHTN8Vh3gO3TvNdIq5qPZ3FyjwJvMPNdUidcpr5MlOQCd1XRLuueWXPEki5pyMt4ys5xvZz16J+Q7JJ5So8gTCln+xkxlex+Ygca0i581DPpGMUTVMNCEiM2z1JyqVMUGlVli0osGkMrNxPR4t6SPVEzAIGjymDSglX/W0yJml9KEsQYs65vPDthJw5LrETuZfVSy2b2N26yRDdshj+pnuQqac9but5khW3/bF6VOLBMb+Jkdx/5XnKpWYrB/0Ou1Fg3YVU8gkXxgkAr4BiBT3dQ0GdIhsGvRyq6h0KutEcMQ5pz0bEtlFVD8O+uP+0Tzw/rsmSFu8eAMGnLPNREiRl/dFnBnSZ4NNUhpinrSxeAH/0cegvu29XeBUAbBxYpLiZ2A61SceU1uN6FZUyTuWv2sb907A5Se6jIji/vf1kEjxgx9rlnMqAaDpAbOfP25MZavi8aVwG7iCwZ+GWxXw8Xa827Yeg3zP09dOT7JM6jsxhfraGdjRqyfJGXCs1GTCbZOMjJT8ZZM41jTWxJkiVkn1j4xMcVJjYPLO8XG04ptks4qiZUKE92xYVPJLd+XYTZGeDLPxYNhTTrbOnO4KakRms2wdc4l9mcGYoyomjEtH4w0KZEbAZ46M0jI+ub88+SAJ2w84dEgtiHXr/fNTdcUm7IBvd+Ke+x478a0Y4sltPAWCp1VyDcgQ8j3K2KkViSHCLCdfVI0jr+5qQYF6wMgEtCAeJHPOZ9rjVrL3CeujxyCXEAAFE1JNbe2ZZ9yfqHJEk0ZeorG8cWm1sQGNgYyiTbWrlEDkvWeZtAExrAOWEeM3UsKB61g+W2ZfGEZvho1o1ip8regqAJYbki+IKIB5Aa6nxd7g7UKuEbxrDWrqbxaxT8ALJjr7a0t0YP/Q22tTE9/feGCJBdh+Jkxmpn2bkoY2Oe8orHoJqCmpmCOap9acovPxn6UBrmICkyKMAXWomsrlZARMFuO73MP+Mww4mdmrD2tmI80GdNTCcwpV8q6ToxX+frwgw+c26jZZ8AmF5xqwOtMQT6SEXt0volDdfHk2TOx1HnWXKcNKP0Z+Dufle8RL9Wo4LlVq3qWxN8s9eJ1vSG5vvrGTFDYFBDw8gvPxZ7RMTGZAXOXlhZirbQeZ86dU26pR1atxpXLV/SsMSA+efKUABWAs0uXr+j62bPkYQAyTx7dF8tyeGgg7t+5G0MDg3rG16/eiKHhgdi7f088efI4ahswHV1QDodUBsxK7itRCRKMMota+y1Y4s9GoTpb5I22saW3b1lN+6eJAJAaC+xFE0E8fcozsLyf9dYNVDhm8ly4jwBEWYaUz8z9s8zWNgN9Z15iYAByg4EPT9LBbvU1EX+V5yQphJ7urjhy9LAA867uTjUTNIlR3ygfAq1NuJTCFDaiNkqxsVpQ9sXxJNJDa1vcu3k3mhrbYnWtrJyVXACJEK5Nfj7IMjSQFwFElwRukeeSKxBHkC8iLrAvmXp69PihJr8npyYlwUDDZG56Ov78Rz+K6YlJNdueTDyNwaGhaGltj//+xttRWFmLg4ePx/VbdyR5BEP3+rWrcfrUKYFbMMCPHD8ZFz//NEaGBwWGIf00Pj4eU1OTSfrpTNy4cUNrgOd6+/Zt7XtifnNDffzp978d5cJcNNSUo7enPYrF5SBCDQyNRnGNGFQXb7/zfkzMLUZ7F6AJ052LcfDAPhGQeM54CNCs4VmqQdFDg2Je+QyNio5OJF9pDFWiWFyP5aWiZFPk31BCeqI2Cphpw4jv6Y6TsIGnn0VsliUJxH3+4FcfxVJhLbo6e2NtfVP7f2z/3lhYXow79x/EemVDDHBNIHDGAoZLsq4aDfhfJF+T0rr92tirrCn2VXl1LUQXSc2y7t7eeIR0CUQayBNrAN14vxQFVnOukFvxrN0U3vanso/MRgLcnOOqIUxemiYt8vRRlsRDWjZLQZp5j3ybVQCcmzquaI8y+YlZ72ZV8WuwfyA2N91wJifCGBt5KjVkIhTfaOggLwgzX41mQP86ewa+9PKL8eYbP5PqAPF3dHQwXnrp+fjJT/4m/uRPfhjv//L9OHnqVBw4eCCq9Q2xOD2tOPXT//6+GhsHDuyKV7/xasxPz8a9ew8k64T+OzknzYdTJ4/Hndt34tq1G1Gp1qgJV4n6aGpp1DQdAYg6l3uJBBTTkNyrpWXkeLh3VZ3zC4WFrelcPhuTYtSv5Fw0gAH5YXhzb8kDaNQhDUWNhVQauc31a9dNLkr+ktx31gB7/NSpYwLEG5taNDXIfqbOZS3PzMwkso6NmWkucU6z1mmeuOb4R+QjUw1L/GGdgFMIjJVkaL3AaZoPIuCkRpXy5JQLS446+Vbw+4DDfGbyF84l1oabsp6kIb9cW1uJvp6uaG5t39Lvr5aLMfVkIn78w6/FwbHBWF6Yi97evpiZnI6nzyajd3gwRkaG5S1QQ825uRmPHj+JhUIhXnntm1vKB0ytzzydjMWZRU5/gcsTnG0rRU2tQIiampiKgYGhKBRXYmp2Llo77WnDcmRa7Y++/4diqT98+ECyiFGpiX0HDsVKYUV+Gc+mptXoOnL8uJqfeGWsLBfj8JEjeobkVTQkhkeGlV9xlszNzWpik+v+8KMLMcc0DP/IWV9Xr9yBBl2eQunv7dG+QA5OGEQCa1kL5IOZVCOMJ9VNluF0HoynQ3sbMttNMTc7r4kK3ss1i6Wf6uuYbunSpI4nyS01TQ4o+bHk16WzD5JnR6diL029A4cOxc3btzxBzhmySaNiOU4d3R+vvnQ2rn5+IU4c3h/PHj+KPQePxdVLV+LQoQPx3/7mvfj+D16O61euxZnnz6iBceL40bhx42GcPns0lpaWo6WzK+amZnUeCCtaK8a0nmEhjhw/HE+eTkRdQ0u0dfTG8NDuaO0fivmpeUm8NbS2R6DuwVkqImFqzBJb6+pjcbmomoJoBUHH0uUmXhFfyNlpUuX8ylLqyE5jnO76mL+L4LRBY8/T3+QdOl+zfG7ysuMRE5+FJzANUVMb/V2dUSv/p4qaFGqEd7bHnQePoqG5JeZpjnH9Bm00WUpjHU8lGhqSAUv+b6wjckAIaXzR/GN/qsms7/AaOwiZ/8JGBb8un7k0LYd0JF8ifTU0yG+IXMPqBKUAPeQ+cs5zL/g5zoAsCcdaM+GqXo0Jzq8VJNn0eo3K9bmvOp8kg27JTu45E2si+/wLGxU7GxD5luRza+ffv2pU7LwbX/33/6/vwEjFMkW5UM8AkZjPySyYg4QkAKDdTE8Mzaz5z8YkyQBAQU9cMhVZigMWAyz7kg1F+VmYnHnTsdEk15H0XTODlM63mHFJmkO6cYk25hGr1S3mg6SqwAxqHCxs2E1BRzFlAIzPwWFs5nLRgIcKQptucU0UzdKyrlbNRlizzhyvL627OhtXquiW14ZB6wxOtza3OiAmEImqTV1tgBx0uQH9Ga1PRZk6zOvrWzrOgBK6VzLj4b3rZEzX0tgQ+8b2CGS4e+9+zC0ViMQ6hAwKWw4ETcoscUEhSoCGcZHvtcEyg5MGtiwHlUH4DHyoUaWi2QcdzCfuvdiTMicz2OEmTWIHJyBfTFSVsKk3nopxseZ1Zibz8fQszSA0WKlPIwBrQ1IzvMeWma0OXBcYLtIte2FZDwOvAHMCktJnszFyMp1NjYp8fZYmsua9DkgV7h49lX9G4rwa1LGMjhokycAW8DIzQjHqFltdkkYAuZZOyMa5WpNbXhgVJbOwW93gKilJhuXB54dBw2HKPaBZR9KSQb0tDUdf6pZsk0DsJJ0jOaB0WCLnI/mNhiaBSjQd+VmkLLh+j1CblUkhxp+wJ4gDZj/YpHSLLZcMZ9VGEbBqOQpJqkgmqVEHs6alkm+FpbrcDAPEc5KbwHU9UCdDmRGvpkZpXQaD7GFJI8kMFvNjJhDSqG/yxLGkBYx7N9r40mrQf5vd193TE9XyhhJWrot9wbPiPe7evZe+16pnV9ooxfISBpiNYkqQpPA8HiFZUVcXnX29YqPBTtP6U2xoUlHHvWLvZBko/o3kURIdNF5TPBNAlQ200+ewDn9qrqUpCk2hJXkrTaMkL4O8X1nvXIvGn5NhHc0Eyx7AJnTjlriL5JxYqPh1KLbWKWZ6qor4aykhaZxKVqRJjRUWNuzWLAfAiC7xS6woyQWZwZiZIZrGIz6vmVUvJlCD2cIU2Uz25OaDmgRbEk5pgi/5LfAaWwl0Knp4DpnRR5MYoFwgapKsygxi/s7vm13pqRXvQe/fDMSxL/Qk1Ky1f4HYg4AsrEHp57pQzrJHFO28LmzWmeRZxDq1nB9gh5mm7N0Msmd5EzG4FdPcKCFO8plys8hTJMnzSSx3T8fl5oY/k5uZlldzzHGQ4yTwc8js6Cz/R+NI/gx53RG7k1Ep8Uf3upYJGv9pk2z2OOfhepwaHxewkKfKWGOw2S9+/oWYc+g8a5oqszDrYOgOS9ebQuvevXuBZJA9ItwklndP1nyV15Xlq7g3MittZurRHgLa9wIdNqMFXeIN5Mhs0E0jRKPapbKIA4CMAK7sB+INt4mGArq/sFTZO4DZSA8BAADqcy8Bu1mbBuUgTbQIFOd6AP4Ad4g1GiPfrNookvWo9ep9hBQI/giSRWptjQP79qlRAfvywYMHsVJcjvaurjTl4+atGPE1tTLPHB0d9UQZTDQaCUlqRLJ8mg6zhwsF1Oz0rBj/nDXWX4eoAMt90xrusNWTdwt7TDIQm5vyaCAmSdYJGc6Wljhx8kSUyjaXZ3qKnwHsodGSTX0zIcMxibVU2ZJ8QP+Y3ACGPeAT60Cmk6WSchvewx5IjmG5mWUWbBpvSZJr/A6fi8KReEkDgrhaqfLM1wJA9LVXvxa7d43G2sqK9PgXCwt61s+/+FJ092GE6EL8i88uClBnzQEo5ob0p59+rjjAeu9sa5MJ7tzsVOzfMyJJj09+/UmcHT8tkIP/7u7pkgH57NxMsL0x0i4sr8bw8IAkv1gHnA9LyysCFCXFIGbepvJlzmFigaTSFBe8B9SY0xlfp3xUZxwNDjW+soQK69VTK9p/kjYreUpI3h4GKFjLjn/IrroJmI3I81RzltnLcib63SLTvp40o/nZ0uhJqOyHYzJBSU3a86+e19RyjWJ++hwVNxSUG9WQz9L4X4ne7pZorLcEDBNBrd3dsV5YicuXrkdnR09MTc0K9GtD3m59TaC1a4kQsDEDUFVTF1OYi7a06R5jjo7EGfGMtQGwAEA5tzgfu/fsjcmJZ9HZ1h6tDQ0i9iDbxOeQrx6NtZb2eOe992OhsBoHDh+LazduaeoCD4qb167GmdOnNcGBjNf42bNx5fLl6OxojYH+/rh86bLY0QCZsDCPHz8R169di67ubj2Tp0+eJo5JNVqb6uPs8YMxfvRAxEYxisUF3ZvOnu5YKKxF7+CoPCp+8t/fjJW1ShP5l6kAACAASURBVNTI84DmRFlrrrWtXcAOeRz7ClAYuQ+8ZQBxiXPz8zPR1t6qXE77ebM2FhdXJBlIXicgqb0lFubnoq5Sid7ujhgbHYr+XnxraN6uxeFDR2JxaTneeef9qKtrje6egVjDyLYek9iVWOfMJOdTskm64DyBLpKmgsqWtRChrWi5DK6JHKq/tzcW5+aiDoJGmvxr6+iIR0+eaDIVQ1rL+rTGqkBMzjmbiPOs2RPUeJLKrMX3h5xy+xznvCHHIDZn6RKRKcrldH7Z49A5imsPfpbnp8lLJKFa3OThi/fh/ciDiVV4ENCk4LUxiSefdNMjNWxT7sOElky2qU/dtVa+9ad/8sP4m7/9L27s1NGgHooXXjgXb7/18/jRj34Q//mv/0uUyzXxoz//gbyPRvfvj9LKsjxILl68GIsL6/Hd774Wg/198e57v4zCymo8eIy8TKMmhP/yL/48bt+8pcZVfSP3ECa+pZa5/4ozNIXxgYyIhw8e6nOzNg4fPRJPnz2V5yTSf4uFpa1alzOaa1ZtSA2jBlE1evu6Ys+e3XHr9m1NnZDrnEEmbH4x7t6562nP9ZKY8TQslYOWSpomRNYK4BIZLJoxmtDiPKepRyMdAmKlIs8KvjQdL3lF515q2kPagAiUyCsiBiRyHGevAVd7Y8ivMREcNFkiedOycnlqD9WyytU9VcZZxf5STp7W0DY2YGIQ2gKA6N3dvZJYo+nT3d4Uzx49iO9958U4vBfppzuxe/eemJmei4sXr8TR0yd1z1YLS7GyVNDevnT5C51p33z9dTV80PWv36xRQ2F2cia6OnrkOTE1Nxed3V1qirJu8bHA92i9XIpppB2bm3QmLS8txeTURHznj76j+obPBHaBrFBLU5vOqV99dCF68DpgCranN0Z37dYZO/EM2csa4QbS7yfPr0EC240G8hWa0JMTEzE9O6cmi30GTBDidy2Tg1QbzWUIqk2KtZlcZNNnSwqSl3pqBp8+Yl2H60w8HLq73NRGraO+UTEYtc3GRk9a1NSCo1jKD+m5nq5ONVs4D1ZXVqKnu0e5Ks0mzrSOzk41cOxR4By5f3BA/iKcN5z9vT2dsTQzE2dOHIzxI3vj0w/ej9PHD8bEsydxZPx0PHn4UH4XV764JPY/DbmzL70YH779yxgfPxmXLt2OU+OHY3JyJroHemOtVFTTgGYFA6pdXR3x9OnjWFsvxsJ8wf5EZcJnXfT2D8fg2L4oljbjs8vXYrO+Kcr4OG5sqPZwPYzc9rq9r9aZ9DL5Ebk+jKKtWuJUQrWS/1P7R16ZSe3CkuTp3yT5atIPNWGeQjf2YL8P5n2tSkDEj6hjura1Rc22tuYmNWIrlVKsbpRjlekmeVk1CsMg3yLvAQdARo4m1kBfn4i9TP+xVkobxNM61fJAN4sFSxFmHMNS5Sa7ZtWSf3weIX3gL/2RfDtrWdeuYdkTrE9qbCSvMsGWxjVnimqghnopStDskr9ba7vqeMUBmrXVqhrd1NrkKkwnbXnkSA3T5Ez+T5NC5xlT65IYzpiY67OMYW2rYfxjn+O3+94/1dCoqR9+aaf2xm/3al/91Fd34H/gOzAGa0AJgCceYLepMZCAjxwEDXoCuFuKJQNEuYCimN+WuLF0AwwWjYxW3NXN0lIKrqn5YeaMQSQOOA4aRl0BC3IQzlI8hATe28ZpbkzwVa3BSDqxXzerUVwxC6i+3kkOiRGJCq8PIIAeLAGdQxRDMAKaDa9txuyxcRf9Au0AkxcLPvia0IxFr5iiEmDZkkCejIBN5CISthhAUma/8jl5/wya8focGBxKXDsgYU7Ka+t8aNPB7u7oiP6e3gC2mZmbjyeTU7EJYJAMwsRY0eQGB5yTeY/wMn6J7r0TMiVcaaQud5sNgBo0yz+jBkzSj+fQEoAh1pN9Hwyeeix764CU7Jb/znvmsW1AyswOBVThOVgKxx1ujS8mUNnSG4jPmGktRmE6nC1H8uUmRwa3thsNWW9++zDI5sECVNNosCUoKLYM/PE+SogTI9rM0W229xYbWQybpGuf9oabeXX2dkiGSh5V96QEr2lJNTMWxW7VWKx1G920q1Gxb6jRkxNbJqJpakWjr6lhlBnoZpd7jYn9IJMo5EBSgy+Ze/P9rNkJ4MNzJhlVkSOzTzPkuR7uPazJLEFj7XrKXstd5UNXzSCB9IDHNK+YsmHMkz1uwFsA8A6ZIz6r5Cq0zyyZI5+MdF/FFBXDk6TZDAbpw6dJKdbzorSwvTfd4GC9Y7JmvW5Yl0gnwMqhGAeQ5L1gGpO8KQ6QoAA+i21TVPHKMxCo1ETD1hMzFKhNtQ0xOjwizds1mKOwvBKzFdCSz0TCDZuJsVH2zezcnBK2rWmDxNTnbqhgagFocVGdmWiSw5Nes9eY5ORgZNRaPsfPeFNsVti5md281czlWSePi9xUyABV3rdiX5Vh9Frij+/TENz6UvMBZqybS4CMXG/2BnJcM7M7Twhsg/BmUuZ4nfe22OkJ7BeQLT8OzIsZ91/TnlRjjgbhBqPM9ZnHvh37txpbyG3Bxl7WdByyCgJQaJAvL281JTzpl2JRYiRLFiexPxWfMBHXPWbCLMlsWYU7SZHBSOyQnFyOi5wPeF+4cVnRdXgdezKBgG/TuBol+8QZPmv279CERWpEZ6A+TxPCKNI0WgI1KTaR8JCer+R7DOSxN9TUknyQ40uWrJO/EY0m+US5MSNJIp29BlA1CZZkmuTZotE79zp41gBvZni7iQ1jjvXNPeB9NYGR5GEA7llrnJG5uWEPqmZNV8KoYv2iYYzhtiQbUiPT7+lzhNgm9iPPH38DznflBnXaq1yXfYfA4yBB4LlSwMVkK+bkJiXPQnIJUSPm8cLCrIoqinwKSEyQs3wH0lU6wzWRwmRM0QbzsLmSFISKJSRHJOvmHIbGpHx7UoOioZamAobJluaSF1K5HL2dnXHwwIHo6+2Ozy9e1O8Mj47E4tJCYota83kJM9q6ejdBqvbS4HnksXP2NXuX9UahBMDh5+tpDkyOIYqYhe/GIsUizQnuB41jwF3AtydPnpg5yjRQbU0y4W6JSlRiYRGZkhblawIdITrQ9E4TKAB5alLKDL4lFhbdoGBNI3nE+fAEs+QkTcZ1AhLrnKqpTU2lJMdSNeuf1xTpIcntAa7x2pyZrC/iTGt7q8AdGJWltXK8/tqrsXvXrlhbKcTjR49jgYmK9fU4ffZcdHX1bjV0r16+qj3MZ0Y+jKK5tb09Pv7o4y29cwx/a9Glr5ZioLcjThw/Fp/8+vM4tH9PdLR1xoULn8XAYG/0DfSqqdXS2hEzM3PxbGI6hkcGtV77B4djenZGrMkapkfqMai1PJgaIjm/Tb4i6B7neKTcAbBIEhg01pD0tOdO/uJ+OwYZ0MvNSMfoNjGdHz58mF4HMMBNagplF9pmtxLd+J6IPSnGs1a6erq1RiSJWDLJIsdxHjb5GU0B2KVInmJoSgFuia9qdHexz+bU/JSUaX3E7rH+6O5AUtJ5Ps3M5pa2uHPrXpRLNGGZCAaALgs4YnLTKo7e08srPhsWFpYlMcZnBZhhupGmDO/Ff9++c9vADPcMQkSFnDniG19/WVriPs+RpEOGojne/eUHsbSyHvsPH4nrN25Ha0trDA8Nxs3r1+L0yRMCVGbnFyWBdPXqFclCkZ/cvHlTckBPn04opu/atSuuX78eg4M2cMWcmH1fW881bMT3vn0+Whuq0dkOSGSz8faenmhqbovFAp+tIX75i49iZmk1Orp7FNdhgQM+Ih3Je+AFw74ALGNvcq3EL543xq59/b0Cf3jWAGRIAA30D6rZSMYG6F6GULW+GkN9vXFg/1g8enA3Rof6o621WTGjrr4pPvr4s9isQWaEptJGNDQ3xdJKIUqwcJO5tc7p+gbJPm1uVFK8q41SpWQ/g01LGvL53QjYCOJiO89GOuUb0dXdE/ceMB2QjVtrApIPuRp/8uyR1SCeaMpasd7eAVv1RppAJMYIDE0TzJYdxbvFRtA6j31i6N7y9yz3Qe6ja5WErfeTACVNspOjbAiMA+RnnYnEsWGVAKY/BMapoU6NiXyppRZbAOc4+zc24kc//H783d/9bZSRcSlXYmh0IL720ovxzttvxY//7E/jP/3H/xQbG5vx3T96PS5cuBD79++Pk6dOao/PLizEvdu35VfSWNcc7773C/neYN5brXq683/+n/6NPJo+vvBpTM/Mq4GKhFipYiNYkclq6+O5M6cF4NJoy/XmCy+9EF9cuqI1gpa96j3Ja9Is8yQzz9qeIM7V+f/Y2K64fuOWmhfE9BPHT4pB/+zpxJbEc55i0ERCTUg2zYPidWrwZfkfTZEnCUjqC54DMY5cgzirBjNm2llSlgZMyZMd2TjdQJ9Nc0UUYf8pd7YSArExT2IrDiZ1h+xd4nM6+XyliWFyNZ4t9T7PVg2TUima5flUo/3+8NGTGOzvj9bm2ph6/Cz+4sffjN1DPTHx6J4m8R4+eBxfXL4dJ8+djGOnx2P+ydOoJc9pqI8b16+pVhx/7qzkiGcmpmN0eFSNhbWVNdU95epGTEzPxMz8vOOCdPUj/viPfxiffH4xWjCtrquVT1dXR0cMDPXHrrFRNeshhIwMD0dtFSylEktLKzGzsBQNrW3yqsBLgPuN1w2fnUnDBw8eyuAbHAPpw2vXrmqdHzt6WMR28gbkfa5euy7pJ4By9qxzy4qaquwBzgjOaaZ6FJMSqZPJ8jw9WVha3iKoqCnb2qpGhSeTi9HR2R5Njc0y0+Y8oKkhae46zhqamLXR0dYunyomdPhv6gieEa/F6xAL2M9cFzLkqvvwzKFew+8Ur1XOZSZzF+bjhTMn4sXTB+OLCx/Gwd3D8eDe3TjztRfi5pUbsW//7rhz+24cPnYs7t24HUePHotff/xJHD92PC5fvhHPnR2PO3cfRt+ugZiYfqwp+hYaP/V1MTTQr+b50GC/1v5mtTYWl4ox+Ww2NusbY7m0GQsr6zGzuB7r5N95yisVzUymcK9dT/g8V05fbzN6kzztpcq+4z6JPJwYjcQizkRNpzcgI9qomqmnt1fNJ5quGY9ir/Kz3D9qsYrZpvL+qKtsRn97S7QS99bX1YzG/0IufTwfpDvxQVxZje5ueyQtLhV0TnMOcH3EA03PbhJviSvGlXi+5KKqZ3LXRcnHztZEupjfCkPd9ubjNrDHmUpS4zbVPTSGWZuWyjJOQ6PO0k80LkuKKa7pTC4mv+SsISfGo4K9SfzhPFSzgClu6uJSWTUEeQ3PRh6VwkFSA0VT9I6fv4uvrxoVv4u7+NVr/F7cgUGKQ4Go6EZuKOBnn4fMnFfhI7CHUXYzrgyAW4N225A51GAgaJLoyDyRkXfJ0Bicy1JJBE6AGPSO+aIwxeCJAI1JH7rUW1rt6vhauocgYGNTF1QykN4oxczcjIynpQUunWoOa8u/AMzKJDsxdRWA1N10gKFrT+JK4Wx9cpokqaub2PEEOIBOCnxAAwqknACRGFJICHxNfgYCZcSa9CFK0FITRixfg7Bir9Qwxt6qA5efhWVGMIet01i7GQcP7I7eji4lkRh1zReWpfMKVUeyChiNra4JkLJshHU5ud/5AEgKPD7kOIikJ+9OPPdEzKMEQgp0SoahGHDZ6Mz3mYPHHWNLE2gSJrFUNC2RDlJpLGfz4yQBpaaBphbsJ5InKAzWbRvdcWEUwHr2SR4lN1P4bPl9UjXtz5BMecUwrjoJ5h7LoJwiP40SWuc7N1oMoloTficwkKZBEttzqwueTk8dqJKK4X2t65qBKwF8SX6JQzI3YlQcyVzchqowxMyiBzR2scDzRfqK5FTmyRze8mXw9Wk6hsN3B4iRTagzw4h9RiIucChNzAA8AUJIGkma2k1a44AOYoDLgyNp9yao1vseNnyDEg49f9geMNtq0aFUR8XAagL67IHg+yhTbFM6lBAwvUKTRAlsuaR7wF6RsSPrH1A8sQ8osMTcSYxyg85bxHHFqkJhydcVoQkVGykyDtsYfQP9ik+w02amJ8UOLq2vqmlK/IIdzng8bB0AprUiIE2rkhUAR02LNTVHfU2tpio21ssqErVnmxulUU7h1traHosLyUQND52kez83OyvjbS6aIhWwnvViHXy0dtv0XIkNPBuKgswO2wannHBp2it5G1A0c5/QBqZIUBnOXkTiQL48DWq2AM6JVZ0aS7lQzyyn7AXAOs0AYQp1bgymUWDAZsyBBXRLKogmghspWXvT+93NSz6D5PKQ0+KaNWFgrXpPTWXJIQQhbNKYR36JS2ZlmTXcwLQDzT6ABumeMgHk2OzmpVn4NIjwDcmSOGryAdg31kdZkgOAFt5HfNknh32U5FTotxGXZGKevGmS14P0YLXXvPgongkflshaE2AwMDQg5tDU5JSKIwBHMaLTXge4kb+S2O02KyaZ5QzJTQuxmTYopizpIom+NN3BexNziQvo6tPM4XKs0GIzeZngJn8QTWjQ0Orq1FmDNAfXjnGdmdqe4iKG8J6c06wP3ZPsGZGSb02WlEvR3z8otiPTOKwBCsDe3m6bfKe4DYiAXi/68YCDjFVb5xW5npW4eetW8iKwX4iBWjeE1UBKyTtxStNrVeTzNrXPeMawrHXtafLNLGIXHwCF0vqHFb5qdpT8YtSEQG5oLZBX0JQCurKKfw1aT+wnscMBxqVfvKz1muX5uNGczewTNL8582GNLhfwe0hge5FCqxo19fYiwKcLcA6W7R+8/u1YKxZjYmoynk0+EyCryS35CPnszJ43MjfdMg12E59JHkgRWRKJPdUKi7i4qoKxsa5BrE209NHJp5EGK5x1CCiA5Cb5F9IkhzHmrFbi4aOHKlghXACacM709/dFV2+3JTDxL5Lkmc9kAIRdu8bcIE2TYUjt8AyQR2P6wc3+BslFSPc4eU8ARggATCbJxCBiHvkTRA7WIIEMljiyI5yBmERKojFJj6GDr31ETlGO+P73X499Y2Oxtrwcl69ciYWlRRlaP/f8C1rD7HW09y989JHOCkCZc+eeF0MOje6PPkLuZln7mGnVSnktqhtrceLowRge7ItPPrwgE1QOubfeeDd6+7rj0NFDmgzq7u0XqHP1xv04O35EUkXsN5pJgEuswaXlYjQ0NqtZQROOWJd9qKSxX1cXszMzykf5Yn3t27dXTGryS6Ytac7Q7CfG6zxn6pkzLsk68Hus5wzK8tn6+vu1niQ/hgwDnk0wWJOZ9Fa+TH6qCUsaWLAEm2JpaVGeJpq+0USnYxXPrby2rj1z5PAhsWwbm23QCaAOPwVwgvUkOc4KtUDE7t390dtF4w0w1P5eAJaAPJ3dA3H/7uM4dPiIpGhUE9TVyB8Hti7SHDC9a2sbYmJywjKjymXczCa+cM3ImdGwXE97F9BqdbkQXW2dcWjfXvkOKOY31EZnN2bzdfHzt9+LldVS7D14JG7cuK21Bmv95o3rMX7yhGIa0ixHjp2My5cuxdiuYcWmW7duSfqJySiuZd++fWLYcs95fnfv3U2EiNVob26I8y+ejQNjg5LAKi7NRX0TBI1KNLS0R0tHb1Sq9fGTv/1prJQxHYY40Sjw6NBh9ijsYUvvMF3BvkC6hHwHEgT5y+TUs+jt6dI0qUgWxbVYXS1HR3unmeVpIhvJmvWV5dg1PBh7d49K7qRULOjeICHU3t0TP/lvb8RmLV4wjTJ8lcwIDFPkP2Gm17hhzGTECsQPCC0ydV5XbsO1bpYh4LS6EQ0wRlMDH5pEPMgkoPuPHnhiorbekpcQSpiA11R8XZQk+Wl2KkxvAB5iM+vCE+yc3847HRP9/Tzdrn0hGSc3dzMpjJqG6Q1ibCZUce7p2lN9R7NLBCZJsZaiGw+mNHlIzJYuPE0NpCIlJ8uUNT4yluCk2dfd3qZmxfe/95148403NMHOeTc8PBjPnzsXb77xZvzFX/44/uo//MfYqNTEj//s+/Hzn/9c3iK79+5WPnxyfNy1ZbXy/7H33s+R3+ed54NGN4DuRs4ZkzABkzgcDjMpkVQiJdkru1aWvV5v1dXeD/df3e7V2bte2T6XZdmSaFGiGIacxMkRYZBzaKADOl693s/nC4593iu56n7RFWGrODMAur/9/X7C83k/72DzM3N2/cYtq9ZhLZdXQ243U7Af/dEf2H4+a7/5zWcKf6eBnyuigPfxTiYT68fzF86rvn306OHB2ffM2TO2tLSsdZO9DACUfYcvGvKeL+V1ltRW1FcV8pWag20UloSc+11F+mxj3esSrzlQUrHWra1vqrbByox1n6+IJOhkEd/HuU+ew0ajvCzXAuUNyCrYw7ddJcOYR7TmalrO7qzBatDpWQbSoWplr60j3IFnrxBqMu6CW4PUA9m9gywT9hnl9kll7G4FHW1k2XQrOHh+ftk629usVs6blQr2B7/3NRvqbbeFmSkb6Om1paVVe/Bw0vrHRuzs+XOW3921dEe7lBWzU1PWmGqyoeER7VWVYlnKsrW5BZ2RIB3uQUqpj9ni0rLqaWx6Z2dm7ey5c7a8smYLy+vW1depxkCHVKTbNn7iiOaj8pJQhVZjls0WbGNzx0qorbJ5BR0PDA3Y8sqKXb12y5oaE/aHf/CH9uFvPlJI+vj4Mbv4wkX7u7/7qdacd955w/LZnGovruuDX/9GzSDWAxH0wvmMNZj5zR62vuF2XrLVzeW0JkTWmI7HOKmSsROdWauVksgW4EBR1mBmGzY7+48TL2OxqpUqjLealJ7UEJzROONSI5KbxWugsoAcwfmIugTiBWdFzi2Dw8M2OTWl2kTKj2rZ4tWyXTx3yi6cPmIPb123Q8N9tr44b4dPHbd7tx/YoUODdu/uAzt//rytLK3a2OGj9vDeAxsdGbObN+7Yy6++JJVg7+EBe/TkjnW2d1l5n3NjXA2exblF6+vv0Np+5PgJy0J2TbbYU4Lls0Wbnl+xbNGsUt9gFm8UGc4tkN1BgHmZak5bc2urGvrY8bKPc9ZwnA1yKmA56pMGy+c8G5Y1k/NiLzZo29uqa2l8YiM3NjqqfYyxTR3JV2QVrJodUD1WE2ZCoyKuRkXaOtMt2jc4W23t7ahRQXOUa8bCz9vC4ESA/+7exLrIeiCCWWbXyRNyPqExgZIN6z9qdDALt4Q9wHfUrPi3NCn4JFGYNlbGnAHqrLenV04vnH9Q4GxvbmmusA4IW8CmLp/TnOfeqYkdSJaRy4w7vbjyFGu2nd2scA9+R5aeNHgDIQPMkXpQ+E5wHeEM92wj5n/WYPi3AsZfNSr+rXfsq5//nb0DPfuEFHm4lFikoWHBfyObFIoWJp4zaN2Tlomr8B7JW2PuOSvWN5ukb/xsZnyJma3XxS/ZPd9gc8AmZNEqlWvW19MpD2c2O4KGOHyxgHZ2dKppweKhBUNy6MKXtjP7BJm6pz62BSryBMYTHoTELWttbc1aRXk9gA0VCRUPZ2MRl4IghP7yeWBltLY2B0Z2UhsrUjkV7E3uU4zMn0KU//G7nV2dbs0QfC4lO8ODHuZwyDygQIruLxsO3sIUlLB9VpZXtDC3cQBJYD+Sk6Kiq7PNeju7dIjnQLKysWllVVnetCHEG89C+UDK79rBbZkpBQkd4IuD6N5B1jMJCoKImSuGHEyoRELFAK8BIx2QMAJSHUjzQFEAN7dXcu9zWW7pUOHsf3+bZwOyHZB61ks/AtvkJ6+gbZfRMY742ag5FlkbRZ8hAtLFJhZ47+yOyFLFVTE03wBDYTm6WidiECt8PIDH2lxLLgEXcAoAGJjRnlni9zFijOvwo0A3t5eJNiP/3C4VxPLEVT/uK80XIBHXSRgiTQLmD+NDAG7o2qPy0KG87MGskicLeINx6yHFCqKjc88hMihNXAESC36IdWKlalPNu0UKBRvXxxymsONasOlQY5DDropLxrF3/PVaZQd9+TyACJVyUQAthxTAY66HUGXGCAce7nd0/zmEMo8opDhQMFbETLM66+7pDP9GHoKz8P0g3hLGC3YDzqBiTaHIg+nN53aAtSw/asIZ5f/K2AnBhDAcmFORZy3BkQCHqCZgf3V0tuuZ8HkonuYXFlXc84wA5SleKrWyAL42MhpyBbt08aL8gEvYcmFxR8gza2ZQj7B+AZ4AygLSy4s/ldIY4j4wPj18+ktwnfHN/WL8RyxADlw8YOYehw8AGw6HfO1sZ/TcsK/Bcoh51Qq4l8l4SG8LNhdFgYfYP+zsbB0031DIqdkW5Kv4hkaWCADZ5OJwvxlDKHtcIWbW19dvS8tLDvxL3cRM8aaiBqKAqYpnXQgYcBVXFG6o8a01Cq/xnF6XdZx5p3HUQG4Kdg9ujcca49kXHiIt/2ACveVt74Us4wmrDuYoz3ppdTmwV+IeFimbIELzsFzxAFaeDc0E2F4eKOmqiWgVZB/ii6aEmqtqgiTc/imNVZVbeMHModmmpocaNDEBdHgx93R1uDIqvy9QVbJ4LBJgSwfmOMAw89wZX8wP5O/+bDw/wRt5jEsYyt6A4O/YG9Fk9GwgLH4ohGH58G/sM6z1HAyjDBNXvpGLkrDdDNZdPsX5/Dw6mgeA9N58LGoOMNdogGs9gk0bwtSR0UeqRJoXvuZVtK8RnOsFf+xALce1uuTZgxClNMNOkcMWqiqaaiEfA6aY1AsKKvWgaJ4B45psKP7s10mOVMGS6WYdgj3A2bMoUEsJmA3qQAA9ByHqbWt7U4cr5j3Pb2BwQPeKOTc3O6u5ys+73UWdrW+scj52G7fARhdrSgcwlIb1YpwxNyE/CEjM7IgVxnhvSnm+ShWQfb9kP/h3v28L83N2/8E9+eV39vba+samZffyB0oj1gieCc0RXp/7Tj3AewiUkR2CN8z42SZ9Zg5OADKu1mNMoMBhXqkhy7NvAOgzSzcl5VPe1dXhzOvtLa11ChBshLUH27lNzQqAUGomACWAExofzEWY2rC5XR3k6jP215BfcwAAIABJREFUCcBz2SHWqmpg0SBlHjOWZL3HMwr2oYw/vq+MCmT12GIBJhXylk41y2qQ+oh1get1+yNveHNorhqB10lrb222rrZ2rSl4cucLRSMsOa0Q4pyHSeOh3dhkx+XBXbF0kmwT32sIDpVFBKQUrAvrzQrZjI0fGbajh0bs+udX7NSpU9bW3Gr3HzzS/D1+CqugBzi7aI1EOXLk6GGFRLOHEnC6tLJmEDtQAzM6aWgz5vncAKSsowp4DJYlrKc0CmD/0jgBeIII4IdnZw7zAFnPAT8Z01j/iNUuEgUgTdJZqbK9YH92lZMIK6H+w4ueeQiTNGqUUDuotopCY7lewlbxtUfRsBfGs5oYGWtrbrZz589Kpbi2sSqmtOfdYANRc+WZQtdp1jZYT1fKEo1YwpJVB8EnYfVNSbv26TVra++2jGyKumx1Y11WJdu7OwKtqXtoUvCsADjxs8byiHpkZuapHTt21Jm8pYoNDvTLAxuwnmY/Y6qns8Pmp5/aD37v92x7Y133m+tv7WiTouLDjz6xQrFqo0eO2sNHk3rtnq5Om3s6Y6dOnRA7HDYoDNrbt25rTjD3Hj2ZtJPHx/UcmYMjIyNSidGoYD2XYqyGuqTZYrWSvXhhwqqFPZs4fkjNm71sxnoHhxScWqoA8pt9dvm6lesSlpcliLM3Wfup61lreNasWTs7mdAw7hHY293dbSsrS9bR0SqFJXsG4bP7BUJCsRXN2242Y2Ojw5bJbCmn4vixI9aJuqlUsK72NttcX1Xj8fTZc/bx5c8t0ZiySl297eX3vUlJw5t1EnISNSiWnai0CTAmb2gvozkX2W7ShZJnPSG/DQ3ONKV+ZR2KxfWsNrd3bG1jzVnuZVfweWJWndWjLqaRo2B6V5rKglVWh46AicktFrezi6kHWCMiZR9rDnuTyEGynAm+51IiuYXfAYGJjCFUnagCUa6iIoDUsF/QHECtwBmSTC7qMlli0iABZKX+D44A1EOoLyDI5ciJaWwUweXb33zL3n//F5aE2JLP29DIoJ05dcZ++Ytf2r//4Q/s//qbv7VCoWI/+Pfft5/+5Cd29Pgxzemb129ZX1+XnX/unI2fPWt3P79mW9sZa0y5jQ/Eje6ubjsxftRuf3ErWNmQkZfQuhNrSNh+aV/ndtZmiANcLPMcRSHnRPaTjs4ut35tTIjMIEUfQF3VrZ8gRbnay7Q+AbRRJ1CXsu9wHwnm5by9AbtYeyr1J2pfbFjdsvHQ2CHNp77efuVAiWAQ9m3GAeArpALmL7UIKkdsbngPajy3knaVjqtfXOnJ+dyfL2SeBu1X5NdwRuA6NY9kkVknHEENEZod6ZSTtHYyXjMV8tpHeA0RzgKwGNnfRW4PbL/Yp7EXuIK2aPFa2TIbm/a//ucfWGNdyZZnp+zQ6CFbX9mwuYUlO3TihIDl7Y0N62hpEWB+9/5d1Umvvfmm7hdB81gZ5TJkgNKM2pPPP8ptysz5+QW3QMyxl7RrPUTxlC3kbWd31zraO+34iWPW29+teoLxR0B3pcQcpT6LWRu5PukWW1xd0Zy9e/+effbZDUslG+yPfvgj++DXv7LHT2aUYUNuys9+9nON+W+887bOdlzn0aPj9rc/+XvNFxpL1Is8ZP7OveDBDA4OuH1XzPNGZIGrxnxcLh08S+pGP3szb7zhqRqijj2rXgQbcBaBvSXP5fPsQeBzGpRmbc0tUtNhl4Xqya16PNeQ2ob7SAN6a2dbFlBqpFUq1tXVY9OzMxpLsiEvF6y2n7MLZ07YibFBe3zvCxs/MmrlvYw1t7dIOcO6dfXqDbtw4bxNTXKPUNo9tNMTp+zRwyc28fwFu3f9C+s/NGA3bt6wkaExy+75mbOtpc0Wl1C4tNrVq7fs1TdfsJknU/bcCxft7p2HNnT4hE3OLdrj6UWr1jdaU3O7zS8tKZScJrUUMx0dqkWFaUHqCXZWNGRwBvF8s4qIKE7EdccA5jbneqoG5hg/09PTbTM0Kg6N2dLiktZTVzg5ZufZfCXlMB40KmpmCfL5kimLYQHHvk/20X7OMtmsAZtQa9HIUp0REcXibqXkGYqoo11d4OQUVyPL6ryhSTU4cz9qVPia/6xxkZ81f7uvKBeTs4/X7f39A6Gp6nZxi3PzwkGiLB7PoClo7EXYjkK3q6aambHN32UHzZkdJU5wA4hcHZijzekWPQecTtTMpuEtrJSGhavldWYOlsSOm/1bPtv/8w48+/v/rBHylfXTbzdcvvqp3507MCireN885NsJENgCi9rBZzFsxWwBxPE/y9IiSDcjpkMElLmEyr2uxTQJh9vIa1ugrcKb3baC4uL555+XBJZr4OfoDEfqB8lJFTLkLGU2OAGg+KErVA0WNCxZNrayijEWdAp6PDEj+XCkqODaOVRTDAAK4GvtxbCDh1zbgedig3tlS86FLB42CAAcnyuEmPI5dN0BzBNLNMiV2WAAEPgenVc2EMKXOMxF/pssMAATFEwAarU6xSkqlDBeB5ujxTpb2/ywEIvbo6kZq6dYxHaKcG8Avvq4AEwVUQruYkNwibVb53inOep682wVEitWkMru8F8fC3xxnwBHvUHkthIOJAaQP+EMVS9MuTYFJ7ifLGyXyI89hETy/jocK5fAWUiyGxNzIK58BL4APkHW9H/BQklFc/Bll19zCNXmGvW6bLIhNJXPI7khDG2UG1x/xRmz0SEmUsu4zZUHh6uTHl7H/eKDdULYWFxgEYGasHmc9an5kPDCOrLkkRd3Q4OYoh427+zhKCsF9o9Y135M0+GQ+UNThX2aQsqZhHxWDl7+3oxzscACYBw1Fjx4M3ghKuywglG+gg+VrYAfaJAfco+TaffYl5VLgs/h+Qjyzw++vXxSwqMY32zkFDIKSpftkkvCAVq5HrHP5VUZGi8hd8JVAe5N2dzcqkNRGQsPchACE1pBfQA6UtbU6yAopha+qdmcTZIjEea+DhAFGFQemBp5znJZyKd5jmJ7b22ITYKtA0AuLMCWNmw7NmT7dvb8ebG8YR9nc/teGMFKSbodHOxplBQpQv3i7o+NvBVgamdvVwAl94lnBsNRCitYnqmk2D0UM7CfPdDYR5vAp8K+GDJuP4MHdZNsMaLwU+YWlg6sGQBw2Ddw/wQAKhwML/HCwesyfmF0cjhtiDd6QzjYs0QHOT6bWGpi8nM4d4u86JAR5RCxVvF5ULtE45SDB+NO4eU8lzovMFHFRMw2Z9Z5aDsrh5hOND0KeYGPYj9hQ8fvY8ERFFwAfmLyS6Dk+4yC3gE5xHLB79wtBvkCkAP4k9ctID1NiQYazQQ08gyDZjow7VkTWasBgAF0S2K6lNUUk21cCApWkRwsTjig0VRySyc8mj3QmWvj0MmzYi7xOxw8YegQ7gdgxhwB9KaJLcubmjc45OGNrVhg+kWfW5kCCrQFjHY2vjdE63WdrPdaD8N85t+VaRDsW5hbkiiHZnEaRR+vA1ipHAy31ePfAPIjwId/71II8KpnCARLCw7JMM6VDwBTNWSWAOoeKC6DzZrAm/AzUUOabUO2b4HQwMDnnvP6zqKjaeF7EtaMDU2AYawlrpCRPD8B+J8SEKkcqmDNJ3Uc/rY12P/dOhBgp4KMncMCIISrgrBfwVoHG4k2hd8KcGpwJUSkPnHSH/fcrY18D4lbNk9jPrCyxM6viUmsAGx8b1GelkpicXsDm7IjpqYhygfUTTSDeAY0ib/33rv6+V//+lcCilKtzWLSppPNYoyi0uSeTUxMiO3HmgZIxxqnBqF82UvaU7O7hGt2aV7JIjI0g2Q3GY9JOSYGMrWVrDu84Y66g70V0Jj5RVMFNm2BdbsRAK5kDSEnjGemPbCEUsWZqVGtxh7H9wB+qWW4N3s0vJJJGz00ai9cvKhnxLNirly+fFn2gvydOoymBDUTX3w+WSCKFMA8ccAKOyDWKamMxGJrkPqyUlez3d0dNe36urs0PlArYO8BwA1Yhqo2lfL1mwUYMAOVAPd4L8daUrSmVNLW1zZkpcO6huqlJdVohdyOvXzpORvq77Frn16xi89f0Pp4/foNAecnTp1QnYiB0uzsom1tblhvX7+A7KZ0s80tzNv65rYIJKh+AHexdlEtI5Y3tjCMS2fp+oEVharXnB4+W/AaUu0dP9Cq3m10BqorgtzahmcCWMTaqPFIlgfWoeRFKUfObfwi+0nGkuxNA4gru6UE6kC3HBWLEeKGsjUgfLAOeyOZMdGSSiqAuT7B5/LmuxjmlKlV5z3uy3KIM0LN+gfabXS4R2skzzlqIj56OG1WYzxsWVd3nxQTNPCw/GH9wPZDYdJSWlcdwAw5cjs7ruRiP2FMcWdzBUB5wLSStTanrYgnNk037JRCEK6As3RKPto/f/+XAleGx47YwyeTIkERFL44P2cTJ0/Y09lZy+X3bfzEKbt9+7aAKr5mnj6148fHNY6Zrygqnjye1FrE2oENCbVmIl5njfV19q23X7Ou5ibL7a5bPIYysKJcudbOHivsY1NbtY8//tyW1rbtyPgJ1SQ0uRlPjdjdFUsCR+ShzXygKUjuTrAbzOez1tqGJR+FoelMkc8Vrau7NyiWyG9ifapado9GU8qG+Czlkm2vrVlfb5esbA8dPWqXr14TEJ7JF7RuYMuFjQfMUTWPoiwVGnClskB51lRshgD3i4DfYb9Jpj1zRCHHCRRLDVbDXqda1XN+NPlEtUhHuk05RlNPn9pONmc5wE725GCXQbOSca0mrVQTPj6l6tQ5BCa9rzWs5RFIo3oiWI1QX7mVnBPoPLPQFeSMR7dmdAWBZx6y5/q+gAc+gCjznIYOa6qyFKhD0mk1LThTML9hDsc4L9THrEn2QzV7+62v2z/+9KdWX89+XLTjJ4/ZxIlT9sH7v7Tvfve79jd/8zesCvbv/vD79uP/8Zc2cfq0Nbek7cH9u7a9RSBxwt5791vKh7n+xU2R4rZ23DZn/Ngxe/WVl+z2zVsCcqtGYzRudfEGq9XXWXY/p5oVMpNAy2w2kGaoGxOq72DVqxktH3XqBSepKceHZiF7dM6Ddqn5aIiNDA/ZjRu3xJBGXfrySy8qp4qcCld9+znRiWPeJKLhgtoUkJgmm4BR1aNNnhUQq1dmVGTFwnOk9oVGF9kFue2dWzTyfdUCkOQCmcKVMZ6R4g2qoIINEExk+eIWhOyp3uyKCCK8D+OA8eS2t97odSa/h7jX15Fb0qk6ancvp/ybYn7XMhtb9ic/fMe6WxqtsLdjLR1dNn3/kS2vbtjY8WNSTuztbEulw+vevXvX2jvb7dTZszpjALarUbu2YeurG8EGrSQQGLKTlGONSdve3FZdTcYC+TE0Mwn0rVZi1tKWtNfeeFm1Tv/woJWzeWtOkeGwYRtbGWvp6LaZ+SUroKI6ftRmZmZsfmFBz/m111636ekZnT8BbEdGRxWYHt0DGgGsPxC7Pvn0M+EMhHwzp9QcDyRVaihy29jD3LIX8NqzTIQfhTkqUio1rLLsWMGpTbH5drsuwHXOwGRzKExbuZXsnSjzPNh9oK/POtpbbWdr21Xw2HVR36RS1tLWqvqVZ01tAo6V2aFh0uD4Qr0TItWcrKtapZCzl54/Y2N97Tbz8K4dGem3XGbbRo8dsfnZedVb9+7ct4lzZ+zxg8dq1n/6yVV77rkJm56atTPnT9vM5KTuO3ZqI8NjtrNdsA4sKMsmi8iB4U41Kt54+5JyjV569RW7fu0LO3bivG1m8vaby9esRtB2a6dNz8yqTozyJDmbQ4Q4fOSwaqeNjXU15Hh+NDT4Yt+AqMYaxvyjNsNqCsUtneLMTka1L03vBw8eSlEhUsleTucT4UJgB9TAkHXBaOqViuZOAORGpdPW3NCkc8PCyrLtQyDhGeeLlqSJSs6ElO8xgfSyxAv5pazJPFfO9rJLDcQwlCD8DnVVVGPyi5Fduc49oV757dFUx4K0Tug9sYDt0pjjPMZ4Zj2KSLnsLbKpM1POidsm+pmLRosrb9wCHlWpMFECwLFjDkRaqQVFnHKiHipRzhWcmaitRXCSUsTxoWgd+u0/0//8J79qVPx/cRe/eo3fiTuAosL98h1gluVAiysQxP4CmwyhuDpA1TwsyzcgWK7esVW3UcALhYJ3C9nInNnum37EQpZFjAJM/VDGgSlim2oiE93GwSxI4WS5pAOfF6iRJ6nLgIPNE6BxAKn42ePj43bv3gMtoqkQxMU1qHjjgBY8yvm8LKYcyrkoXgMwCmZS1Axhp2UBjhjD+ULOCoRhxdwjnQURNQqfqYDlhsK/HLCj0OV6VSBR0MtSxz+bLFwUCuqLvdtw0H2tEztN3sldHdbb0alFkp+pWFxFCrYDSMrZECjcOKg4GOTgPGBJ9J5RE+FLpYMfNNW9DhZQ3sWOonq/LP5hUjkLAcaN+3QrO0DMJj+IR4fv6GAuACf49ch6GFYPUuKQOSCVQRhXkQpDFkKh6fBsdzgqPqUWkeWUM5a5dg7SHCJkqyNfVgfbxeQIjCCuD4BcXuQhWM83I2+U8HPaQHTY4HAfgXxfqlAiwE8gvXpa/ntiMMOkLwKUfvmlgliqCi+io8YI9xgQh4ILqxAOP1EmA80wabeVDO/NooMGCnOF/4PR/YyHtMCW0NSJnpN+jzJP9wINg+k9KSK4pii8HGANIIADNnPNmyweqgXo7ffELSfUpOG1uEfcf8nCCaZGedSiRgMglr++F/dcJv9VEUXRik/t9qaafmJUB4ULwWCNibi1NrepGKNQ6x0etsXZOVmdTc1M+70A3C+VZQ2HVF5yfgXzJWwFKfv2tuxxjh47Yk8eP1bhyvUBsvf19Qjkwh6FBgIy4IXFJZucxjvfZcxqkBI4bjVLAYbArI8lbKCv327fuSNQQpJO7I32nfUnmzJAPfxPA+sdEKwBxpFftB+IQj6Dg5DYccQ9CI61IgDN7lvp4CcWAxwinb2OusCbo1p/ATPDeGeca23VfCCYzg8KPE/5+of5JKArrKFqWIUAQ89F8IMgRRmNIexc1EQNdhuycQpha1FjTGul/KKdjaNmcC1YjYRAd88XAXZjDMEsLAjUjHx/oyJLzJZy0RspQIEC5uXJ5LZZjkBrneNn9WfZzXnRGAcYrydMdEeNQQrMbD4nixwKRQpGClAY+oCsW1sbAuEA+COfau6vH1zrZCnCGo3aR0WoeV4Fv8tzU35Edldz1NWEkRe8S5d1CNbc9TWPtUP2FcGSgsJ5YRG21mAItNN00s+zftPk4HAV2brJugXgp8EP99F4YR6xb3jYYL01J91ekPdnz/GmoasDItCauYDiL9HgChkBTSErBeACwJ1NTdJ+hSayZnswtfawAGhzXwkxZO2SCkL5QSaVliyigppFQGwqqSYNB21eh6/9/L7Gi/JQQgYJz5QxA4C1tb5xcMBiXxDDtlq1XKlg3d2darJCkAAQ4XmLVR6CWJmHNCl45uWiB3ICWtHQi2wkpMLi+cMi3s26+jIFQIhlma8Hau4HIBkLBGfdNnhz49lmoBj89WqIzS/NWW93j9jd5Gy89fWv63D3s5/9g/X29VljKmUbGzuWyzrowl4GuO9rva+XgDg0t7mvkQqOA6VUJ1qPyamg0evNCJ4L7DGa0owz1rB88N5mj6TZyufwHDK3wgQIAaCKBzYZTWjPIPI5rVot7E3Psu6jOo/n6P7gzLF9O4ZtxMUXbHp6UsHkqDwBKjhM4+UPO1xgvZr/4b5yvwW8O4A4P4e6LSn2KHsIzQiafLLmrBZlO8Se8ebrrwt421jfkNIOBhsADtYQVgOwSFpfb59bV0lFlrL52TnLkF+UTlv/4KDmERYAqGESdRzQy/bKpeesrlq0K5ev2WsvXxJp5Nr1L6yjq0vZIrPz89bT2y8A6NEj/KqPacy1d9JY3rOF5VXL75dEImHXlVUcbEMpfnwtlHKUwF2s7Ry90VpNo5n3cxs6b1ryDKSKRJnFXhAy5GSJKEu9ehFceI3VtVWNIXgUB2HdobnLPKdOoAkJeMl6CYizGwg6rC+MD9XXyjUBB3OVMF8o7lhbDh8aVRAm4eKoJFLNLaEBGhj3AnlRCOastTNp5fy2Ggu7qJaaGqwWa7AHdx5YvD5l8wvL1tnVe1B/8FkAowXMA0qTtZLNK2QeFjDA4cLCkp09M3GQr0HgJfWEfrdSsW1skVpbrFwo2PPnztlehlyHpNR1AGvp5lb7xT/9yiq1OhsaPWyPnkzJ1oSfWZh7aqdCo4K1+Oj4cbt2/bqNjAxrjk3PzNi5s2cF8rEOHTl8VON6bGzUCoWiraysqMHJFt2YiNmrL5y1+nLeDgN85QDU4tbU3GK485TKMYsnUvb+P31o++WYJVvbLLsXmi2tbUEFsqt1jfwQQDs92+DrT621KkvLLtny0NyBcFEolK27q0fNn46OtgCSQ9rat+7ODjVy+rs7bW1pWRsO4+vw0SP2yWefWwxlEJkqqgNRA5bVNNCooEmCxSx7IfUXewA1f62s9y8VCtbbhS1ORvstezHXCtBfzBV8zWpIqA5k36OhPjY4IuvMpbU129zdteX1dSuz/4XmiNs9OfnJaxhXCFEjaN0MhCLWfZGcAhmK+oB9EcCZtQ5iA6AdKgTWeM8j8jpLLP1ghwj4XiqiwiRrq85Gh4akUmPOEVhMsxJ7Xc/RADT1+oy1lnVaNmPVMlpwa29ptm+8/Zb9w09/IrVfLrtvp08fs+PHTtpvPvzUfu/779lf/uX/kBrp9//w+/bf/vwv7PnnL8hS5c6d29rTAca++c13BCZ//PFlK1aqtrK6JcCRteTP/vRH9vjhI5ubnbf1rYwlGpO2VyDgthgyljz0/OyZM8o6WVxc0L1jz3jhxRdlM6dcL4o8NdyD1Wvca3junefMUSuWrb+/T2v57dt33PorVm/PXbhgX9y4KdAzIpNE+Xw8b4BnvPwJRsZ+hTnCFzUK9z8iXTG3OR9EoKSa89g56+zvY0l2rE0otv08EzWj+F1/npxBg3Jd6hkP3vawZ2c1SzmqJieKRM/qiyynnMjnZDD2OM/b9LGnpn0CxjRniSbb2t6x9tYWa6ivydbthz94x9pScdtcXrTh0TFbgiX/ZNpOPXfOOru6bWtj3dIhc+7uvbtSd2HvxeuSqUOdtYul8+aWQN/FpSXllMgXv84bfiJwEBJerdkWqq5yyVraWFv3tIe+/Y2v29PZpzqbQZyBYBOLNdit2/ctWyxLUZHd37eRsSGRG3mt6clpGxgc1prL/Hj46KH19PVqT+d+MGaomSCbULt/dvW6QFj2Y0BmlMisUV6POynLg5C9mFGjsOyB6RE46yRSP5+zhzN3YbJTZXuWnUKNbHtrx+IETMvpINis1XGmrFh/T6+wDc5+stRWQrUTG2nMgJc4USwmG22IQ+y77R2d9vDhYyfC1MqGj2Qpl7c3Xz5vI72tNjf5wIb7u21zadFOnD5tszPzNjg0YJPTU3ZkfNzWV1Zt7NCoXfnsqh0/fsSuX31sb7xxToS34dERm19Ysr6+Ycts562nu982tzJSlTSlE/Zo8pFdeOG8PXhw315/83X7+598aK++9rJt7OTt/V9ftnRHtzWkWm16ds4GBvots7MjElI0DzjXUC97HktJtbuywEQwxC4yrzqHfQSsgzqfvbF/qF/XQP0NoY7g+0OHD9v8/LzO9G6HHDAg4TTy6bQKXA81KqrWUKtZe2PS2lIpnfM3MtuWK1csLxtoyFPeJAK3cCKs17XUrJB2ePYQv4QTqvEQwtitTuOQ+aQckrDWK5uRPQYsIuCGfpj+bb4CbhKaJNS0qMpouop4KyvQRd0/NWHDeY3ro1HBmiXsBmvLvexBo0JE3XA+6QQHUMMNp4CsLK04i8rcOASgc56N7GdlU0gGS6EgzELWp1ly5IJa8F98rEC3+20+7D9TZDyLmX0Vpv1b3b6vfuh36Q6MwcQgWBWgDWlpd7esPCKQgk4tYAebg3IjWMKqHqLJF5tOFMAoZm348GK5w/YqFHQwZFHCTgn7IhYvAEd2FF4XEJFNGLar8gjqnBXHxkXh6Q0NL3ijrAqKZLcJcVDUwz69wOIQ7pJgZ7tTeLDooWig4EJCSWHIZrawsKIDhuxUgtUBwJQYl0WY4M36rFxHe0eHCgMWfy3w6hw7IEgTQ0zdimckiGWiMG2KWbfboXDy0FwsSvgsDpYJYENGWSbrAtZmweoApSsl6+vpsu6uDhWaxf2y1cPqzrglU1MKEAnmS1ye1MUSTBEOut5McBDKWTOyUwph0AqwDQslxQAgkQ6J+x4KGoGc+pmQ7xABc5EnfZQxwdgQ66ladjsoPkM6FawJ2KD2VZRI2gdQgXdhCE1m8+Jwwo2MlBl+KKMJ4syXgwN7qSiWlYpiaD6h8+0qQd+gHACohgBR94CWr23VBAZI3quOvzdkuCY2D3lq4599YMeTl43HXiYrv2gOWWy8UZYC4DXPiwbbxtqGLDS4hhzhlG2tkkL2sKGVimIuAU7z/GHJcBARwIyyIHiVI3eGPaV7A2AkYNvvgcAsZX4EQDo0KiI1CffWC0P37o2YCLC5KCT4PQ4aFImyQttzKTR/ZxwAWnDfmFtix5MpIHa7Nx1h6Qq0CI0c/ivLmYaENeCnX9rXgZo586WlDvYV9ZYr5NwmLtHoTN+aNy/5/Pki8yJp++WiQAaKYr7wTm7r7LTrX1xXIRw1vQRObWzpfSncx8YOWU93l37m08uXZfWB5BYLEBqNhHACZNZqZR2mUUtsbWzp4I1n9erGpq2srenZyI4IO5VGMjlSKqymn0xaMtEoie3W5rbt03Rpb7XFtXVrTafF0Fzf2LAjY2M2PTurMQIQNjM7rzkc5U/owER2RLrZcnlnqZ2amLDh4WG79cUXvo5KdhEycQgEpXmgws3nAvffFT8waB1s5P8jdpiUU+YMVGAEwGK3EvpyTMhKgdcKjGn5mjY2aE1LCzQaAAAgAElEQVRUE4gGX2CYuIrGszi4KsYp94X1g3VnZXVVzaL+vn7r7evV2gFzb2l5WcweMXSCjVjEohboX0OSvmc9Pb2ay2EoH9iN6VAJW5ZDJOxNbBjwIEblhjotEwLyymXrUW4B1gQFzS3WX0BuXnNhYV7rIuwZDvesQczdzU38WrETADSNa37A4KOQB4xpCM0c5gXrBk0JDvNq6AX7Q3IDkGWzbnvOgTNg+T4y/gxWgnFAFRQz0Z4EW9/tcmDj4nff3dHp+5QYsx7Ixt872j08lfEjZiMWNRHzBwVisaTGKI0Yz0NCbQaQ6aG5/FtTQ4P2cRXSaoD7POYebm1thcZcXGHPs/NzKrwBXbo7u4L/rbPfnTXkPuSS6+PJCitpdU37Wlc7AbFNahLRxHO1C/ZhbinB2IHVzn1iH+X1aChqXyzSFKQ5TFM5hMyVqwL2OYBhbcA8gv1PUw9gBSXD8NCgwBH5ZEuFYrJLg+XKPjs9M62xQKgkXtzUEABS/DzgEw2nqGEGSO6HhpoaRIxfgnJX19elQIiUGtxTZYoEyyd2G547c4e1vq29RaDxrZtfWE9XtxQjsbqKffOb37BDo6P2xY3ryobAuq1aYyx4hovsHzMZO3PmrIBP6oojR44YRAhfgyvan8o1f/+1lRUdSGnUMFcBMxizHMaYMy3k5uxu2z6seAXJm+YMa0FfT4/GPDUW4xlLjt7ebrcAiSesKZ3UfXfwx9n+NBa8SW9u24FaAJWcml9l7fMAqSdOnbRLly7pECiWPjVhaEBQ0zx+/EjAKf/Husx6C9AAc1p7fDxhT55M6rqUMyVYtE5KNg6G7FE8a4gaL754SQdzPjvXTb0IGIltEms9exCWPqhOxN6MeR5T1ODjmll7mZs0KzZWFu3I2JCdGB+z+lrF7t+9LfYzIMsH7//aBocH7diJ4/ZkasoaGtNWs7h9ceuOXTh/Uk0tGKbYFhJauofHP8AbgdYhr4tnQANYFoA0hnL7aswCqsbr66RwYVxGllAorlSvVauaM3zfG0dug8aBl32cz8/no47mGfI99mzqGPY/1lnWAAf3nO3n+Rctek0y0Do7O0JtUZHizS1Wg8+0cgJQ8+VssLfPvvu971oht2e5QlZrm2y96uNaU/HyJwsmhyLJinb0UL8NDXVbZmvDUq2wj7GPqbOpyTmB9DTqaNqhcIQ0xP6BnVK55P7WIm2ETIBojgI+qm6QvQws/TqBcxNnzsljnRJ+a23Djh8Zs3Sy0ZrxtCdzA+s/chEaU/bz9z/Qa588OWF3791TUDXe5lg3HTt2zMiXYj0+euyYwFwaVHzxPmRUYJ3BvGT8YEXFWsEai6JClomASQ0x++bXX7PBnhZ7OvnAhga6rZDPyst74NC4raxt2+bWnj18+NQez8zb2NEjOiNhuzY+Pq58FcYJjZTBfhQdfp5gjdrbzeisQFMAxRD7N2sIOT6sTYz7SBVO3TC/MGv1dTXr6e5U0O/ywoL19/Vov8NSE2Xp1es30OdanWwWC7K4JKcj3dKqP7PP0VTA85yZmWBdwg+fJsV+XlZ0wwMDWpM3trdkfcj6DtlNXvQw6Akrjdfb3NySVVAYjByRFdfUwpzVYcPCPlcoWB4LMWWzOItV5zHq29DUE6kqqELZl6gPIhKRyBgAzFZnO7t7qjVo+rKG6wyhXAUUnM5+jXL8XAlDnezKYObBodExERY4mzKG8lJ/osisyn6QPW91bV17VFtri9REMdTvrc3KM/jWt962xnjMbt28YffuPLSu7ma7cOFFu3rljn39rdftL/78vxv5Pd/73nfsr/7qr+WBT/116+ZNEXUgEX33u++qbv3ok8tWqtRsaX3L0s1J2A/2pz/6kZpmV69ct43tXTWa9lEZo8iMY8HmNeMbb7yuMGAs8tj72Z9ZP7+4dVN2tzRaRTQR+OwAotStUl8HC6dKVeO8s6Nde5STRWp25swZu3XntucdhVwrnalQFbIuK3D7lIDi/oFBe/jwocYp1lrseSL9SB1RFogIkMoz5D5DBvDsC68juUZARM9bc/vByHaY8c798kwsXzOpQSFdYAXk53O3ImYNkRpDinDPAVImFTlOAkw9J9Kb536m5J5hedPZ3irgfG19XZBsS1Pcsjt79h//+BuWTNRsd3NdDfIHD57Y/QfT9o333rLWjnZbfjpn3Sg/6+rs/r17lkg22plz5zyHQ+fFditIEZXX2s75GXtgzqLlQt5KhaLNzs3b8eMnbW5hUQ2KmZk5qXhPnj6phsHg0JAtrSxrXceeKN6YtszGjk3NzNt2Nmd9Q8NiynNGkJUiyhXmeKpZtSZjhToYsBZ1F/eA58H5YXZ21l544QW7dee+zc2xfruDA69DrUedSF3hpCnPTmD+8jxQM8piOVjfCgtQLqjbmpJvBBZA4xWVhNU5cY8AcRoVOGsolLi0b8kU9VdRaifOHY8fT9lAb5fq26HBwYOagHMK95H/UZPRmPE80jrbzmT089RArIt1lbK99doL1t/RaNnNZWtLJ6yG+r+lyx4+WLDRsQ4p585fet62VldtdGTE7qNKOHzY7t68Y+fOnbZr127ZsYkTdvvGLTtzdsL2sgXr7e6VMwDql91d1vsNOzFxyh4/eGRvfO0t+6sf/6O99Mrztrdfsb9//3PrHR6wWqzRns7PW1//gO1sbUnpR23KfkRtiguCCGlYoFUct1CjQniNZ05R47AXDY+M2MLKkmoX6j/GPbXn/Xv37dixcdXIsnnDLlLWXU6KxN1BWXWqGXC0KFsDisRE3DpamrUeoyYg8wTiLpZbrNOMFVlS02yqT6ipuI0NV5g/ItfIYrZRY1B2yWCKpZLO73zGyGFD2Z8h6F7qiODw8S8x1WeBeceMXBkSqbsYc5xDOHdzb0T8qa8XmYqayAnRbkWFGohzV2TpDRYaKbTcOYE8JrAVVLwpNfYc54EcvK86VWM7WH1D2xo/Nq7mH3UzjUWuh/vHM2Td5dwaZe7KPjzkxfIarFVua+sEQ77PV9S4jRrDUZNW5/9nArq/alT8LiHwX13rb3UHjmJnoBArQjDd55fNH1YgxS9dQm1OodNIsYGEPmL2il0eGMlaRMNEY3LxGthy4JWtMJq4A4HPdkoj1m/UdecQhJ2CXlds32BYFBinEahxYEXkU1ibKoCLe53jfeie4O5/6QsjXxTpeFdzwOOVKXzEnhDzzP/n/ugOVgmwI2Ba6hEvhgXIwPIA2JY0bM8tT+qCV7i8lv06AFgAeLi/HPp0LUGpojBnvIsbkJS6pLOV+1Pat8LerkKZ2MAl20bqTpPHWOhKYvpWqhHbrs62tgDgeI99bQAe2lnUwYHP6LkV7itPYRE9N1mgSBriMmUKEGUjhJBWD0l24CCyAhPoqEaNZyOoAy5GRUygLPePwovvwcQHqIYNEYXg+qHcg13Z8HgQyjcIXXUxBkJIr4+LqGwM1xIYVXwDxl+0gEfjj0LZGZwJK3I9khp7IwhwkuchxmiwtPlSHYSlGH7rMDtqYmHzOmICi2Ho40OMZSxbxGKMGlN1dmL8uArA1ZVla+votNzeXpANwuKoqlg9YLaiaDEPvWNDYmzx+aOsFFjH0f2KJrJY6FHuSGAbiYkULJ64NkA55ithUth+EFJGkcKBK5VM6z1lZ7SzLf9rgjTFaiInoqXZ7SVoeASPdq6HA5zsxPQ9P0BQ6aQS9Zao96BgMc/TLQIGqC0AiKWukGLJN9pUY9pSTSmF0iHDBbwFZFHWQWDwSw66t2OtFMpYv5gXZcheOTiSG3Hk6BE1NJBEc8iH9UYDiGtFzcDvFQo5a4xje4U/eVUH57XVNb332NGjtri8KvCJgxKHxqiph4UU1la9XV3yZIZ1jbVHGQ/q7m6BpTRRpZYpoXjqsc2tTc8qqSP0GQWVs4hkX8BhK0Y+gD9nnj/yXQ4F6xtrahjJ/gkvfrG/4mIEUSrqfsOcDs0ovMB5VlJIheLSPZYZS+7ZzPiWOob/C8wmPa9gzcT3VAAeKB1cOSa7NgVxAjQ3qFkdMU4kw6+4IomDJkHbHO5gT8KsZ8wohDFIvQGjAacBv5krPDtABclrc3nr7ukRSMj6yTrAerG6vurWVhxKCAxGCg4rOVyT5oY+mzNRWF8Ax7BryOX2bWhowE5NnBLzFnuDx0+eaJwyZhqTqQNPYwA2qYUU3Omfm4IfCTUS9JakB08DHnKozRayWkNphPH+XNsyh7lgS6X7SYMj+CerYGTNZE0M2UyRCguwQJYeKCQYpzSSQhNdAZYK7WbNQiXhtok0iwi09r0C5cj2wdhjf+bZMQdc/ecBuAwEfKp5vc0N7A8BOt2WSet7aK5rbwIsDk0MDi+y7dovWHt7p49p2WWE/RXATGopD63kizBFtwHzQFzWWEJX/Z64As3Vbp5jwX1nrOCD7fMl62qFeELgO4dX1izYYXwBMsp+IezrADnLy0veGIIFhYUEnz1Wb5ndHc1l98x2/3EBMOWSdXf3eHaVPpMJKIGVj+94a1uHWP/cP4Bx7rEsuILdBHPWGzVudydmcDqt56H9DpAyMNOYyzSsAKqOnxhXM4h7Ojc/a3Nz87LwwI9dIHMDHv6AM1j5kCNUZyMEbSqjZ195DjSqxKYDdJNXeNky2xknHeBrD+ASSAbsZxub63J05rOwFnGI5PN0dfA8fa8A2KHO43DFM0A14JYcsL329DzbWloF9LjSwhmr7LM0nhYW5rQ28N4AAVwHh1BZehR8zlMz8T81FfI56+hu0xrIvsnBmX/HDgoQTvVlPG4PHj7S/Oe+sAhyCMZ3fyuzrbWQwyL7tgOgXs9ov4T40pjQmsHc4j3kh11x9Vm0J7Kv0yzGJmtgYEBN3eXFWctnt+yN1160WLVsv/6nj+1b3/iaDraffvqZ1usj40eV0ZHfr1m2ULLZp1N29NiY8pa2tzIiQmztZK0x1So2rAAKZR4lNaa5Xpr5zAsO8zxLxi1rNGAz1x81ZaMmMfec8QfghuUI8ySy2WOO69l2dmi+8z0mGusLYA73M6pnmUcKzU42+XpYKCqDQGQQsYqLnrEEgUOMWHI7yC3yIPmNtXXr6+6zBPVjPeAU4fTkK/HnYMeiGpPmHGtU2c6fOWZHR/utWMyrCcnaUKzU2YcffGLdPUO2tLRmhw4fsamZWVkYUfvBHoexnGxuVo4La+fc/II+P5kYMHxRX/K8eTbU7xB02ju6LZ6AhLCpnIBsZstef+Ul29na0DhjXDUl01Yo1+yTy58LOBsZHRFwSg4TwMPTGaydTgjE4FmMjY3ZRx9/LMsN1mksofi32adPtf/STLx3777+jfPB/Pyc+3FbVeqRSxdOWVsyZv3drZbd3dQe1Ur21G7B2keO2M76jr3/wUdWqtVbiuY2Xvx1MT1PDxoFJHLyBHOJNdWZ9jk1oWgM89mwIeL31tfXVGfReAEgYh2gyd7X2yOrLvKWxo8etdmn02pUs4byOVD9PJmc0n+ryuhTJ0DzDQUKzV8IZLBgUdMqHJt6AzVcad/On56wunLFdjY3tS7OzM1asVqxdEva9nI5kX28sUnjKG0z0zMK3r545nmbfjpr0yvL1og1GOSj+rjARUhqUomHcRw1owHOZKkaQE8nYaDAieye3F7Q99+QhVcHaSOl5o83mj0rTWtE3O20lCknSza3pWMdhwSQz+6F84wrFsmfoVFBA5jzpkJ5G8g3w96S81TJmhrqra01be9+622p4Tu7Omx+dsZyWZjoKbt2/b6aGD/+8V9bQ2Oz/f7vvWv/5X//c3v1tUs6q9689YWeIeDWe+95o+LDjz82tBoLK5vW1paW1SGNitnpGbty5ZptQlprTFqRkjxkfLmpTp29+eabNjU5qfBcd0eoU0P52o3rB80vKbmoh4I1rEBmNZvczonPNzI0rKbmvXt3VSvRqLnw/AW7dfuWmseu9nWiDfsE50maBmdOn1YeBOMakDuygdZ4xgoZlVtLi/6LApL1SK4CFVdyR/71PCdwgwOb0YOzWHQycsIiY4KxrXojKHs4V3H29pBuz0GiIRsR9RYXvZbg/bxx48xoAZUQhHT2qdrwQL/qpqXlFRvs67X8Lvkvu/a//Ol3rCFWsszmmvX19NuTJzMKSz538awNDg1aMZeXPeDq/IIU3M1trXb85Ek/E9VqspHNYhsorCJrOVj4jQ3WQMMpKIvBRGjqz8wuyI5t7Oi4rok1sau3x7r6+tRAIY+T80w8BnCNPVvNcsWybYvkUbGB4SGbmp5WlgT3g/Hx0Ucfa5/FUmxgYNA+/PAjWf+9887btjA/L3D7ve++p9f/7LOrquG0z1SqwiHUqKhPeA1SBhPxPUi4juaa26vxjOWYkPB5DnGV9YucUog0KPR5X/6Mmg7QvLgf6mNhLTy/gnV1dGhOax5T8+3s6KwCUcwJo2SgYjtLcyMl4lCqpVmKiqdPZz1nA7JXtWSYj7795ouWjBVtf3fd+jrJ8SlqTyFzqjmdlPJkYuKkSE/HTpyw61eu28Sp43qtU+fO2cM7d61/oNeuXrttExPjtr6esZGRIdUxjOmGxrjW5N7efpuZnrdLL75iP/3pL+ziixdtfSdr//DLG9Y10GXxZIutS32ETdqSGqV8FvCrkbGxAwIICjWRcQuQVNztwOt0nEn21QxUfmFuz5rUtGEPjmn/WFxcVug5TU6WMc5n3LsDLw1lzbn6k7GZiJnwk46WpKXZb8icKldtHcWLiBaOj4EbUC9Tk0h5EHc1E7Ut85s6DBU6TSwnbKDC9gaAqzpCHuaBGj0oe2Xj+a/DmFGjwhuZwf1CdtDuLsD6h00hDX0U0TRFWVtY37hH0fkKfIpzwujI6IEltVTpEPiCU4FIWxDCAgZKM5t1hDoyOvtxodR0fDaaQ6Ojo1L8Qipg7pD36HlTWJu60j2yvIqUtqwBnvnmZ9Tos0WNiYh46M0MV65o7Q4KyQOc6KuMit8K+/7qh36H7sCRIIdk4AMi+MHOO44RqMAmxL9TUHMoBwz0jdZxU0nbqzQp3COZBUz2ToGh4cWdF5rOjiiIyeR+gS4F/LJriEe8y9EE+IQMCIFz6oC6DCuySuAgwcIqH9MgpT/w2ed6ZKcAk6Jo29sZt7BAmaFNEUYYMruQuSFPfZcUAgKxkHrOgIfkUkixucLQY1NQHkcA+NhU4vLhczsYrp3XYcFzcOhLnzov6ABTCyqKYFVkAd7KBD9iPVK0RsCh0r4OG3hiUjTJ37xCg6ImJhoALAd0CuedHUJTsXyCcet5B+4JXiegg8KcDVrsZHnP+kKoxpDyEzygTosfnq4csEMR74i8KyHU6ABUC3YfYtEHRri/jocGMw6UeSCw2RnbkR+zNyJc6cEmIBsXAbrhHgUQUTI4jSFvHnG9kpeHRoouK2QzCNQKYaSMR1g1Uo5wDUF94TkRHvArW40ADvL+/lqwrwAvPZAa1pn2ydAp8QYVYI/fi4hx7ECyP2+FBeqa/bDg98cZ6ljZREwVlwr4QuHMXNhk2Do48AyDjrHvNlcub9alhOuJ7v8/28yC3VZ0yVQjXKveU8EOrjCR3URxP1g0+Zj37A/3D3XFSQjBgoXGHKUoekbFotcxrEXc+oYvmDasExxkeK4cVgBNmG9cOSBezOLOvmBNqHcAmHHJs9ja2nQQkzGTSKgByDUBTDAHM5m8jQz3izksSWtjg3W0tgdwqt4VAGIXOCOkgQJYqixAwYSASQ7QqZY2BWItLq/oHlB0M2c4/AOswLguYJETi1s/QYA727bP/YvHsOS2GsiUQEosMNIHzKFojYxCkSOAljlAIR6Br4AiNDb5/srqiuaJg0zOCKaI4f5Q6PHnyCKERoVUSaGR56A9yjO3DYl8e72QQjrsa7QOj+HZsO75ePKmmVvgwDBk7PuAjP4uUCAErY6OeeHlIeyuDOH61JwUm6RykO9Dg5pr6ezqVIHvbEZvgiqwNSjMOMSIRVcs6Zmzt7DOApDJRjB4UnO9MG8AyNyvHVA6o0MNIBD/RnHe1tqudZGxzBqtcRiUgsxNZQw1BsCOJgDNCBrRqaR1tLTb0tKCwEXmAPNQAYXJJssXaV6xPrmiQd9XA64iwNX3o2DVQuM7AH48E4BzZQ4c2Bh4IzAKmvc9y/MQuD4YwxwqZJ2GkqU5rWaW7AEhCTQ1BQUL6kNXkmgfUT4J2TgetuzrvDfnOWDQ/Pbgyqyz5mHtSIWIx70HUMKOxkaIr4hZr/Gggtgzg3juUXOUa2dPInScfAHuB4dInj1jBMDbfdZdrYnqiu/xeTggsB5GrwUwzvWiShNQUHTvfdYDgY1YKYaGCZ+BJsXWJoCmH8K4/9wv5nPExuQ9aaQAnLA2yI82JItzlIG56VY5WAMA6O9ogY3qHGXjaO/60l4wWou538xhrGW0F9A44LW4RwKN4/bSiy/q0Ap7F7XG5sambWxt287enlj4Yv1XKrJr8CBIvHLb9QylAuH5VLwOkYIu1DP6PeVIJDS+V5aWpDBTsGIGQL0gMgksVAABxs1A/4Bt4rmey4tdPTc/Jym/N1YTClalxojsoXRokrIv1E8hNFMKDykvYjqEMm9pWKjBRo5IwfNjaFKgoFPuAXYEAMsxE4Dqoek+p2lKwHhkj0c5cev2ba3haqa6cExjQDkMssbExisp9QAWRNhMkaWkgF3RODwvSfumAnm/zI6SVWKNoOJVrWXd7Z0CLGZnHtv5M8ft8OiwffjBL+2FCxetqSFpV65dk/qrq6dLe0Uy3W4PnkxZdnfbRkcHxcRDnUfmwtrmtuXyZcvTnFY2GOG7CasUPd8MoA/QgS+t4zH/jDqEBkWwPKODlYZnRvmaw8Gf70Xs4ohcIy91rKREmHGlY5TfJmtPmpOoWwhIl7KKmtABXp9bgP3e4HZwvKq5KuUeVkyQPerqnQxCzZVw8Ezey2XsOgK5p8o+gz82Dahde/PVi3ZyfFjgrdfDJYs1NtvNq7csmWyzzc1d2WixB9M4AoCPLMBoKm9t72qsbG7tCOxmfYRlOzDQp70QULmnt88ePZ4SYGJ15GfVWwWlWUO9nTpxTCAvhpkAdLBUM9l9sdNFFOjttcknT2x07JDu6dOZGTtz5pzAVO7DyZMnpdIEaGTdRil0+NAhAUg8M1SWjx49siOHj+iZ8n1UbNg/pRri9uarz1tzomaxWsFSjTHbzWxbe0eXNaTbbGsnb3v7Vbv8+Q3b2iva0OiIra2ua/zSkKF+5znNL8zL61ys16DsRnUBs52xODw4oL0KcIS6gufa2tKs+cFn5DWYJ1ub6zY6MhzIDTUj32JlmdyALq19mT3UNRndR9Y0xltmb8caGpKuZhCxp8ktVTnrMQ4gqTTG7ZtvvWWbrGtLi6rFJmemlf2HbVSZM1loVPMwAf+fzsxZe2urHR4etaWVVdugsVQuqbbSc/QI+KCgCDZB1NqBKMd9iOaHAzXU8k6mU66SbDBjTvSQzYhn27EG0LjX2o19bQiTB9RylbbXSCJ01dVZZ3uHNYkgUtXezf5D/Q7RCHssamnOV0xckUc4Y5X3dXZjr3391Yv2q1/+xi5cOG7Hxo9aS2uzLc0u2b37k7LJ+9k//sKaGlP2/d9/z/6P//rn9srLl7Se37p1UxZtXMd7737bCrmC/fo3H1k1Vm9PFzetszOl2vM//vGPbHpyyq5euWHbENyoJdEUxbyRGOXOvP3WWzb5eNJmns4cEOJeuHTJrly96ll34YwiopOU3DoFaT1Qk18kiLyNjYxp3N25c0f3h6b0ufPn7MrVa1rzHdj0LB5vHvu58szpCVedtLfLbsYV8hAh/L35XZQNNOVVn9UYnygt3faL/YEaTSTEQCj09Tw6pzm5w+tbtx/i9fiK3Axo0vrPuIJD9b7cFVhPUVkkdW+U2RHU6/x+VFdJlVPat86ONmtv65RVDZkvu9ub1lRftP/wR9+zumredtZXrbuz2yYnn9rK6roaFdQlNPGwgNrd3pb1UHtXhx0/PSHwlOtqijfY1sbGQbh3lUwIAF3skIpeK3Lftnd2LRYnXzOrP9PooVHe3tWl+dHQnLZYjMwYzp8xW13Z1J6UbGmz1q5uW9/asua2Nrt69ao9fjxtDY319kc//KH97Ofv29rqqvJExkYP2c9+/nONxffe/Y7NzEzbjZt37dLF8yJ6/OrDj7TfQGjlGcqJQPuJrze4BECuYM5A5ImIRtxX6jm3YC6LqASGASmC+oKzUWOT20A5IY05iVoyzPEi+Spuodrb3RksCuukrKepA+mCWlMqEQK2ZVnK2R/Nrqv0UIhNTk65ohxL8oa4VUsF+9bXX7FKfstKuW0b6Gq1cjFvQ0MjNj+/pP0dYlFfX68tLixqLl/57LadPXPMpqdn7dw5twMcHB6QLdqJkydtbnbZRkaHVe+B1aTScY2tkbFDtrK0ZuPjp+zDDz+2cxcv2tzSmn14+ba19fZaPNmstVgK/HxejV/OMqrxsVYKezRjs4WzAONBTXsaM97ko35lvWttb7ed3R3VUfyegqsbG2xniz10QJlLzD9hU5ryjr1IhdCUlO0R631LOilXj8a6quyZnThTtN1sXkQ67iVNJ7A8aoqDRiKqt3xBTcze3h7VJNQvUtmV9lWPcGbhPdl7WNOF84UsExFHwxyO7OEPQIbwh3+tUeFYEXiiE8fIG8T+j7mG/Zw7o5AbAR7mRCRfBGtSSaBURjHOfUClK8WVrJt8bZO1Wfi/KEOHcUdzlGccWQtqDMoFgAZpkxo0EFVQXrDmzc/NC1PQz0u5DG7i2XBqUKhRHzJm/5Vci4hYG+ExwsCeCeb+SlHxL0fLV3//nb8DF/v6go8+3dOi9Q/0aRMXWIX9RjotZQRFNDJBOtQcPPf2PGAGWS/FgcvT6ezCRncff03q+pjUBxQHgAVMxqiYEpMreBZKugbjnY49dhAHILJ79gIgRuC3qxXcmskXJ9icaf8yetIAACAASURBVC2O6ggHYJdr4jOw+GcyuzpMc03Y38jaimyOEKJFQSB7lRh+lP5aXAuLluRfQZ4GA1OegKhKwiFMYbcAsjH3vVTAJYs+m8OON0e4j7CZMmRmJJvEEJFXfLWqIo1CmMOlDqgspljj4EEL446OuUK6qyrMYZABbBL+KSZXDOCZRY+mROQkU6fCQWoInYUdQFH3WgFADgyyCothq3aHh+LyTHiuYv2FYDT9PEw72WgAdAUv9mBJ48GYwVMytMEFdgdlhA5Q4f5HfqT815UUflh3Fsw/7yYzweRfqd91Gxo+u1ixganP68o/HVApAhgpQBXe5MHWAD5ePDXKDkuszFBc82euRaG/qAMqJfn8EgZKsKDnhPvmwYZCccBzpAHhzHTAccCpiD0CE7Rb9w8Q0O3MkDTGNQ4A7AmQjIJmnVngHfyo2ca49UwNt6mKclqiBSfqqEcNMICtKOCdsajASRU3HiLlvr4lD5cGuNjLKtOBjZz3pqCH+eGMzoKeh0KBA0MKlgsbv4KyZM1TEgOVMerAJjZnLiVnU2beCwiR/RRhhBXL7eWsWqpanrnU4J7vFLOwdGF2MG94X0CUxZVl2SEIOA3jFk9p1iEaG4SEUThxD1054I1KhU/W05CqExukxLqixlSdNynS2AlUrXeg3xYWl7UuUMDD9OEL9i9ezN3t7ebR4HU2Pb+ozwLb0xUVrvJw5pZ7ZCsInMOUZOluWca4kt8tYBNZCkElwTrI2AJI4Lr4XNhIAdbQ5OVa8EIWOz4UcXq2+O8CBCjwL+4s4+DnCS+GAxxzIb+HFYE3Ivg5rjfyLtecR80UchNUGAVlUNQwhp1E0S+mfFAlnDpzRuGAH3zwgT18PGnNwVKJAx2AJ5+TMQVQKfuh0PyNxue5587rfaYmp/XaXGtra7utrK7Z6QlnmDFX+OxR4aVwRtkLug8razxjgfWWsZZMNugZc7hlXFMQTpw6o7HHGJ+ZnVWzESAssk3BI3hjfTPkecA8rtrp06dlqyObiMCaEaMP73D2ngQWOM7cke9uU6PAJYpYDj2AwcwvPruuP2Q5ucUa1omJYNcS7OtC3oiAYBjigWWja8znraenW/eC91ldWRNQy89y38gQ4Q1Q4MnaBHZ0CKhUsKCaij7m1FShCA5CLJ4nBTKFNd7quf28DpnRPsx49swgb3z563hegR/+Q8C08oocFPX70aQGEM9BAAO2i9WKmvzekMcruqg1hv0Eu7V4wvc6QArZM4SxTdNDzG/2uTC32trb5Fff0o6lW4tNTs7YQH+vDmbMNe5TtP4IUIVQkEpqPNKwognC9WANh3IGgJ/9EtABoIL5QKOStZkDsQLJa25jxet4I86b+Fwbh0gOsNozxQKNu/KA+0TQIA2cXNa+9rWv2eEjY7p/i0sLCjHFY3ptY1NAO+/LQYZnCJjNHtfb0x0OfB5kqpZiGHfKMGlptmTSmdQl2IGsqwC98ntuU/PgyvVr1tzqLDfGBPeDjAwYkhyWnr94we7dva8GDmttWxt5A7DiKzY0POQ2WexTuazeR7ksexkpDFGzeKh9JWSOuLKFBiNrJ40H1iXWBBoqWEoQfD566JCaOkMDg0FZlbOpqWnVRyj+aBxBAvn4k0+8+RpsPrm/WtfL2I85lgYgyyGY3RcLOK5Hz1F7jis7djPYJtBEc5UgY3dpaVFgMvOaZzKCBVS8zuamn9iZiWPW29lh7//j+/bd974txuHnn1+1nv4+hbazH/X2D9uDh49taWnFnrtwUgHfPd29trq+Y4uLK1YXbxQzfBebN+YKqsygzPLmOTYr/nkitVIq2Wj9g0M2NzvnILNINc4MT2PHpZwiMrFi+jNMysgKhZ9vaWvTnEUxKgUT2SFq7GAv5ay9qKHJOFtb25AajvlI0xjwKE/waDpYyQH4SvXUpPeSpWO5IguXphBWLoBKzapGVylVylYpASrim521b7/9qh07NGDFEnYtzI2EbW3v2eXLN6y9vdt2Mnnr6uyVVZDnvpR09oBdTJONpiesx2KxogYaKgKshQRmViuaI7FEXNZRaAe3d/Y0xyElrMzP2tnTJ62JWgx7CRTMjUmrxuL2i/c/0Gv09vbZw4cPbGR0TM0gbNleuHhJjQrm+uHDh+32nduy6aN5hr8+Vg6EmLKHw5YkhBZLHPZxFA3s23W1inW2N9vJY6N2dLjXOtuStr2xJHsg1uv6xrQ19w5bfm/f/uZvf2rxVKslgtoX69bRsRE9PxqlPGPAdV6fOiJiiPNvkAVgc/LFuKKG8WZ968G4osZQQ7wAiOUNJs5xjEu3ZzQp4Dg7KFOIcxDqwyYsoLJuPSM7Qc9bCQEoUnzTEKoVi3Z24qQNdXVYo9ixBWVNcALY2t2VBRqAFnkOPFdUpA8fPBSA3d/bo2e/Q04aqtFkUiH0IFXJJoBmiEkJnVvEqqd+pjZU09zrrcinnX9njYI5THFKY1R/xhoXZYQsTr3OZMy6Sh41kxuVylpTIJ37orOGY6eXImcsWLFq/adh2pSU1ZvyZmAQZ8k/pA4sWKIeBm+jSGfffOsVBWZn98o2NtxhX3/rNeWHoCoCDPurH/+ttbe32Le//S377//tx/byqy+qHkGx0Ex9WirZu+++e9CoqNTFbGZhwxsVlar92R//iU09eWKfX7muMPIa2Rw1ztr1riROuM3TN77xju753Oys1o6W5lZ77vnn7MqVK6rRBG4B5gbFrggWOChojcKWEWV8zo4ePizbkrt37ohJzD0/c/aMXkeZOWIle9C1n1YcSzh79rQyKgYGB+3xo8farxmXjC0AbhrkUSNZQds677DOsT46aVK1Xx4PfvKKIDSS2YY9qKs2HLB0lZ3sWxsI6fWmBXWHqyE984K9nPtLE5lxwfxQVofUZZ5zyC3heUeOCtQ2NPqxfmIdwzJxoK/XYtV9217ftP/tP//A6io5293asM6OLnvyeNo2trbs2MljAmm31zeksCSr5+bNW9Y/NGjHL5y3/NaOCDqcqZbmF9xWEuKQzv5k+uEW4Ixy1keaA5xFyUGC/ML45kzL/KA239zZUWg5SoTcHjltRcvs5qyG3/5+yda3t+3EqQn76JNPldXX1dVhL1560S5/9pmawOPHjwvMvXnrluoRrPjYX3WfEvVqttCY2t3NWjoN4FySvRHPKlJU0MSQ8gECYhGFUZNUFYw1npVcDJoadJ9W1lYdf2AuG+fDsg0O9mrt2y+gbqLBKChWexX1IlZEI8ODIiYsLy3rtTkPcb7VuTkWs6ZkSuQvvqhhRHJMxC2uLJ81/TvW3zSUsXn6zjuvWTW/ZbXinrWlG5Vdwb1eWdmw/r4OPW8aFZmdbdXl9+4+tNHRYbt395G99NILNjs7Z8Njw8pr4YyztLBiQ2OjNj05afXKasmKYX/k6FFbXd6w8+cv2GefX7cTZ87Yo6k5u3broTW0dVo1hsvBnrV1tEll0tdLXbGm8UuTCMKeSAiB4KBcjoAfRTgLShmeC7lZqIs7e3qkOJFiuQFLrYzqO+y8pFilvpPrhRMimI80Raht1TRG8ZOo070ie4eZncvv216eLBzk+x6uPtAPhuhZa/wee+za2rqaGCh5la1XpsGV1p+pUZWRVl+v9YHvaRqHM5YUEQFz+X8DWJ9tVvBzwkQO8KqqtTY3yzYWvIWzHcourM14cc9ydBU6WBx7Amc5ag3WNBpT7j7gVsTCOpPe1CQ/TXsUdbsU0SXr6u4OKnzsvrHcDXgjxMeg4GLvZo/GNhnMBWU2z4x6VKYHwTWAjY/5EDnPsA6yPj5r8cRzo65zvOhLsqiewFeKit95XP6rD/Av7sDzvT3OuIaNWKmInSNwKzDU2ThYYPC7RUK6jATu+DFbX9sQ41kyrkrZbQBgFYXgVQVwU7xj+aAwTGegMvmZ9AIjQmGhZkMIaRaoSXMhNBz8EL+vBVWe3AkP/uLnFThEEVJiEQRwJTcDsNptMgCI8OKMgGgHXxLy4XN7Dgp5GBym32HBYOPjM8kyIvg0Cygo+WbKz8IEYIMWk1ne5Q06KHEYoMHhTRn3apQEMZlye47A+AA80EaPfUg9C2VawDeFNGAKoVgw05LkAEjGX9VCymIG8ETgIJ8pmfYcBq4Nz3wOucjxVdQLpA6BpUGZC8BLs8MZM+4/GzUNvPh3UITvqXmyD+PRmUVidSuzwBdUCg8KVDYsqR34txAGqWBcvYf70wJcAGTBgOT+y+IFmwYYewGM9U0mUuF40RG9RgS2aKEOxvaR57R7uXuRyX1zlUjRw3Sjjnk9GyxgZTooKqINH1C0KpCcN0N9wstjmwQ7FksfimIOWhS9nGMA2WBZw7rr7x8QS+CffvnL4BOd1sGbMZvNFQSSAXSqUSGPfs+AiVQrHiLp2SkU49HfXaEU+bM6u4Dr4bDBoQIGasRc4nd0r3SQonuf0ve4v/LilP1R60GAO9fH+8tWI3i/81z5TB4mR6PNn3PU8FPTCjA4AB88B+6xVYrWIKllxAqgMPPmDIU+r6lmCwVkYC4RFCw5KmsCcsl83tpa2myfA1ewJVIeCKHjQYkFEANowr0DrKXBJPZVjgP3l9krjEOKWwVyhVwNQiQl8wf8J8BO3vawenrlWSoJM1ZReJ7roFWTxQFs2/1cXn7FApFoSprZzt6uihkPt6t68FlggzH23MYhqH+Cx6QORvv5YKnldmnKRGlsdPujmomV7offrFQb4JisL/hGO0OE5kjywLrG56577+s+qhh0tRFrDUWXLIYam1QccVBnLfLn4b6/FGtiCsL8b27ROJK6p+DFJNciz9idbTtz9pwA0s+vXNEzi8YqF3/+7DkddlZXV1x5FjITYCzSDOOaAAyd7d6gdZYxlN3LqeErezXWXnJ+GhvU0GX9FBgbmtfMT8AQ7RWsywIcXD3hNXO9nTx1Sq9FMcqaDIAT2am5osMD32CvA+qyLvHsAE9paPA8xIZnvAc7JdbQaK1xwJgmjFvauC0GYyuh3AauLdXcrHUrAgKYk9zXiPEipYGYfRU9S147UvBxTxg/ysQp5N0PmiyRhkbtyxETSYcBclKCN2lkQ8U94/qYP5HqQ4HbfBYUX5AOsnva7xcWFu3b3/mOPX7yWIe7G1/cUgPdrR9YF6PC2RVYfDYF4nGgDqx6/q58DylzAKs8YykCLpxMQKC5g6+shfwuX3quKCqwPYIBrBBPb1ZGikjuLQBlS2urXhPAeG19Tesrz4dnGO3tYk1iAdDaIjYUqhw1CiE1cOiX7zSMcbevYvweOnTY1tc3dV+mpmfUFFUQKJ76IcgeEDxSz0SNRz6L21dhN8kYSrp1RGC2xWWjuG/nzp62kydPqIGN7QljfGVjXSxlmrOyfUPh0NsnwCRSrahBHFQcvIfnEXijPzpwcg+4VwD2HNS5TtZIxg3gqmd2+XoQMRp5tgqb39vT/Na9FoEAO4eE1G2vvPqK/eTv/s5ee/01O3LokP3mo4+09yh0uVYT+1I+6lhE6aCKT3ubGjvcM1eR0Xiq2MjQiN5LykmsFpDew2jWGC3IQofmCPcTsBT2PE3Fu/ceiG0P61Oe9VK6JgQQwwSffPJYKrZXX31FbHGerUgG5v7KrK3TU08luVfOAwzBmjd5C/t5PYe52aeWz5Vs/PCwba4v2YVzEzYy1G+XP/rIXrz0ku3t5uza1evW0d1th44ctqWVFcvvl5UvQqPs9dcvUjUqv8hicZuZWbDm9i414QFw8JRm3VetpzrXnx0HWHkhK7jX5zugkJonagpjM0CuEwrDbR/j5KJlyNLBVtFrKsYE+yVs5a2MgxGsI6wvrBuey0Kt5XuRs82dxBKpNNV8p6G3m3HP/nrCmd26AKIFY1vWEFW3fyPQnMO5N7SxI3O2M+UHfIXWNvannL3+4jlrTdVbMtUo4JTn15Bqtxuf3bDu7kGbmV20ZLJZzwxQCfKP1BnUPAq+pWFatemZWRsY6tdco1lAeDX1MfeSZvQXX9y0hiYUXJ45UMxl7cLZ09bZ3mKb6+QTQQSot5b2DiuWzX72i19qPIyNjspvn0aFmudTU1JULC8tqb6GdQp7vK+/X40TGgPkR8w+ndU9Zv0kZ2h4eERrLTUJYFoiXmfNjXF75cXz1tqINUnRmhIxZXUMjIxapb7RdrbzlivV7POrt6yEurTiHu48n+6ebu2JzCtADJRWrnjyecPa3d/XZ5NTMzY42K+9na+VlWWtZ1wXnwEgkdqLcUKWBGOM+yNf7GBTyDyieUKjglqNxhSvz/wolQt6zmqSxpysJZW0MnFiyNqtvlazrfUdG+lut2+8+oIz0vk5ZerUbPLprECsnZ1dO3zkqL381juWWVoRS3txYcFW1tcsVypaHiUQzetyRWN/sG9A44WGOnNIgBgkIUJ9Q4YNY1gNeZ0rJQvQl5QOamR4qDe1u+PYEDVQHAX1t8hF3uBX/VSjmefrFg0nlLTUPtH66IzmmJpeIt4A2EkdzN6MSo81NGbl/YIdGh2x3//+t21jfcUePbxn9+9O2XPPjSv3pFbzHIi/+D//1kbHuu2tt79m//W//LW9/c6Lun+E3YrJn9+3737vexoLH3/ymRUqFVtY2bA2fPwrVftP/+FP7MnDh7J+2iEHIN5gxaoTKbSvhubut7/5LWWtMCbYR9g/J05PSFEh+xD+h/Uen1nqKlcPslZS1/l5p2DjR4/puggDZo+gfqXh8emnlwNRByKdk/xUm4Uz5AsXLwrIheCCTVEErkESYJ/iZwEzxSLfLypIGOCS+lkhwVKRub0uf9C6gDVpyEVkz2Hs8uwcs6A55W4PYAx8RpEuY15/8vPUqWo0AXInff6wvrBuMr4iexjObLLBTSSsrSUtVwOeC9kQXe3tVilmrb5WtD/74+9bfS1vxdyetXV225P7T6SaPPPcaeEmm2vrwkYgVj1+Mmm9A3124vSEyAUQGxOtrbY6OWUFmhDkkXGtzSmdPZQt0Nkp4tQ+6s8yeU5x1eHcPwiX9ZAg21pl4UYzYXVl3Y4cHrdctmgPH09ZfVOTLa2tS5XTNzTkeSLUDZmMVKTYsUY1M+pEMjy5b1jjDQ8N2fipkzY7PWWrq+v2+ZWrej7MB54XuX3CJCCWqmZ0hwfqENX6nJ2bIHqEJii4CnUSlpMBG3L2AU2rejV2sOAEz5D4qcpSQ11Bg9HVleRS0NxhX2T8bK67JbDXQ05+8zo3q3MPigeAYayzyCSMwsGTTQmLlYv27jfftGo+Y/G6oqUa6wXM86E2NratqSlhW5sbNn78mNT4sjCbnZeibnpqRoHyVz67YicnTti1azft0ksXbXlxzcZOHLfV+VmLN6HiXxPhraWtyxbnV+zChefto08+t4svvWQPJ5/a3SdPLd7cYbVYg21BvmtJK1idLC+de4N9kmwMQ14La4/sreu/VN6yDgJ6s1+R1Udu09ihMVvfoAZqUe1D03twcEDKEm4m2ZiydyuXhGP09XZLAUVNTP1RV63YQE+n8inIp1pfy1hra8q2d/Nal0t1pnqIRoUyzERmcpILWRmMDSka8nmtPzQKlQ+TdjzsgJRZqRzUv9EaES3qke3RvwRuI9ujZ/+d11OtQWYoZ9p0iwiGrHE0SFnDGA+MVSxVozoCIhQEXC5YZE7qJwhA+ZzGC8pCKXubIMi644KTJqp6RpxX3aEgYZ0dndrH2Xu0fkldwns1qIaGKMQ+PTwyrHMe6xPnVUg0PD81TMiYjXAknrXWR5qnkYLM1c4RVqfmxFeKiq+w/f8/34GJlrQtL69Zb3eHzc8vWl9/bwCoPAj00NiYJiWAAYcf/kuuAD6IML7cWskLaQpGLw7xsHYLCSZ7GdAtyNz5nsCaoGDQQUpMagAS5LReILCSsmiwcEcB1ALnAoveGTYOFFGgRkWFii0pAhqlAAFcQMrGwVxyLLIraiwwMOibbGN9y8EiWKHBCkXBO8GjmgWO15M1T9hceS8YmACIkZKAglfWQygwFAZIIZQUyAfgxubO4Z5DszPe/QDO5+fwxIIVBU0lwuKWRHFShoVL48VDDsXeDYxXpIUwx4Gt2RRkOxR8NdUp1730gGQFnMr6yaVxDkQ5u5XPJRZjkAjyLPncsNoo4lmlud902JVdwaFXr++WDQLS3afJbRx0iIDxHUCt8PPO+Aumg5HMLyyyDji6oiAqJHnlZzvH/p7+5YcUZ/ry1u6/7Wx//V2ScA7pfFAvRpGWkosg9mtdnaxDdDgJId/enHN/1lKxIACGTYjMFA4o3CYKXoAzOuhq7tRqajKxIQMoLK8sO6Mhs2ub21vu4YoNWsgHwQ6H7wGkOisIOWzJWbSyb3Hv6IhNLlVIYItEGxWvpcMrG2vwf5fFSrA+cWaSYiC0OSpoMwQ9cR8EdmV2wmENcg7e3TndI93bAA4p8Jjr5jmGcFnPOsFDsmK4PuFdLBULFiCA3fUxfT6BIYBXFfzLOQS5DNUbXDUfL+qGuBUG4atInXkf5khzq9uKuCLIrVvkdy45rLO9GdtqdOGnCVjV1ORWMbGYQFeKLULNKXTlyV4sKnCuWaBe0dY3N6UQM7Er4haDes69o1laKFq6EQZWWqBuAiVKS6usHijGKQw5LBBky/Pn93lPfpZDf2TbxdqicLAqDHGXxkf2cBQ6XDOWO7B1pBCDnSj7EA8yln0TczNkqyhEUCzFtAp0njVFF58xAhMp5GHbqBnJOtSEggtJK0CXB+oxVmSTFOx8+DysEbKTqplAQcJF+TwEuyGdhtVO40R2e7ISw8ecPQCQgX+nEPUMAv7OAZggPIAT5iuSb/fediUAayprM6xrgBPurR+CYOa7NNfXPfemlmevFFY0h8k08PntIPq+hwXv7wdmiyuSVOjCSisWrYTtVbAB0BhRAG1FtjgAsMxh2MPMTeaalE8lD6lTEz6oFNQ0kRIA2ysPd2S9c3s3ABD3i+dZMZ+R6XOvBEY+o/ZTYc1Ph7wRPhMFvGyOlDsT0/05YMzAGOW+FQo6eHkD34FIQClulhraUQ5JYBhpddefIwsuX0O5Ro0FqdB8HdKYCfvcs02hSJ2oewYjXLk6/v4cdGDS0yyLDoxqHEvV5ewgHxdNB819WT3q2bnFFfOMGoG1J2q2yUYStRx7V1DV8XuM4cjS0a32vrQHomZQ+GBTUsxGAbaJuNjjfAYOgYMDAwIXT52aEKP58eMnsl7EJiqR8Ea3Wwc5U5TP4TaGkdLQw/kAWfAF5zNyMOKw480uB4HOnJmws2fPaAxjFUPdA4jRkExpLeO1yVNgzNJYZdwAbvjBB0yKccdnd4IHY1Cvj+Rf1kox1Q6RopPrZr+p1qFAKGmuRfuEW5w4Qzaqz3hGsIcBcmADb2xs2csvXZLyAxXa22+/ZTdvfqG5IasY2TS4DSigBM+TfUSWiAQWhswuzRXmWamsewnoCLuQz0ejJLI9YiyhbmLthCUK84zPCghBYDw+y/xSe0e7116qD6qy0KL59cZrr2m90PiO+/ivq0+oUfPo/kMx4BlTzeRtbG7a6iosTOrFssCUN159TfYG165+aodH+q2vp9s+/vXH+twcFv/+J/8ga57e/l7twWsbO/Z0dsEq1aKNjg7YoUOjBhN+Feun9W3bL8EYTWlMYE2XbnZbE9RLKMyiZ8G4UogjTURY7ME/3W343E40UlCxJkWEEsas3zsHBWXvRI0E2BopR6kjgnozUkLxvjwH9hDGhZS7sm1w72b2Cq5VTbxghca4jA7DzalW1ZDsY8xZZao0JgUoSe2pbbNkTU31tr21Ym++8pz1dKRwSlQNyvVldwt25fMvLJnCQ74mK6Sp6Vnr7e9R7QtIBnNfIfB1cduUd7k3ZCJFLc9e/s5Y/iXiNj+/YHWxhCUavMFVKRYsVi3auTMTap7IEiORsPbObjSf9uFvPtEz6B8YUKNiaAhLpJgtLS7ZxMRpe/LkicAMxvqjx4/s8JEjqoFpkpw8ccKe/N/svfdz5Fd25XmRANIAyIT3rgCUZxVZLMOiqWbTdLO90YxampEiNPvD7p+2ihlNS9pZ9YxGpkV20xfLW6C8QcG7BJCZyEQic+Nz7nsgpZj9A6aDiGCwqgBk5vf7fe++e88995yHD4MBd6fM35m4gCUOA1Xa4c0NkoW58PopG+xus631RUs20oAhj0pYa67b6k0ZW1jZtN9/8oVt7+zZ5OEjtrCwoHXAmUte4jnlpuXa2rW/XMYLQpZPCC0tL/nPBoCOeMHehJAiTznlj+SUZevBG6WAGT0NWm+sylNXBtNOGgIMpbbwZlnVdiquGy5VDNVz5Fth2pO6rOTTtXh5DXbk7PzJl+SFsLS8ap09Xdbe1amzhue+srSi+/nS6TNW2dwSe/zWzVtWAGgt79h6Ycf2+MzyIEIWqOqycazxpoSmYBONELa82R3zIendh+kfFoWk4gKfn/0dPfmYYqLZybnCOexeO56PI2vE+ucs11lGfgo7trNLRI8oJcjPUsNyjyBcceZ7g8KljJimQDKGdQmI/f67bymepjNJu3ntinV3dkjObGFxzV49/Yr95f/91zY8MmAf/OBd+8f/+Y92+MhBrSPWs2Tatrft5z//hRpBn391xQrlshjxuWyH8oi/+I9/ajN3p+3S5Su2XSpbjXsTpruV+4uP3mA/+MEP7OIXX2gymYYjfgZTU5N26fJlz+uR3MKjQhJfPk3hcHAgGaqurtiRQ0eUS7MnqJ+5n6dPn7KPPvrIZXHFfg7eV7xmkKF89dVXlT8OjYxIGkfyiKFejMREal4ZorMeGxsFMFd2maZwKWKxngOhK040qnSg7mUaRLW8SySxXgFDqT+oF0ReUB7swJ4mliXV7NcZZYCdlBBkw8IqovbgBakZ+rq7rK+vW42j1bUN62zP2vZG3hr2duz//E8/s/rutlWKW9ae7bCrV2/Z4vKa/fCn39c10KjoxIcmv2nT9+7ZwNCgTRyc0hriySqceAAAIABJREFUmWQActfWrVwse0N/Z0dS1Bi8K78X9lAWsQpJKe4T9RHnQk9frwzos12d9uTpM2tuTmlagTOkWm2wm7en1QDMdnVbgUZqKqMaDSyEpivAqwgcEGvI1yRnhvxoKUzL+oQKd6u7p1cTFcjOwQwH/4Dw5Sx4Z6bzRa4kHyQpQCBHlwvkTScjKP8Nvqexec52pFHBlAdMfDXrG3ierqIhecKEExyGBnuVlwM+w4SnGRLVMCJBRSShRIP19fcp3+OcxacGEL5UroiUK++k6q4mKrbXFi3TVLeOtozlWsmvaraxmdf+3ykVNDmHhO1Af6/NvpgTsYBpvskjR+3Gxct28PCU/f6TK/bWm6/ag/uz8qpYXlmwZIam/4aIqunWnK0srNqB8Sn77Ydf2vkL5+zJ7KI9eL5glm4zawKvAhdoto21Nevu7rLt4pY1JprVROAhEHOdzIOiAdKfAPJOFCQuMpXP7gWb4EzBZB0pLXAM9gKkioHBAXv48GFoAkVcqWq5XJvl2lu96V6tGR6ZPNH+7pxlmhKWbcnY0OCQYvyL+SXbwdePvVeray2yv9RUb066t9Wa+zZCauHf+bwtbZ7fiXgnHzaXfmOPUgNKxk+eY+4f6LWpkzD/V1+xMRHzFM+ZnezE9/p6etz7rrlZjUFhj8WiS4MJP6nJexGfNRp2q8vLwg0hAHhOBsm0LkUY1djUPVGSSY2XFj0D4g75KnGUHIqzh9fnvnAvUIFgT8XcCuUKro3nggwlsqBSSKhWVe+hMvDg0UPVLCLxSK7bpVAVFyUFxzS543DR2yLeo28nKv5/l8y33/jf9Q683Nku4IPg66NOsKqS2rBxdC7q8ZPw4k8RWYawBEmoOcgIcHzBzPVx3AaXZiDhDWa/sVnh0wFeRItJHhinAqoyfngKLFZx7Zs0JhPOEPOilUCnJERsDqfV8POMY2VaWsU0EjM20bSvgQnQj3yLM8vc14CDjaRAAPceEhFZJTIux9SgxJkRQIIXACv3K4InjAMzUoimaU9Plw5lgpVkSgIYDiDkIHCE2d3LAQYTSTMdVox+SYQl0wMzO58XiwO9Sq5HYFXwDiAVjaa6JLX8XpyCcakdxvJJwHf0ZxkPCihnXNAPAW6Ag2aePHLfkAHhM+owpNjRaKePCEeWpG5c3RnDMoLU69Qlt+NmfDyFYEiGDI/MuX06QtJRjAmTPAYwnUTjm19ivUu+w42CIkgXE0kHYynGnAkQteM9eXW5HUZDSWr8d4OZsYBGN+mTXjwXIaDIgXd+n/XpmukmJgXgMcV9d2e30XXnsONCSGLofo+MjtnUwSmtNYrth48eW1dPt63nN8Te4N+kw6nxah8xd+DBJTc4IDnAfWzZZZMAaTm8JbsTmEnxHvAz0nYM8ibcE58ycsabAMowDeVFPUC1a7hLiiIwykjwKL73p1NkQu+MZm/0eQPGD2HYRy6poRFqklAOS7TC00k3kGxpszImqBSzSVgo60r3aVBEg16NdIfXR+MaJIFnIKADeQEYazs7SoZ4xjQqYHwAvOW3NqXdzn7c2trcZwhHvw3JLUknGz+ODhmwApKT0I4MD0kuBbCNAx0GZ9/AoCRHKGg2C9vWEHw0YJZyH1KwQtIZSyYabWhg0Gbu3bMEjSWKHCWLziAjRko7N6whiiwASAD7fbBTU0cuZ0URpYaU1qkz3/iCZctewhS6syOnYo0xfsnJAZgHpja/F4Ff9Fm5H7BMYbq6dJTTjrQWNAXljL99iSo8BNqcbURiCyAfDXUF6ofwBFiTz8Pgh+lZs/HRESVGMCRh0HsjzPWdmSyiwNbUE5MigcUNwA/oCtuGhI59I6+f7YLek7MknXKTV66FRpkk2mD2Bt8f/BpY35ID1GSWA95ivdMUaHQXGO4/MRmGCskuay0aRlM4qSEifdKqJltio0XJaKUioCYd5BLwWJBRePR7aaiL7ULCzXvDBCcZ5rOQZA4PDdmN6zdsYyOvvc3eZ1/jYSTpkd1df0ZKQBe1NjhrYryOzWo12mXu6XGLfxcLKUwouH8AUhwwID1mRjmv/fgZppc8lnjTjftGqi8px+Cl49NqDdYJ04wJl8K2vZjza3RzauRfvCHmjWWfdgPkddkYn3DyRB7AmkYkxpOeRCvGhrivIiGA44AHKjzZr8QnmNhqvJQ1DSeZIWSFNJ3hwLcY4sgvQJSo7wl0BmwHvAYg9EkJnzQkdlIY8POwmCgwWA8YAbuRM5NkRYH93OOx8Qmxpq9fvylAc20Vxh3x11mZPDtps8sbAdamF/L8WVIXrMNdl4za3twUe9DZ5QmNhyPlcu7sGd3fzc28Jj02NgsanycPYX9yduODICPfvbpkmFxCzjSaD7uyoclPKPYR01yaKCm5PAX3hdwhympG9prTB4I5epA/UT4VWLdxzfBMW1ivpYLOw+HhITt79pz9zd/82g4dOmyJRiDWBhkHSz4rS2OkGHKlqoBcgA/A0jhpybOExQggwJplvRYrNNe8iM319NpuoSCm99Wr17UXurt6BCTyGXm+qxurNjE1IeCD15YhJ9J9Gr8X98BOnjyp54zhM0x89hxg9ybNg5VlgWS8HsbAExNjduvmTek7a6KjWLT3333PWtLNdvvWVevpbLPJ8TH78Le/twtvvSFv9EtXrtvg8LCKWQChxsaU3Xv4yHYrJevr65RnAgDSwwdPbWVt0za3S9bSlpOso6ZBdf7G6VXPZ/QVJJrYNzvFknvpINUkFrCfvz6p7FrskfErxjRN7AZn9XE/KjR2OtoFnLAGdL6E/FivFwggIgKhOR+a22r4BfNJTaC2ZELsxrvLpcjUdGzE6wBtanJzWPdImfLZUMnwPBGgtrCdt1wWhnLFfvS9t4w/sna3tzct19lppVLVrl66Yel0zsC3kGMCmElmmNas2MrKuvUP9GvKEcknznPJvbV7fQIpACYrUpSSekviZwSInbRCAa+SnG1urFmuJW3jo0MyMCZPYRd0dvdardZoH374O8UvpJ9g9iOVQnzEY4JGBZMV3GsmKu5O37WxsXFN3wG6MFFBvUMTjXMGZubk5JTWpsgsApIS1pnL2GunT1htZ9P6+9ptd2cLFNC6+/oNRZPdepNtFit28dJ1q9SbrLd/UKxzziRIGlHyBmbx0OCwvUBuSjkcchrLqk14v7Gx0QCYJ8XI5FkCeKyuMiHWos/oEm4uL0mM+uT3n4pV72uQJgSkngbJWkFAQ04l05axtfy6CE+cNexZ5dRMwtGohcwQJiqI0wmMukeGbH5uQU2spiTN0LJ1duXE5O3MZa2ns9MGB4asXCjYi+ez9vzZnID/Ev47NADzeWuiAVCpaJ+lMilNJTVnPOcq77ikMLGYNc3knhu6m5NZ1KBEgsiZ8sWdgiawaE5QT6TTMHg9TsuzjtdJJTU5RL1JTg1QxtlP8yLb2iJmrM7P5qTNzc9rvVZrTAC4DBQxzpmybjROHox8Wntbm516+Zhdu3LF3nrrnGIEhIp7M/ft8ZNZO3r0kP3mN39v3d099pOffaBGHoD11atXbWbmiWW1h8x+8uOf2OLCin351RUZZc8trckYlnjyZ7/6Y7t3965dvXbdCuWq7VI3BMASzX41IBqb7I033rB709Na3+QsxKrDhw/bl19d1HkouVk8fWgKhfpSOXlDkFRS7m82NjKqM/Pho4eB2NVsZ8+dsX/58ENl8C7P589Bjf3QdDh29Jj2MDXRbPB/UQ0bJsAFLDJVEUC8fWmnZsiBLvvJfogLlp8FEOeZRJCSNc4UkBNfkDHs2K8bpURQxqvGBD5Sh0c5Q/aE+zA5ZkCe4RK9Hq95PYH3NI2RdOvq0KQH+6KtJWPrKwtW3y3Z//Wffml75S0rbq6rsXjjxh2bfbFgP/zpB/KvK+W3JBmLmTZSpF29PXbo6BGtS2I/BC0koKjxWY8un42fV6vyIOp79irNvjt3ZzRBRz5CrkbujERssiUtPx+kofBpY6qiVsezoGC77PNUyjZLJesfGLYHjx7pWjmzh4eG7dbt2/t5PHkycQ3iCv4i5L1zLxZsbHzELlz4jl27fsOu37wVWPI7IlRF6SfqS84CyWkzURGkO1vSgNNOWFAqGfAc9q1yX+EO/AepzmtYzm+a1YITmKqW9JNGa+RRIRIkqg2BqEfeAuirxmxvr3IpEZZEBNixnq5uSdAtr6zpvhPrOLOSCbN33jpvc0/v2+hAtyVqdetsTyM2ZdUquW3V2nNtql3YK8TSezPPbWpqRPEOn5Y7t+7Iu+KLLy/bG2+elyTUkSMHbXb2qXX1dmuygCmkLjyZNgo2PDRuH39y0V4+e9ruPX5mD2eXLJHJWmm37j6JLRlbW15WHraeX9P+JGZT67BGqCk436khnGTpzQvW9jP2mM67LknMcY4xVcrZQS5fLO5YT0+3Gu40kTTBSE6BIkoL5tCdaubw+vmNLevv7bQsvjvNjdZQq9nkxIRNzzzUOqsjcQluIXJFQuRN8D72EqA/06BqRDBFQYOc6fVMRvU7azhOeUK4os4jH+F1Y9OB9eR7NJBRAy4R9+X/atIixgTWIOsI2U0IS9wzYgb5NGcnE5ysFdVINDwb6tbf22/zmmLM7TcIhIXVmERvUe3IfmPyPsob67OIdJdUrRtJlRCeaLap8RvWeKz5iS2sS/YgwQaZTu4RcQsJaKR9UfDgPJC6RWhQ+BQ5fngufUgtET1GXMEvYovfSj/9K0Dx27/8YdyBgykv4E+cOKFRP0xJ2eRsBgrgjfV1HZI+IdGgcbqHjx/bnVu3FZhcz9KlDpD5oKPP5AAFNIkqRdSOOtPeUYyAOyAf4B1fHGx0fvk+oL3AwiBRo40e2BLO2nCAWqwwGT87Q9nNlly2hqKGAM6BtZEvWi6LLq2DAQQu9CJ5TZLw+XmSf9dV5u8KDLW6GgboDnNNFHEU54C/aD0/n52VUVJz0sf3SeLdk8OZneqsIuPU7qAKn0/gpQCeMOoq0NkDM8UTSRBJMMmoOqWScCntT6t4QsVn80RKElTb2wJLYRV6Y8EZ8G7UCyvUpMdNkRnlcDRVEZJ1klWCLAcJyYSMzMQMc1YrYBKJIUAFRQTsS02M7NKBz9kWo+IwgFtaBNr4qJs3Jjho1AQJI8YEZRndheYIkxpiNgU2Cwmh5LZCMc/1cDBTVOigFSvaD5fYWPEd6E0Gmbmr2QAT0GWnSK61LltSWhuM8OnOwUCmUEH3GG3rwP5U4oyOLb50GH+2ZZXQA6TSfGKPYAqHJBSmZtn2rADc7W0AVYqotFguTFLIlAq9WMzYgqYuhyXXCMAGEO9MILR4G+zFC6RnMF9CmqlRz0KMrlAc6jX2TZ28URcBR4GacZoiACGSPJExs+vjwwjgi0KXvcxBp/0XJlgceHZpM/Y0hzssY9aXZEHSae1N9C2lm727Z525VnkEsIbYlzRYWP802VxKyYE99iJ7iGdAgsozKKpZ6QVVI9NAhZKYbCdeekmFDCOsrC/2N9fOf8i+CAgP3idqVAZJrChHAzO0q6ND8gKAauiQqzkmqaiiS60MDKqo4dkBtPGJiAnod5JUIplV2MjLuHB0GGO0RU1U1DGADzrH7HsAggMHxu3Jk6cCHnk/fpbmFoljTKb26lVdszcn0XhtFSioPRpGSQGaAAOfPJu1VKpJjEL33PGGheRCFO9osHmTFSksEieR2pA6wIydRqskzpyhBuDEJBFjvwA83FuePUkXQCzPhGcv9kqYsuK5wJqikcP6xRAYaZy2bLviZn4DlpBLMxHrKZpojPBsXDKubEcOH5I297PnT2XkKtAtNGaUbFVJjtsEBMX9TKGY60DCz9cq65QkkTF1MU5g4ygG0eAu6h7QeIVBT1zlGgRWClBuUNyLbFT2Jixd5IbU+IahGpJM1jaasDr3NFVQV/OIMWmavRQ2/A7JJdfn0gquvUtzTVJsxDz2kEBKPEnY6858EugNGNja6nsAwFisG5d0iswjQDD2F0xeQDnW68WLF6VHzr7k7yTh6F2zdnmOPAfWk9hfTLUgsRe8m7jnADpoH3OfuH8yv8TXIZNRc4vnS7LOGRSJBaxl9gx7in0iEFX6yb5WJFUSGqycvpIOkcSVn0F8RTNsl42q6XNKHkRNpIRkCxW3qoDZNSXssA45pyNDDuIC+4bziQYoMQTQkJjBeabGVJBy4jOSa7AOiFtIpEhDVkwnZ1UK6MJ4WRrWPg2J3wBsQT5DfhMWN7IIkC68ec/1RtNi3sNl9pyRKa+kJgCBTevt6lKzgvOCCSQAB+Tczr9+3q5cdtNRni9gdt18KhGmPa8tc+NyWTrxnLEA3L53yalo7lT0HiMjI3bs2FFdsyZvMhlbmF+UnEVsIHG2aIILk+5QPOrvNGyamDDrlbkqf6epqwYf8ai+p31KTHr//felU889RJuc6SjALrSaaRrTbPApRlhySCtt636g28+EGa8rqYRchxo0MMOSGZdi5N6TC/WPjNizhw9lsIvMTbIppf165NBh7bHd+q51dGalbx5l2ADK2DNMeq2urNjrb71ly4sLdvvGTU1tJZpTOt+YWkGigiJ9Y7NoA/3d8rVguo41UNjCb6NVYEdbC7lf0d58/YytLS/apYtf2fvvfaApt8++uGR9A/0i56ysr1lHV689wwhxY9POnj1ujx89siOHj+jsXlnNmyWSahwAirhXDQQSn3hyw1embmlSk/e6ZKbiHOcnhtGbNMrJQV3Kki+eK413ZFejaS151kZ+U1MlKT4/TG/5tnkzk9dbXFrSOag8ir2BVEZ1T8U6/0bzjLjN59kU69NlRCmw0cSmoKdhgbmvT9u6PBiApKZgkBptcgIM7NSmBF4VTBqZJipyLeyTPWvJtclLZadYtenph5ZOw+5slJcHwAmxh8+azXVon2KqzPUQm5BZybV3KCfifsCQVZOHfZxJ2d3pGUlPpNItNjV1UNI7GyuLNjTcbwN9PdpzSxhk5tqtra3DPvv0C9UkAPr4UfDaxCPW39Ejx6Tlz5kDg/bWnTt2YOKAfLsAW8n90Nnn+8Qo4jTvSSNBDWQIQc0Ja0s32vvvvmkDna32cOamjQ732erykpplHT39VrWkPV9YtX/6549tq7RrQ2PjOpuJP4cPHdQaIO7SZCPXpxbyPYNnyI7WOZ4aI8MjWlc8d4B0rmNgoF8/5xrjPmVQq+3KA4bz5P/9b79RLSeT2UBuYq8hDURdNDY+Zktrq/LsQsqwNZvV3madCOAJ0kiaPAgkpFaA4nxeZurjBw7Y8vKiDQ302+LCC0vUG61Wqdjxw5NiL7cz1V7es6ZEWszsaqLBXn/3u3b3wUO7dvOW0hpqpqW1das11OgGaDqpsaEp+C54DUAui2wN8X19A4PSIP0TJP5kQltDJoiz3OSXk860ivnNPYv+TxHYog4rl8l1vSGNrxk1D/l/JAeQh6I/A9vfpyldcnVXjX0+aoM1J8xGhwftrddfs//yn/9KUxXHj0/ahbfessZkynaKZZmk/9Wv/6dNjPfau+++JbY4kjLkG0z2Xb1yy2q1hP3qV7+05aVV+/ziZStWKra0XrKhgS6RSf7iz/9MMe/Slau2DWHAGq3a0ChCTKmwrekXzqG3375gt27eVt7MF82XQ4cP2ZcXL+reseZ4pprwUv3kpAT+E+sZ6aRS2Y4cnFJtMj0zrVqIZvCJl0/YF59/Lrk92PDKzcKECzGB9z84NbXPomefEMeJbzSFykgZJmER+5Qi4GX02UM2FxISuYwkyGpIHbvfBOegk1UcjHSJTZepjMQO8jcHRbcUfx3cjI0Pl3jxGtd9DCTJF/Iw5ZnhZzWVo2mmioBcUm+8dsaHB61c3LDezoz90U/fs0pxwwr5NWvPdtrMzENbXF6xc6+fEymIOqJzcMiKq6v2/Pms9Q31W3tfv22vrWvPtqRS9ujeA10H01LcfkDPrc288h78ePBUYC0jQ0PcpvYil5w8NOU+adTSjUwM5TT1QWPv8aNn1pyGlLlnNSZpw9Qhkk7PXyxYf2+XGv1Xrl7V2fXqKyc01fblxS91nUwV3puZ0Tnb2dllL508qTP1xo2beoaq34KcMRNtml4RyQiylJNGWVuaiJb/oE+HS4ItTJUr/1ODPmnZbMYyLWnFGa4Trw0wFpH6mNRlfL8OPtSuCT5ej30NUFwI9QX5MdM7IniJeFfT5Ei2tU2f6/ncoprtrCcalLvFbXvj7Kv2+P5dmxwdtIbqno2P9lmlvGlb2yVra3F1Bhpt2/kN1dJgQp1dPfb4wUM7ffpVm55+YCdOHLUvvrhob7/zXXv44KFNHpy0O7dvWW9vt34emanOzl4rblds4sAh++ryNTt26pTduHPP7jx8Zrm+QSuU92y7hGxTv+SiOjpytra+qtyQupvajGYF95Zr5oznXOdsFrbT1CwiFOcb646aFK8l9h0EAHJE8kYm8e7cvav8nP3eyDSMpk7TxqNbW9+0zq521Z7IJmdb0raDssZuxc6cPq0pyJW1vLxPKpqo8EajyL3RyzN4VUYSFs9QZDmkz9MZn+Tf21NdA3Et4kbkhcQh1ot8lFQDpvbVMyC2COcKk9/fnKRwQpVjgSKIVXatI5B6mHYktwZb47wQNhXB/Ya6CDI8Z/JD4sDayqrel7Nfk4SQXBudpOWKG437ai08C6a6kCbUlFZjo3ItCEURywKD0v4NPpNOssWrF0UEl7Em3hF7yK27e3v3cS5iGFiQaqqgIBFJ2pEoFifaIiL97URFvBPf/v8P5g683NWpTh6JLBsxyk5Q1NBdZ7PxvcjIfPjokbQWKbJh/5EIcGhQjAK4AjZIMqZeV9B0YzPfhOpghjFDaUjTKQ/a1GL4BkAOJC72B10v07XvfNTT5W6i/q6ztKVtEQz+XDaHn2fcH6NHknGSdxJMsSODvwJgkrqfFW8MAOT5aB0MzMAmJzABUAKac+g3wFJ1c1MOCLHhoxlq0OGX8U2C4N+mg5drUcGP3ErBzamkj6dDBnaPvy+HhxiwyOds5JUs0mkleaaR4Sx5b9aoWRGmInyIgRFML07Uca86q1XMGQyCZbTrUwUkX2KKJpGpctkUfleMFYppFTgkrzQqguQCDFKaCZo6QOsbJjnNDNe8VwMpsCc5aOQdEBI9sbvDFweUJhpCQ0LsCAH5bpj3zWvUeLIAemcRx9G7mKSKLRj09vk9TQHIbNiZwN7x9kkZAU8AuYCRMn/z+87X5samJTDDhtEhc1Y3ouZ6MXZnqoX3J0EEIKXQo0BubGoQIMF4ZqalTU0sRtUxDKsnEvYcLd5FgGRnurOuJHFTwOhzV+wz9gVrmWJV2vVhokRFRJBFi82ZeA8d4PPEex8MDyAu90wAJcwqGTJ5ocr7yCwYPdpmZ+KSvMQRee4LSZE0f0OzgvVKMgjADPCkdQeDWgbXdTFxGf+PDUS+L2k1JS9IfLjsDr8v+QkOap5TA/cPk2HXpt8pFi0LGzmw5rQeEkztfP2c+F2ZfMKOkN6jexnEKRhnfzZaLtcqQI19KW8OmeNWfGKhUFTiNjFxwErFHU1Z5LeKlmlN6/UAcWAz8ey7cu37xeqDJ8+0flo72m0dFl7aDXABDiiYiXlu4pqyubl5FVgA+gLw8BjAMLSKhjWTASkBzg461cXiIzYBDh89ctju3b/v+rx4R4TpJp63GIHS+PS9AlNcsULTNQ1iILIHSJKGBgZcW1z+He7lILCJtdqEnvoTxYvtAkaT7kEAGEQzlpFzV4fy/cNnhqXEWDmTMIyHuyHyjjOgg9QITSo1DwSuuSEkUy2zs8+1DkhGPc5585P7L4moIAOlxJtETM0Wl62KXgIe7wIDKPgesOacQVzWtAINdMnSUTBxf8TI9wYnz0GFNw0Zg2XnDH7iFOC3JnHamcTptMX5BV0DzBYmg2g8Lq0seZM1TDnwZyXNgd3iY8TOtJf0GNeH3nAT9zXlBpJpJAmYxFpzZqcMBl3aiF9W8hw8iOJ+5/mxZ9WUpDCoMKXhRrmS32HiQY1+9xSJsZL1znompkuTmBit+4I5YknnPID/+ddfV7Pj+eyLICGGFAxG0y5ryPkgECOMmwsgDMbeLuHlZs4OYrqkXJz6omGhJjommM1uBscX1875Q8OOWKBzFNZrKiWQmwuK55q8NpoaVVzwfGngaqqT5nGKQmJDbDMao7yHDNdbW8Xu8mlLB4rJaWC1erHg0irE31QyrbWKnBn3sVCgIYW0gkvzcb0OksAGcwlIPiD5BfeH+Mgao5BmH5cKRYH+xBAeJ/fuHYrXhw9sbn5OhoovXiza2kZeLHVej2tisohcwmM+Jsx+Vkhej1hryCHldB8ASVlL7rfgppUy3KXoCdJKxBvOBxo5/CzNTK6ZHETkAOVmsLauOSDEBC0yk8HzhubrSyeOW44JG/a0PpuzIqt4TTT6pBcx5c7dacvn191/qbtHE7Y9XV2KtYcPHvLnzr6p19wMvrtH+SBrEzPtQweP2PTdu2IoypesWhUj8DvfvWDJlGunAwpTvD188EDxdXBgQPutOeWNiWf4i0AIcDU6yco8m53VtX/wox9qXUzfuaPPT/ENu5dzY2cbv5acpVMJe+P8GZt7/tw+/+SS/eQnP9TE1hdfXRHw0d7ZaU9nnwuUo7BeWVm0kZEByYEsL65I5391fRv9Givv7ql4J+eiaS55ETUOv86BiGcUwG48X5Ksjcc9z42UCzIJ0trq5Jayr1lvXnwtM8feouFMs5f9T6ymuQfIKg8MySh4k5CcnM+hpljFCSnkxUg6ET9iDppqRsKtbLUqzQ9fY9lsu2Ij0xFcE5dCzoz8q/I1PJiKmygoWmNiz86eOmQHxgclh0K8hVG8PL9iN67ftbZst+1W6pbGOFtm8EyFeqEP4WariEdD0mU6Sjvay3xWQAMaFTSGIa6o6dWctKVVZNJ8UgSwuLsjK+JRgg+ZwDC0JFPng1MqWr2FAAAgAElEQVSH7crVa7pmchqYrkxW8MV06eHDR7XOyC/Q+L59967qHhpzxBf8VJ4CemWzIgjcu3ffjhw5IjIXOuDclLa2tLWmGu344XEb6euQmfbO9oakXAD19hqaLZFstbXNHfvi4lUr1xo1gUO8JWazt/GNIF/lzHJvOwc5iG/oW3O+M1lBM8UnwhNqVDjI4Y1cPh9riAlR5IeYBhkaHrG/+Zu/tc7Obm9Yq35rF6sbYFS5M0A9HoPyvOLZ+ORznPBjfWlaO0yQAjK2ZtLWhPQFeTEyGvL5Qha0wWjVtRJbmD4lrrGm063WmeuxlfUNayCXa2uzVFubTT94IFmW1hwG7zXb2ilqHyvL3a3LWFjxLvgGQDpy76KaJudU80AAkIQGE7uhZtBUoKkRpkaFojN1EnWdn6nkHUyAuhxQg6ZpaWISL3g2Pi3ouRN7272EQo1B07sR+VKaF2bDgwN29vTL9g9//98lJ1zYKtjPfvZ9TV1n2rrknfJf/+rvbHS0244cmRQT+4//+GfW0dml+3/3/kN7cHfGXn/9DXvy6KndvjujiYpVycIkLZNM2Z/8uz+yG1ev2vWbt61UqVqNuJloVn6DBBsHCK/1wx/8wH7723/ROiAOIAkzMTUpbxfum6oiRltYnQLKnDRF/e11MDJAZTt+5LDWB7WMiEWNCRsZGxPjnrPQSWkh14iN1waf4uF84rkhV4aMCsQ5an15KlF3JlwqmhjGs3GJTeJYYV8G1+sRJ7Fx7kr+LkjC8m/44LgiAP4NLWr6MHkjHzBNpbkigJvaUkP72ojegFH6WDBnAB4iDsDUQHdnzlJMziQabWFhUWbw5cKmmpJ/8R9+bJXShpW2Nizb2m7TM/cF9p47f9Yy2VZbm1sQo39+fsFm7t9Xc+HAoUNWwjcJgkY6bQuzczI6JraQg5PfADbzf64FWVfOHa5Bnhvk7sWi8IW+wUFr7+5SM4J8S7l7vdEePHgiQkQVhjuyUStrsPjka7KwuGJHjxy0iYlJ++TTzzR5fubsaU3P3bx1WwS3N99808B6SkWmk4ghR9Sg+vCj32n9kz+xB4klnBOSeoPg14i/ZvArUBOLhhD5vysBxHpdRRZ/F6ZDXVqXRwVS2cgu1mtB0oZoojwZMtWu9XR36tlzbnK9nHVgTyLUQI5TM4umQtK6ICZg2t4MiXLHdiq7ts7kayajWoUhjdMnj9ujmTs2Nthn1Z1de+noAauU1q1UAoAuKfcZHBoRltTZmZUsT09/v22urNnkoSN28bPLdujImH38yU37wfdfl1fIsRNH7eG9Gevp67a5F/MydW5qbLXtLRQDhu3KtTv26hvn7fbMQ7ty54H1DI+pUUF9hU/X1saGdXV3ak+Qu7IuqBeUG+65TBmAP80L7iPxGfWBF3PzWhM8R0i5NNdpTDFZoYn4rW2bOHBA6xATRCZFpX5BLdWC/wL7nrwDqV6ICE1WYYo11ahGBZKJC/PLtr2zK2WBje0tkWWooeRZyBRUyN+JCxFDkycpShFqoue1x31deNNYOYsmxjlvXHKQHFhT9GEPE0ui9DU5ZcQ/iB3fbFi4UpTLjvX3IPloVtx2X8CIAwo3CXKZkHGZXsHzTBO7aRpmGTXqHfOkDub+4k3qeJGkvITT4SFZUtJJbiXpJmTJ5HkLKTuhJj/7HyIX5xLvEZtEIg3XXdotTp18U66YmoAveT4qNnlwUl4X7hN//1rJxBGibxsVfh++/foDugMfHD+ukWMHvbx7zaYhQfZuuEtvwPwkkNBJp3vrnQQH2zSd0Nwspi0/o4kHNnS6xYFuOqp7LgMQDT8FtAczUhJFgjEbWBI/Ykf4+3o31lkQHI4CccQuBpSCAcvPR0Z90LxWUHftUYI2ASeCYux1wGUCJ/8Wtc0BD9VICRJAFPKMr5EUwYykgJDERTA8pdnBAcH1eYOhWUxmmYpKQzyp4ESiwb3RREqQ45Cpbc2NhDnEAVZhTUirO9vmASl2akKzIUp/eJHrMj2uV+cmy/7J/YvPEz/X15JLFG4ut+MG1pEF7HJIfB6BcUG7VJ1jkv56VcmAT7JUBSrx55go8gzExg7m18gBSDc9NBDInBSYg4EZn0/yTSQoQVvR5UxcjoT3EEAkzxJvbqkIFdjtDR33yHC2hsaNKeKRKtnzpgkHBMCFGOg0WzTC5xI8GOJRnEf5KxVhPEtzdpQD8ElraUlafm3DGF1lhJD9ALOBwx7W19ShKbHCAMsru5i2IbMFw6BqGeR1SmWB0wIY4uet1SUzIwYB8iDSMkfipSoGA2skyj14U8ElYHT4AOjJfBcpjcYgs+IHWdQk1p/DNQPQc2/8vjkIzJ8Bl7mvAJQwhzURxWqA4R9YduSQAActLel9rwAB7sF3hnsgdn59T0Zx7Fc1OMT6cNYaiaGY0ZIXCGOcYpI765yRUU1cME1RKlknZvToQXJvYKE2hsIz6NfyHAHnNNkDG4wCNeyzfZZcKmn9/b3W2poSC0iAp6RpSMJM4DIjsTCFSWZ96grfhZKDAUm00tsEam5tbFm6udkZLmjGw3IFpEQLvNEZWuw9AFp0yokNAGPzc3POihUzy5nzFN6MNUd2t/xspEHrgHNsKMaJG9fE3FGBJxA7yOLA0GWtck8V34JcXWz+cH/4/NxH3SOSpSZvhjn7xmxoeMiuXrum9yTJJO7SgCMZI97RqPjmeC0JsccuH9vmNQFCATjkTxMmpEj8AWv5Kybtufas1urKyrIKFzdBRCorSI4QTxQrAmtdZue72hs0f1xyxxmTanKpMRq12T2eu1+HaxQzARJN2jFsJx67508waQaolv56XXuBz8LEGgnwwMCgAGbk3Mhz5ZECeMMoeE+33X/4wFnPoRkLW4aEm89DkRcN0SPTnljDnojNWO3fIDVA4SGZrCC1wB6N8ksUUGpwhTMjbHzdVwFXLRntM56B4nyYAmQdanpADWeXRBTbP0wgRqM4nqXMzlk/zc3eLKTwp5BgMkSSb67zChgowAf4gP2tAj8UD0z8MSAfgFM1x0MDVBMjIWdQhhDWLwm8S9CxdhslkaUGR5BV4uwRs6uVoo4CwGXG+OK8FFChM69ZxQD3BANq1i/X6ewiP3u492qapnwf+uRV9I/w+ybJqMYGW1/fdECw4kA/+Y/nAS6B6DKTLkFAnOY+IOWF/4HHWydGECuJdEjUIaXhXhB7AjiXlxZVdNLIBvgBUPOGMM0v09olpsqTCT+rjJtOUozvVtm3znAlTvX392sSiQ/FOsInQ+zn1lZv/OgpOSGEBh5xk/1DfCIeyageA2JMDZEhY7KTaw5gEPuGxueZM6c9FjY12fLKknW0e/OHa5I/QZhevXjpsg0O9KmgxESQf6dJwbqGwUZRpUkUJpkSjQJSAdf5nO4nQzMlbTev3hC4pkmncsVGxwbs5VPHrTWXU5FNLEGCDy+U06fP6Cy8ceOWNyGb3KSQZiqNSo3G5/M6g/79n/xKEwIrS0v2+48+tA68MDLOTk83N1k+v2qtmWYbGxlQMX7xyy/tu999X2aaH392SUba/UODIh0ANsP0r5SL1t7eKmkvAH083jbyBdup4G+Tsd26S45ojwfwi3hCc5mcTxr8Ub60XBZoR3NMk8PBo83XsZMKJB0ZiCkC6EMcZA0oD0wyOeTnO14fUQqMf4O12NfbK/8FkYOqFREAAGQF1mCkHu47QCKNO+ILzGUnE1WDeWRGEituMOka4mwYnleuFc8VmvU0wcr24w8u2EB31ipVWNBI90BaSKtRgUfF5mZRrNSFpWXJv1lDoxjvgLXcZxo/xGp5voXJahoVsIiZ0iPObRULtraWJ5mXVBTrbQ097ra0TNEr5VIwNK9L231iYkoyY4BbgAdMJSAzSQyHsDA1dUgG2dwL7hlrjbOS+0sjg32MxCH7jPMNmQ3MtPmer0EkaRqsM9di77593loa92w7v2TdHW22sbZsmdac5Tp7bXunZisbBfvsi8uWL+xa7+CQzl32Q2cXEy4+Lba4sKhGCs8hTp4y2QepbHkZz5gez8MbGwVKEX85l5iI5zOJBCUG8469cuoVTZH+9V//rfX0+F6NkmAQRSS5S/2SzVkZecNv+PGRi0RJUe4Npr+8F5OnxGHlmJx1qgMcTJPUXlODMdfIiqbayKUyAuAmxsYsv75ly2sbNjo1acXdqi1wPb192r9inWOqvLEmh3bOK8AjWNOQtSS7uLdnm8WCE6fCuUxuD4irBj31YCiInH2PnJL7BCKvx3nHPpNkbjCJp1Hh3nQ0M7OK4yQzkuRBijNM0qHNrmaimms0apiU37FadVdN0L7ebjt5/LD9/W/+3vp6c7a2umm/+NkHtogcTy1h3b1d9j/+xz/Y0FCfvXb+Vfu73/yjvf/+m8qR2PMvnz0n4g5yqDev3bKnz2atCjAt2dNt68hl7Rc/+aldvXzZ7tyetkJ51yqcTZzICVNeTi0BeHvhzTftk08/dQZ2EtZ6zrp7u23m/j2BwV5jep2APLM85RRnvPYgv+csPHrosJpaqtGCXBO5COcR91RTkSIFNIkg40Cy4wgC9geRT53xSc50Sp5ukvSMdYx07v0ch8jBhZDfuvyLT986+cyJN14/uyQjX8j0RI8Lr6H8zIt+duQDfN9Z6K7iwLmkfwu+jJLRq7jcD3k8X/73PevvRY6FPL+gRkJLJmkNexVLJmr2f/z5T626s2nVctHaWrN29/aMyE+nz72q8zW/umIduQ7Ju+EjMXlo0oYnJ626495aTMgszs1J8g+TbCb2iXt8dmqP9o5O29PktTOq1fQPdSBYTLajw1pzWZudmw++QUxDZ+WZtFdrsFK1autbBavUanb42DFN7URiZZxW1KQsgH82p9jHhBvnFO9PvCGeMFXIdM3HH3+iHAwpbNaM54teowJ288wgJAg/aPDaU5P6oTYEWOc8i75bPIdkCqJLJEsxMcIaJH5RXzgJlZyEydLhwX6tT+4ddRr120BfX5C0dFlA8grJVguLKVtXR6fyJXLO4g4yh+R7O4pPJ44esmeP7qtRUdos2CsnDllDDQPjhPIqJk+qlYTl84DyNZufW7ODB0cljTQxOWUz0/dscnLcfvfxl/b226/bjes37fSZU3b/3rQNDPfbytKyzt+9WqOVtiqWSWft8tUZO/vWWbtz/4ndvPfYOmmEbJYsmYEAR0N61UZGhlU7gTfR8HTiIdNo7inm0lpNqqXBOmioSWaqtUXrlzwF6cIXs7OSSWWtr6+uS66WNRAlhCPhtjlBk5CzB0nglM6h3u4ua26g3sBPZdcWF9ccc0niIdRkPf092q/sx96+XlucX9z35iOnRdqRyVUwD0gA5Hn8nZhOPuSTFE4+Eimr5ookUeZIUn5h6jQSKeKUAvs15kTfbFTga0T9yz3ivvGsm0MzlLqPtREnPJxI6zLlEKHkeylSCBgaslUtmqBlT0jWinNNWAI1FueFk6AkzUh+B5kZOcNy2afHA3bJPeOZ0NBhj3HOCPcJcY1cUdga00ZBvltk51Dnx+la3j96AFPr0gR2knaQXdcu/LZREW7Dt//7Q7oDb09NScJERjgKUK7n7MU8xfLOPtAltjrmZMEwOiYSJHQEBEBAT2ScZUFQhREoQ9nAGI0M8ChPodH0XUx1MgJPCaAUywCSAnoE0LrsDQUpRYyDt252KUA84UkMhVVknvH+21sFBRLYypHRKc1suqCNDUqOnjx+asjgYfznEkM+Nsp7ScsRWQSYirC/ag4Ixf97oHXwjKRLhphBk47PDUhIIOfaAUM4/NHhg3UEiCJT56CvzUEcdRz5Hgchhy3sRjGVg+RTDMoAL2IFEQyrrnGpwIluZdCJ90aQ+3tIgkn61FV1l6N0A0k7r6lAWfXmixcdbkItRpVARfcLIdkTu1njdJ4QiPlP8BVw6ZMIAjGZagCIDT4YcfJDxXdgY1Aw+DSIA3sky1EiQUCt1ZXweXKGgVTKzdCk7+2fw1lAzi4TeyMAkFH/fC/4Agj85l7Jo8QbbDLbzLTKI6EU2J+1PbTOkxpzBhjeKRR1QHS0d2g8FoPDodERMb4eP3kqjeVq1UcIadwAwo9OHLD1fN7mkeaBBSmteAdveB4wTwFslFCXdpxVF8BkTY8EbWnWl4MVQTc2NLv8YHPDNz2zAApG7Xs17yTptSsgJI5mutZmq4pb31dfMxJgnLkxLkk+jRP3peDZbBfRR3TQDmBWDSImHJAVCcCpZGT0Odx8HkDfTdacBQq4RDFLUemAEqBLkxpB+EIw2RKZbiUmYcSEcvM77g9AVmSdRqk2TKyIGVH2iCYFDSeN/lJMktwD7tZYX1UVcNXKnp08eUz3m5hFgiAj1+quzc0vSGsYnxP0mElM7j54am1tKUukUlagoYSUVaZFoB/MRpmF8RowGldXXU85mAZqkocYwRSVPCdchkXa+/L9CM81mEyrOctEUxif535SoEa/kNhI5oGTHLHXASEpAPj8FBY0j3i2JEsApjRCBWx+YwqHUXvukTRPYSuWSpJ3IVY+fzYrQAgGK6+/srwsRkcEydzgzj0qmB7hWuOUE9cFc5xrZj8Auks6KJ0WIEQ8jD8vE9VsTjGa9/E1TMIKEO/sOjEemT7SdIL7crAfYI2yVijomJKB3cprAb4zlcKaQTIFcIvEHHCKtcC5wJpxw0dn9OMzgdyDG2r6fmOdc/9IyGFuu3G0F+rR84I/s+ZJQGluCFBS48mN/1g73P/YFOVc0VrB+LQ9pzUAiErcB4Ti9Wk2aV+roYver4/98rvy9Uin99lpDhK4lJTeN8RB4gn3kOvjOcPoYg/Q9JGUhRpnSe1jng0FLzEqNu19utEl9CL4r7N/fwrOG4wUpPHZtXd26HMw5aBmcpiioyBxM/IQt8PEF7GPop81TPNb8nt7ex4fw3OhoOEsjIxNHRXfaH5EeYcYC4mD35yoA1hFYoozg1hFsaeTQtMvFM/4DW3KIJXJS5oJADCc6wLXZehZU9znDAbQ43ni58X3aXxSaLG2sq1ZAXRb+bwKaNh/vAdyKovzc26WOz4m2aXnL2BEM94N2x4g2KUbZdYu01v3htJ6i74EGIWG/IT1x/Nymcma5be3VQyPjo3Z0iLN8w2djTDCye1obsAK96anX9M3vVCifwvxCyYryUZvT7eNHxi3ZJBKQ/Odgg6Q/dKlywKJYJ7TVOS54dtEI//F8+cCWtjvnJ00AD2mJRQfKYK5x48ePwogVF3To0vzi4oz7dmcdXV2WLGUt3fee0s/jw/Ysxez9sUXX9ng0LB95733rV5BqrJkH334kV9TII4ASuJDgxMKTZETJ0/amxcuaO3eunZNkg2vv/66rmt1adESDTAuAT3q9vzpM7t2+Zr9yZ/+qeU3i/bJZ1/KW4C1+pSCv6tL93N9fdUGB3pEBjn9yqt25cpNnS8sY4gQO9r7zZI4iRKlLoMYNItD8c0ainkP3+O+aOInNMmQ+eAec55oAomzOMgwicnKa3I20rAM0hq8jib9Otpd7nJ3V3JfMmwOZ6jk2SSP6WSXf00IYkKrYgfGJwSsSb41R2MWAJE4z3Uw++hnM/Gf/KoxUbPmRoDIhJ1++ZAND3babrWsfKi1q8se37pvX168bgcPHrWZ6Qc2efCINNuRVs22Y6LqMhdouCMHA8ihKTzFTGJrXWAIUiQ00Jjobk6l7enzF2oOMQGHMgbASmuGBqWDCfgqcZbikXD75m3FUfbDo8eP1aDmdak7Jg5MSspL8p3d3fbw8SMbGx9X/kaz4MSJ43bv3gPJQ7DvMCQ9ceKkJLmcXLNnrS1JS9QrNjk+aCcPj1tnLm35tUVrzxID61bea7COnkF7/HzBPv70kjW35Kyy5z49+1OBarz45BzAPeQv1gN7nrOfaRDkoYiTagJDqtjcUuyQ7BNTFx3tdvjQIXvx4rm9mH9u5147a719/fbrX/+tfIk4T3fLPnEVm9iwZ6lLmKZASku+GwnyrrLOEAA/EWJUZ7iWPHkMLNOtghMDRMBoBMTftSS1CZGksmuTY6NW26nY0tyCHTo4KXY5bNxdSEHZnAxamdR8/fx5y7Z5Q/TuzLT8f5D4Km55Q4QzS8akyHYiB9nYpD3Oed6Wy6lO4AuPDSbfIdTR3EDzG0kzfgZvn31AXuBqi62uLluxtK2J1cZA7tHchQBYvIFabX0zr9chz+P9eT3Ofs4VpIGI+XiUAKSeO/Oq/eVf/tra25os3dxoH3zwfUkML63k7eDkmH300W/1PH78xz+1ledPRdz68otrdv/BnL10fESN2IG+fvvdh7+3BKTAJnxNfCp2anLSutra7KuLF212dt5qTGun0pZIce0uJ8o9ovamoSbiX/CI9Omsst2ZvhtICdRdTgYkJycWIY0JyclJCzVJ87x07LjOOGSgOTfYI9SZND+ZHqVWiLmTJoFrSMxm7Pix47awuCig79KlS87SZp0ERQL9uTmlOMl0N+scDyrqiQjOifyFiXxbm/Ie8lVqcI+ndeUQ1M7e0HBZWOo6AbCa9naSFK8jbxukFoMUTSTGiGgXqH5VgNowWS7Cg/JmJHtGNOkln7RqxRbnFm2wt9n+/Fc/tUJ+2XZZP5k2u317xorlin3n7QvyaCKvzNKAffhIMeOVM6eto7dHExWpbFb55srT5wYZvak5JRk2NY7rNeXO3FdwCnAA5GxV51SrNjA0JBwDT5e+wSF7/PSpmP/I8jUlkNLqsd99/KkVK1WZaTdBYuro0HPkzJ6+O63XxR+LOPL4yRPV9sgEkdcRU8i3mXJ179AW5daff3HR/QdUS7BoXEmBL/AT8hYn3fl9Tun5bisnEGYT1llgf0hel291dOb0PAGEXfHBSRzUcD6pwXasapoFPy3yOD5blJOmtnCT+6RySvY6z1WT3zQmyrs2tzCvKTzOO/mZJZN2+OCkPX9038YH+mx7Y9POnDpu60tPrbOjTbne2NiI4j++BDuVoq2vb9vE5LitLq3Y0ZeO28ztaZs8OGEXv7pkZ8+dtZvXb9ir507b5x9/bOMHRjQpMzTYR7ZGRWeppha7efueHTr5kl2+OW2PZ5ese2TM5nluMnJuViN64sC4rawtK2+mSUgj2c29nQDB+mYqU9hAIPEuLC6oUSECVamk+odpf0mQoeLA1F5vn91/8EA5MORO9whl9SMDV7edXc+T2aPJpoRkLruyacn5IWvc2Jy2/FbBeOK8b2trWp+HewwhAE9C6iZqTZoVTpShObmp95J89PNn9vLLL+vcpSkG1qQaVtP/ZeWYrEnwFW9M+nP1CYuvpXRjLRMxMeFNkpNziWAm44jvNAPZT8QK6kVhiUEqkxtBjUG9r9qPZkUg1oKbIB2pWiydcmnXlMuIc3ZGf11yM+o2lxxrdpxCObzLYjHdxdSz5K/k5dIks3RIWdQYyvlDzSSZaibf8a8JU9zyx2tEZcGJzeAwEJSIDXqQIhhHZvO3jYo/JHz+22sJd+BIm5s3is0bGM4CguVd5OOhUTLIGd0OchA8XG8a1jYjlxkVEQQLNh3JMAwfDhjpisqrwXW22bhsVg4zZ9u6drEz/zAijaY6bnQcGaCA8dKMJLFgVIxCS6bDrmEZjUrdQMvBbOl3V90kSyNUsDKa3Mia6QXpUQbwlwOaYEORwLUK/GakTTqYztAkAMvcFpkqXiuR0EFMEJZONCyMAFJ5EoxkDqBZl8BDmcYijyMpBZ8Q4brVIS2XFcC4HxgE4oGgjm9gc0r2iQKTzqvAYMzckvu62VEqhHvrjzCMNzPKD7tYusk+9uwm2DW9lhhWYve7TI3LelTUfKDgjlIEYrkI0HIgmOJCYE5gDYq5UvcuNcmlyyuhffj1ZIAmHAIz2QutMBEhrfLAoqPAEKPe9dSj74dr0TqbnLUpiYLAvObzRPNzXgfdehpHfMn4Dh1ang3rM3hv8DqSiAE8SaWsq71DxX9hG4bbrq0ubVlfT84Km/58SXJZMzR3CjB+066rvbpK0dQsIJcDfHB02E6/ds5u3Lol4yoSX5J5HgJGUw5A+SQEa0vfEwBH88WZEm7s5s0Adcy15n0vxD0WGdP6XRlj+qHHsxMoF7RbAXBZG67n6nr0Yr2gVc1YZADkZMwFQz0Aw+wvitUoycbn5pmoQON7gVHp0zL+3HlTjUzC+AimyHx2YgvFPGa1kvhCAg5tTZm5ptUoYvxSEyHhGbH+NK3UhJyUgzTflCKIEydi66cYraS56UZoklsIZzfMffaJ2A8U/aVdGxzs1doa7B+wYqFkJHmVXeSC3Ig3i4ltzWx8YkIm6SVkCzpy0ijmw/NMJUOgphyNTH+GJNqZVEbX6M8MxhH/9/1Gwqgkp+jG7AC5US/aGeMAziQizvyKGru+FtyIy5nHX68HgDlALmID4CnxhwQVxijP2OXnXOKNtX/u7DndZ1huCwuM5NNkwUyt1xPEQkGMQjWRK5j8bSrxhRVNXOdZU+RoCkVSCz7ZEEFr2J4RbJPUTJgI4t6Q9EeWd2RI0kTzaYWqYinJLEkirw8wyOfm3shsm+fQ0iJ2uiYu1tfE+MLfg8+F/ilADkxnNdTE8NrWtWht7wUWihp8TXregKOMB7vcjktT8Xy5Zpq76OtzXngzxieHNMVVQcrMmTGRyad+fM2TaZJabzK6+bZj5C4dJOmDnbKYXXxuNZiZhAv33JtBzsSJ0kM02aQdD5Gg6qA+n4tzhYQ4yp9xndEsEgJBiqmCIB/jU2s+8UEsZC/DymIdk0xry2h66mvN+zhZwYbyaQOmAFoUb4ntJP1cK88IkEDsJ5qSQX6PNUUzibXLn/msPJtqfU+xN/rxEKcozrku3gfQnEaTmqk6zZAydI8S9oDG/YNBdCxWeF0KINYlk2+AyfwesUfG62ESgXhEEcLkEkU3YC7nSXdvj83PzTtbuDHha62vT3r5IiYEU2vATnTuidVIatDk5uzgHKZbDzMAACAASURBVKHByf1dW1sR0QGmN3477733jnSH81voTyNZ4aASMlAwKQHEyBkoeojXfHY/F5yBFY3lid/cAxrmN27e9Cm9YlnyPIBIkY3Pc3j65KlWHebW8pNSDPTDhqYSDGx+J6890qD4xXQI00aTkxNilZeK7Ek3k0dGhM+JeaWTTFyWhmethmJjQpJpNHN55uQaTOPy8/s+Vo2Ntra2KqC7pQXG+brtFHd0Dpx65ZRkFu7euWa9/R126vRpAT28x6Wvrtjsizl747vvWFsqY7WGhH328aeScgKkhHk9PDYqhufDJ0+kSwy4jbcHZ0Rpe1tmvjTumKqQ7J0BihXt0NQB297asKuXr9mZM+dse7til65et9EDB6yjy4FrQDTuORrSExOjAu85P5qaUjY7u2iJprT82GRwGnJFn1L2XEgAQyiaiQ/yKgr3zfcY00NM4/oaj3J1NLMAf6N3TzTfZu3xPsohNX22qckheXzQlAgeXXE9yASeSdWkPzcaR5o8U7zwWM8u86aP+9Aof2tiUoOGE/kzshxSOhJoTZxE/jGdarTtTbSdE/bed8+Z1UvW2dNl5cKWs1+TrXbpq2vW0zNkL14sW3dvv85NzLkXlzECbxHzneYF0xVI5QBiqBFW29OaoHHGucmezLTiB7VspQpTeJ4Hdnd2WL1alu9IKt2smgQJKWRShgeH7d7MPZ0zyG8+efrU+vsHdM2sz8nJg5JEZH8A5j1+8tgOHT6sySnuEfsdGQ/yIRqXi4tLaiJx3tLEJMesVArW29Vub55/xWolfGtarVYp2mZ+3YYnJq1c3rNipW4bWzv21eVbtpdIWTLdqjjnk9utOvtXlle9wdTba8vLK7oOZAO9ke0eFLy3M4PLmuIk/vrkqE8Uu/41Mqc7du78a9bV3WP/5T//tfJiTU8jn8OUQTrtXnm1ug0ODihGsEa4zniGQ+zZb54HT7vYsGBPl6tOKvHpOZdkRFpEBCFkl9IZa2pgSnXTjh09bDdv39DUEf4TQMSUmbXdmpjng/39du/ujOIS18bnFQs/v+HkqeADheyTpEBTKclzrec3NRGMRI9PsCb1fwe99/TM0dL3STaf6pV3D98XI39PoLKAeIAmNYx98o0zCE86NWxUQ0BWwCyVWgRCnuffVEKjI8P28ktH7b//3W+sI4vkWsW+9713bXFx1RINSRscGrC/+dv/ZkPDA/ajn34PcR5ryWXt/t1pu33rji0s5AVM/vIXP7LrV67Z4sqqpimQOGMvvH3hgg319cqjginuJrw3aFJosgRSnxMMNVVJLbO17fJh3CukjWt7du369TD1CPDnOYmAriAf7AQFvPocODxz6pS8yB4+fKS9jPzOoSOH7fPPv1ATkPvJXQVkFXaAoXZTo7300gk37E4k5LniUnf4LrkEEzGQ92QCjxjGemZ6mThAbOSMQIaGHEM+YZJ78vxFdV+cTK6UtUcigEsdI1P14MunGhn2tDXodXg9pL1EFgw+eo5Z+ISzPleo/flcO6WCdfd0iPjIGp88cMBWFmettzNtf/anP7fN5RdWLm5aWyZrt27dVY3w1g++b+X1NZHcILyRxy4uLlvPQJ+NIT1L44/3qDdYfp2p4RaZPXOfVlbcK4t9hLF0d1eHTU1N2KOHj+zwkYMut0pugt8gOW4yaTdu3rLW1qwNDA5bKol31ZI9fjZnmbaspduytsXETnOT4hV5hAB97vfaumILxtqcL7DyyeGQCEKyksnh8bFRGz8wIfAabyQk9EQOkVoA09iOHVHLQ3LQ5xMWQMPKCTmOowQvFNnsMe3uyhiqc5oTqrkAtPl35Pw4i6RGoGlucjfyGAzl/fekgmENyi3cKymhz8QZLYUQTfObcjJ8T4pl5J8gTWXkuwX4f/zIIXv64J4N9/bY5tqqvXb6pL14Mm09ne3KB0dHB5U7xFocCWRkniF+nDj+kl25csuOHJuw6zdu2mtvnLcHM/fs2OlTdvGjD+3w4Ql79GjeBvs7zOo019osnWyxR09nbWhyyi7fuGvPF1etexhvoE154Mjfa3VJgD+yuTQZINGUIbZJYtaJm2Lui7SV1B6kdkL6iQlw8vCNzS2dWaynA2q4z3ve1t5uM+EcFDEJgq28s8ya8DSFCIUZOrUmORLer5WydXbkNL1SYmo03aI8lclSkR9STC3vBqngZsXLhcVlTWQAqOs5g+fg09fSqvraiWk+wel4Go1ybwI4YaeqHMXzWVfz2JehDTWSN1OdCMiX8phAmOW5k5uxFjnTiM8QgiCdyI8mSFYT72mwkXOLNMh1t7RKTlGND+4vsqkd7S73K+nzr4m6EHEiSdSbR04+juuP1+A6IkZDTBJJWyokSPR9g6wYmniSzJIULeQUJ4fEiQtiV4xRktrSjvvXX99KP/2bG/LtX//3vwPHOjr8IIlSOiRfSK9QsMhQ000vnaGwJ+YP+G9Hu7M12LgwtwFaAD/l5cBEBYxaNCrR/6zuqrPc0cmB4ux5N9J2hpmMY4venNCURgOJMpMVLldA0OSLok/dQ8j++rP/H1a+QBEAmdD0oNjiMxCkKOyVpGzmxYgH3CHjAnSem1vYH8WKGniAAgP9fTa3MKeCG7MzwC4OTRJnxuqUpAamIGA3waWtpU33jL/DNCHxioFJslEyn0UWIQBdYkOnBPpt5Dek30lgJJB58PUpAxJyl/sIQJFMb12Sw3W0ObwoKF0+RcwYAdp+f3zyAAnlhMs8ACoHySCes7TGCfIaH3ZTMpft8WaQnjMGwUEeTCPlQTtdQZOkX+vH5Yk8YXCmuA746D8RmCuSLog+GMi3UK40uGQHX1xrZM7rOf+bw0gHghpFPrURmafcC/89N0DlXgiww3A1MNcZpdSBFPwvOAQyjIszng6rHvmZ4rY11N14VRIZ0v50oJdfBLhi/apI2sxbsVRxBj+SZMhaofmILvPquqY3AGQ4jPl5kiruKUkGvxOBzEKh5AxHxjnFGnB2dmQTR9MlnzIKcSfoQarM0OQLrFyf8GGMs1LZEUAJQzAm36xJfh2WDF+s62juRPEKg00AdPgc/DCvqwSgFtaf56POUA/yMtEg2b1PktoDcTJGpUyYMGJsV/I1+zIlehAaz4ymt6556kwKJaBKpgBJ3DR8f0oofI+CPEqWNdBdMIAWb3JowqTufCmtJaupgEPnHIAPA02AahoGy6vLlkjQyEDeoqJUOZvtsNmlVWtoSlgSCR6xuvBG8LWFYRx7nDhJvAPY4N8i250kl2esEV15xHhBT6EPM5RrIpGOUzMAJWrGNDtYLu354GfB93i2vI4kmFhrAr5Y8974evb0qctilXaCHr/fe+4p94hkd+qQFzvRyJjn4V4eu7YpbWzYNCRLda3Rrfym4q7WAgUHRXzcT6GBwsaI/jY+CUPs8HVJTMbMmdegcctzlrYq0h5MpyAJJGZwRVJKkqMK0jToccd7E2MbcdsTP9ajj+iz7tWgTTSo4FIxyuh3uSz9dn4GPwNMdYm3AE1MkPBeJO/cZxJhNeOQf4C5upG3dEuLFcol908RY6fZqpWq+/4wzh4kBKR5XCoJ5AWciM1nAGL2Pteg5vS+14p76ez7NIQmrZrvNAyJG5IvpHj2s0aShzqbnS0cJds4e70B3OiyCEhaIKWFtwK+JvJU8Ek4MR/FyPLJxej5xOfg53XOJpjQ8nOABF5MTTwdUk4kYO0BHtFU4EwE8ERTV9JbYQLMzzqfAOF30HQHAOTnYzFCjKMojrKGXCPnNTEKwJVYLm+nUPg2hSaJDDg15cJ9xofIC3cmtGh+RXADBAmGJCCio2EObmASTy4Ae6zG3ki7YR55Bs9f0oIQIarOroygRWy+6GzBdFVNO9dI7u7scqaV2LsuIchEB0caa7lcLtqF71ywnTKgDCHP/ZQofgBl+XnJQe64BIma/AFsE8sseMA40cAnRzC4ZzKOnwesJf6wxpeX174hG+QAOdcB8A0jj/scJycBGOKzokHIMywWtuRpkm1rte+++46lml1mjuugAYqsm4NOvFazGvasSSao1lZWVBCyr377z7/VfuZeUnAj08J9Ix5BUCEmSXqwZra+uqafPXXqlNbQ7Oxjm5+ftbcuvCn2aLaj0+7fe2gXv7psuVynJIlY05tb+f2GMOe8QHlk9eThk1Jj1PcCxeGemiHcr0MHp2zqwLilko1W3imKhf/s2WO79OVX9vNf/FKSYB99/LmNjI9ZS1urvZhfEEMbUJrYcWB8yDpyOSsV8FFhAhgQhnO1JENtnhNnPwxu3huWu5uKenwBLCFnoznIOSAwsYoHiINIPH8KZuUZSffyIRYI1AlTioDWxCNeQ01AeXR8LRsqPzIYg7rvLkOps5L8Wqm3n+eeJzrJwPWdq5IhAVBQoxA24vaW9qT2gvTgk3b61dOaKES65NLFT62tFQ39hL35+is2MtpvW/l1b9hQN2ztSPopmWqzvT3829rtwaNH1tvfo31MYwRza4yruZ/Iw8Bc5xxl/fMZ/BoDcUWTWXUBTwgMcb+I4QDMfb0wbeuKS5BqaBIi93jr1m01wYmJEDTGx8YFmJILUc/Q4NReYZK8UraRsVE15mDrEouQSoFhKsmyVnL9mvX1dFl/X691deZsZuaWLc4/t9dOn7JcstF2CutWryDp47KJzZk2a2rrtBdzy/a7T76ynT2zw8dfsts376jRAEgvAFy1ypZPYQcJMYBiSZoS73aD8W4AZ2guwq6l0cjnKhS3Q+OQnLJir5x+VczpX//X/0fybNIC3/M4r3OSmqmhQcSy0k5BrGhHB33SWhMUZOmqsZxkJbnUMA3vJtWehxBbxNKt16Rxjuk2/k/cgrnnczonCoDF6ZSVdsu2lt8OZ1oCRocl6iF3qCNp640I1mmOqZTqnoAtYj7XrM8VJGVFhAnTdsj0whbmTHbZS5p3rba+npf3WaLJwT2ucbPgMqY0Kbh/TFpBFiPmkTtz1tBQZq3J0xCzagDD4JWF5BeyKNzQZFOjTR4Yt6mJUfvnf/wHSYeWd3btj/7oxzZ9976lM0jrdNk//MM/2cTkmEx4r167aT/72QdqTiJx9/g+zPvH9qMf/8Du3pq2O9P3ZKa9XfKzfGx01N658KZN371jT56+sD1LWJHYgzSQWLw0EvckX3X06FG7euWK1hJfkDnIa65dv7GvCuAxg9QsoTrcRQ99ih69es6486+d1bQbnhQ8dyZ0aRryOsT0mN87McldQFhXTPRBBGD/L8wviJDAecGZz55THJG3nJvtejOXnIea3/XuYyNB+X+oH8lVPA5S71ZC3HJJTF6bC1LOHciAyr0U077GMrguyfHJDNeJecQWyVepmeV1Jeu/q6tDgC2fHzY5hukbayt2cKzLfvnT92x98bnVd3dEULp5465+7jvvvO3gIjkYteCLOZ0hIxMHrGdgQJOX5PHsledPnlpTI7Vm3bYLRVtYXJJED59pYX7O+vt61Gi7cvW2ZXNMs7TKXwJcg1qTaW0AerAFzsBisWJLSyuWbs3aTrVm5T1V2JZubbHbt+/Y2nreXnrpqPKWq9duKG6ePnNaucjDB48E3J6DaHfjhi0urdqpV05oWhMZnMmpSfvnf/qtpivY9zQqWAMOnjqRUETGANiyDqWUQUNCZ43HEW9uuXQsjSvWAPkGe8Drz2CAHmrcWNMNDHBfSvL1Qr6QfIS1wRe5Kvt8a4tJVxq2nI0r8thjTSDRSBlDXcKZy5p4+fgxm751245OjtjqwpxdOH/aFp49UENkfm7FRka7RWLivKYpSaOGeoGcuq+/x+7eeWij4/325Zc37bvvvW53bt/WRMVXn32p+/bg/hObODBqywv4TbRqNOTR03kbP3TYbk4/sKcLK9bRP2yrmwVNbtPsIf9iQhbyHHgV/mSJ4DPHmpBKRcB4RDgNcmyPnjxVM5X1DvFkfGzMpmdmbGxsVB6T7ifRYo8ePdK9iY05XosmEXlr9L1TvbBHvkSOhpyfy3Zizo5sI+cS54QaJ/hkrW1oPWliAHJWwHCI2ZzbcSJd3nXUFA796YvzXcop5GxpnxJ2byAa2U5S4n00QVqvq57iy9eRSx+pHlTcchyJM46mDxODrEXqcybCHB9EGjyl/a3JmtDkpAGkhkoZvNI9bTkwIAxHHI88Vk3VTEuQG8ePDD9CX4PKQ3Z3ldt9s3HKn6VCEUgh1E7R38In/LwhEfEb4iA1nte1rsKgybeAdykfj5J4ocmsW/Gt9JOviW+//rDuwNFcNoxWecEa2doCtsKBAuOBPxMEi9vb2sQUKAR6AWth1Apggq41SQrJiRiegSFMQS096sDU2O9CBsA8Nh7EDG+iaHcWtDccvgbdFZpCYsX7+OhhdV8eRIWvWK4OsmjMHQYMnhuBDcWoL3/m9WFJELQZEaQoAuAjoSH2uSZnXcWjM0Awt/SJD8AvmQEKeAHYb9Z1U4ATRGCvcADjPUGA5c98BjFdgmE2n8tB5aQKYIBf7icJFwcBvwfbGDCcEEQxwZdkNYJRqsYppauZdk+D0LiQ8VIAliNITUIDGKj30KgZ2r5uREiC6waPnjTGpg0MViWG4UzwHM7ZN/H1Y3NAQBr/HszQ94fRIrAuwzWXDRFrCeBMgJtP4agRo6kRvw41TyJT3xHZUGBEc3VvULlPhQd7v0WuOyht52BQGU60/cNRywjmI4BwkLtCusMnEQBS3BgVMKawjS5pSvcNUJkiqRNwUyyCJmlEV82niGB1tXd2yVANFgv3S6OZZRJqU8IpcCAYukctYQ4trjWCsTyLyB6iSGedx6aP2Ajh4I7+MN9kBvGZSeDTaWdFwlAGBOIQp1DgsGV8l0OT/cFzEnOl0RtAOhBVx/lUkifvFLeh4RU04HlmJDTR34Wf83Xk+ymynOUnIx39JoE33jBgf/nhrbHsIC0TwT8BdwJWKD7caFjPOnga6JYw8ROaInGtsUISTdxfT1q0jtAVDmsPYJnrhK04MTkhsBUwgqYOci3cs831NT3nhlqD9Q8M2dPZeVtFH7i3V94jfMZexrdpNu3fGzfFoliITNY4CSNfHoBotPeDjAXsSQACkjyuiZ9R00dr2acHlGCJ9eWNn8icpcChGAKU4UsSUDXWRE3j5Uh3SLZBcnU+eaE4HTQ/Dx08GJoXFHMuEQVjlYRy6uBBTVAwsu/mus0qHpQYNzVLgiSCWtKIVmEIMxZQGkDNr0lmnADKGSZdqjY6MipWD2xrXidOqcUiw+NNTcVSV3eXaxRTiGxu/quY5H48DXbo8CHXvF9dkazJ8PCIGs/sDaSeSPRGx0b02Z2Z4tJcAFbywejoUJOKYk+msYwEK6x5sGJfu4ROVWzN4aFB7RGeLSxXPm+U3pG8Qmj0a+pCwL6DimLwB4ZeZMJwBnCPFK9Cwq2pIxUgMb/wpJZ/2580LJWcWaTGsO8hAc6hSRQ9UXyUmNgJeIyJ37auTfrd4eUFNOP9E+Q6+JlUmikFPneDtbd329DQsN28dVPnkNhMsLBl6O5APqx7GE/4FyTTDt7TmGHKhURdOcReXVJ4y0srAuvcqBvAFzPEtMe1APrwWu7f4YAcz4R9yKWStOOjwv7a28Ug2MFdAB4KKTTGI+jqY+Jpa0on1ZwHdC8wyRNk0tS05L62ZKx/eNh6Bwft7syMPX76zCf4VKTBkKV4gmnr0pQCPwA80L1lf9IwCIbjMjLe9r2vQowzTezWJoHEFIGvnj5lW9uc5XWBYHxeyZ/lcmoYsxZpJGhqlIkK5T2M4zvTMza7KDbPnD9nM3em7bcf/ovyBQBKnovWVMJ1uvnM8lahifNv1qCM6NGOrtXUPASkZE/wdyYFeLY875dPnrR3333XFhbmFSfUWE2nrDndLPalJLtqNWvPtisXunfvnlj47HfiIWB3Ot2ieOKyRm7+zufxaVhfkeSVFIr9A86CA5jY2sYUs9lOvXrKRiYnbfrmtH300cd69nt1L15hWhZKW2oauHQmuQQNKQgf3hTxfRjfykGs1taMvXnurM7+Zp0vGEIX7IsvPrdXxCAu2leXr9rE1EErcJ5CHEg2yWCUvdDV3i4Gf39vvwp4GJuAGUjS5JGQVLxMqqFJQ4Fny/3zM5O17UQH6RKHKWTifvSbcaDFPchYz/HMj81JTceGZjHgNoU46wYAx6f7gn+FSCGQgzxvI5cFUOIzcG/UAIFoE2QVvJBOCNDg35BlYcpodGjQ1tdWtRe4z/T9Tr7yinV1dss8Ob+2bEvzz6y0vWFnTx+3vp6sF/LI4SVTVihU7OpVpJdgJhatf3DI1iQhEowkK3vWif/C6qqIBUgs8mcYwiJu7OGHlVH+pClcq2tNAbqhHd/XN6C1392BN9WeWNA9XZ1qWLC+Bwf77dMvLtl3335D9xW/CUDvM2fOaqISk3aum+kbztsX83OKHejDoxUe2fXIVPG5Yemzpzs7sjYxNmIry/O2kV+2g5PjtvzihV147Zwl9iq2toL0557lmAxJNMmXYntnz7786rolW7NWkNwgRAyf5C4VPI5xZhF/kWQBVGNanUZxa1tG5zM+NXjFkGDC1oaRiiwVZyFkKmLldmFL5sonT55Q0+Mf/+l31tffK/nc2BxSXhUMQ136LW+1+q6ATSZRAZ1YS+5Z6PmhTwa55Ch7vlL2BhZTNzIuhjxADYS3VZDEJK6tra65L0jdbGVtzWoQ1JhQ15StTxsJrGK9VytBNpgJVgzb3X+QBguyrOypjhwygXs619dWV5WXQT7Rek6l9HypVVlPy/h4oIdeLrlcElOr+CaSRzN5tFNWY6WpiXOXhgjyv5wDxCtAdJ9Ixxye2sxjD6xxPlfVGmo1y7a02PjoiE1NjdnHH35kHe1ttr62Zd//3gW7d++RdXT06h797ne/k2fKkaNT9pvf/JP97Ofvy1Olf6DXeoaHbOnJY/kdXLpy02bnFqyhsdkWVlZ17wEwf/DB+3blyhW7cuW2S78xFUIfXpKqNcnA0ZCj6Xv10hWR4MgX8GEhR7p9m98LEoiSiIQYQ/PaJ7ldMilAybU9O3rkiDWJLV/XfScnov5lfdDIFCFMjHlIWQ1ed1cquver6xuWyrRofyEF601+yHcOIHIfiZE0V+QnJfKTg9qaqg9T89ErihpTk7Kq77zm43dcqjKoL4SzUmxqGn2h3iB2EKvVnBPRzieh8bMD3I5yUzGnV21d27MD46OSuGVibWFpRc91r1KyybEu+/c//75tLD6XZwVNh2uXbilf/OkvfuzTWvktmTo/e/zEnjx7bsdOnrDegQHl6Hy2llRG32tsaLb2XIdko1ZW15U3gwnQBNvbJc9pVhO8sFOxlbW81fYSNtQ/YK+8+rLlOnPWmPRmIlJde9W6TU/fs3pDk/UOjFi9sdGWyWVrdfvs8y9sI79t5187rbrwo9/9Xo28733vHYHZ12/ctra2tL127jW7ev2mYsjU1KRNTE7anTt37NXTr9qnn3ymhjK5W7niElCc8Y69uNyNky1MU2LUPKwr9o+IIEEqSoTBBp++4SzkuUIOokfqe909x0RECngMTcQdiGRMFOdyihXsC94DEi3nVnx98irWluTjCgXFn+h1Sa7KZz5x7Jhd/eorO3PysC3OPrN33jpny88fW19fj83NvbCJA0NqcGRSyOGt6bXx7uBcQa4KaUAaF5xtr33nvF27csXeePst+/ifP7HTms6YtWNHjkimDek4nuGDJ4t26KXjdmvmoT2ZX7bOgRFb2djUdAwxfmsrb/19fcqviANMl9Ulze3TUjRHWbfUa5I/8mrdnoUzjYYHdRPTsHhD9PeRozDtCCk2J8m2iHlBcuKLfJ04y/NiL8j8PMhrMcHH3uR5ScpRfmjsW5rwDvoj6cu+B/fy5rfvb/Ienp9kdBMN1pbLas9zhpLfMsX39Kn7V8hzET9ZEQHxXyuJdCLQP8irg5vsyx45PKGvOAlOrHeSb10xkPURX1d+gpyxOxDKwON2/IzBeLsfeS7TdBNECTUJ8FEr+d7r7u21p0+eWKol49NzeIdQB5DL0bTZc6IEOS3ECF07RG15h30tpQ/xmXskXIu8t1TS76tmC42XOCHi1+XTj1EWPTY0vLb3yY74c7G2+3aiItbQ3/7/D+YOHM62qUMZO54+ou9AmCYr6JoH0IVNDzBEMBkZHlZiyeYQw1YNhQZb29hQ0GHzZUkkxeKEkeKdc5oeEeSRjrbGc6segFUsUVw6o8G/t6cEHrDHN6szD2PnVx3GIIfDz/OlIAPoS5BQQefFqX5HeuoEDjSoMbwFfCL539ofz3fpBQdlSUKlha1A26hmDSN5KMCk084m4T1ybTlNX3AvJWVF8fs16uQMOfS46RYDAgQZKBm2dnW6EU/Nx/YFdFYoCGEW+KHkjFkHp2SoLFDLQR5AFXkgyHTXPT0ctAkTDWL41RX0OaAJ/BxwvK77EnhnXGyXwFzhfaQV725WDpKEpgw/p+AYJhpiwikprCBXJHZOMPn5ehzPp2nkbRAAncquB9z9DoL7s/sBLPmTIB0T0YbA7Prm9bmhlydM/LuAVAGALm2133HfP83C0aZGkalAocEijoemiLzbThOL+9+ec71KAesG4wEzqDbdG36uvbNdJtonTr5suY4u+5ePPrKtAhI022JXUhiSEPBM0Y0F1KUw0rhyEyajztbh+zx/Bw9g+DiD2keX3RQYUCgamXM6e5Ou4uOF4XnzrChU2XuwogQiiR3hYBvPGCkT9yFxQENAFoBGuM9uVNisQjgyL2S6B4s8mLizDgGXHOR1hrD0HQXSBaNkngrvseumn5qCiqbIKgRoJLj/CZMIxJLYaPJJjq9ZOGIlwEgVuzcMnUtX1zVr3VAXpq1rlouRHNgNmoAIUzTplrQ8ArhmjAsPHDig/f748UM7dHBCSWhxc9PKxYrGndc2tmxtu2DpXLsVBDCR1NUVE5iucZPNNmmrP378Zfy2ZAAAIABJREFUZD95js9SRRfAcEjs+FmZzO9WlORqkqheV9yUhJCatIBpGHSVBSC6b8me9Nyldz86qukcGgwb+XUxBXmWjIer+CsWBXryFQ2/iJ28Pkw73pPineTb/XsabGhoUHEwMuFZWzxvPofGc5FKIqEN/gn8n5+VVwW6xcE/ARBUmqiwQIKZrpoXO2UlmR6X3O+GzzM2NubMttqePZ99rnvK9cJ6d9mq4JWAbFkWL4Ame+38eRVymDU+fvzIkIKAXUXhLCkLFbpNkiyQH0MohPp7MAtc1Fj0tatXZfRI8c37x+ZtbCL49FmDtXfCtgVA88QRhiUxlHMnMu6J+Txvlzhq8aJXMcUbffysj1pTwDmji6Z2nBxjH8iPATAfWYDA5uP+REDRgWovsONej3HOTam9kcL+ZG3wzNw/xU2hiRv7HhlIZ0jawpveAu9JvmEdcp9bs7a97c3zpaVFsZO4Zm/4U9hkwtngEy29fT3aD8QspHV84iih/cMawJiQ2MWHZ4yaZm9hq+jTNJKgQ4oRE1PPGTY3NzDZcQCCu078asno93crNWtry7mhrChEFAk7Mg3Ed4ICRc3Whpo1NjO6TrFg1tPZEUBWb550491QKgtY3irsyER29vkLFdrIESFXAnCm6TCMIZua9R4UQ9wXNXp88NE1bpkKI9egoSd/Aicmcz2ZlrSdeOm4xuXJDa5fu659ADCKwR77jD/DeCQ3cI8dlyeJurgwE8Vyb8nYr/7jf7DZZ8/t008/tRezL0Khh2k1jZGaJBccWKTR5b4nDuy4ST2fWRNDMsn0JqOYdbmszjmaeDAli4Vt+6N/90ux+GSAuQeI51MjNCUOHjyoswwA388Ypilyilm83uVLl1Q0w+h2rxLWuE/tsmZl8r1X0yQYn0XSZk1N1t/fo/yqta1lnwV+48Yd29mpKvdKJjNWKtMYSlq9ARlNn+4DPAOs5H7CTiXOCZQNxSv5BvFqcuKAnThyRJOzNCrKpZJdvnzR7t69a3/yJ7+yBw8e2e8/+dLGDoxLQgyWa0d3lz168lgTOrnWrJopRw8fs5XVZVuYX5S0TBVJToDD0MRXwz6YX7K+iU0u5wagxCSc77mYt/JcOMPU1FRD0Nnq7B3PvyAUOBPeGxwO9NCYI+bsVpja8rhLvs1kKDFXe115oOehsMs5JynK9UxbW8Ry5rUBsIhVrBP5N0yO28kTL9nuTtHSyaTdv/dAetXf++BHYSpo3bKZpD2YuWWri/P23vcvWEeGScOiteaIBVXLb5bs/v0nVq7Urb9vRKAfUwvbxW2tla4un6yAsQordnO78P+x9x68cV5pvudTZDEXc86USCpLlmzJtiwn2T093X2nw52Lnum5mMUusMAC+9EGi50FBpjb0W7bcpIlK0ukSFHMObOKxSqSxVr8/s85lBfYL3Ab5qCHlkRWvfW+5zznCf9gPb398tWJkp/sC5o1yieKR2o6ZtLEKAbqyNoUxX6lGUNzD5nJVE2lao6OznbJAuLhcvHSa6olnj4bCSwUl9hjb8iL7vBQ+tgt7a2KPetrK5JJwaA2KdNXtNiPNFzr6+2yxtoaNf4WF6essJ+3uupKq+S5pqqsrq7aVmYn1UzqGxi09e09287k7ZPPvhEKvqu31xYWlmWm29PdFZr+CXlfdHZ26QwkX0CXnaaKZCFlyF4l1jtyGWiaR68kMWYTRZudm7PaWqRnt+yXv/w7DV8+/esXaqKWlcLYKeo+cy5wf0Az01jJ7e/a+uaa1gVxB/k0kouI5BQ4jJAHY0KsZierUUswtGWE5MO1MquprFRdw3nAWsfkXYzig0PLMHTnLAUsQ/7PUL26xr0BM2kFThgOzkhGqodmtEv4iF0egAd7u1lrbWlTg5y4Aat9c2tD60T7yxIabsE64t7AwFnf3rZ9ak/iXX29bW5ti1EDA454zkf0+sgRtaWl3HdHjJPH42fBGalhonI7ZND2BF7q7uyyns4W+/TPX1hzY6Vl0nn7p3/+tX1961trbe8W4/LzL760U6eH7dSpQfvP//yT/e53v7bv7963nZ01e/3Ka2K88vkePnhqiyvrlqyo1HNjyEAO/M71t+2727dtbGyCibvkZguiipSoxuOhNDU2yXtrZWlFtTTxBMYS5/fTkWfHzVyXiUQi2Gs6/szaQMaJOAlD+fKl19TIA9TFGcCgjPUGCIRciLPeZXiRo8mqAch5MjQ4LPk2GqdTkzPHDBjisnKB8EV+KQnUo4KkhjxfLtGejAPaOKQ/RhKHvIo1KOYEMqxB8or6lNjG2lOuGpUWAitYTKHgh6U+QKkzOb2m9XrXcyMHvhHzYDXwc+Qz2WzGsul1Gxpot1/94qZtL89asggavNqePxkVW+v6zQ9sH5Db9o7kfl+Mjdv4xEt7/+OPrao2JQahasemJhu9/8h2tjNWV9dkz19MyCOmW4N+gBplYm1xT5+PvbDV9S2rqauzzM6uFQ+O7PqNt6y2EUnavKTBJGldU2ezs4u2uLJmpeWVlsnvawDS09dn9+/fV12Azxa1BxJ3fPZTw6fC2YJU465yKM5/1juDruh3RdP2yVMkylYdBa/HCGjR5W5gtSqXjf2IEmfWao0FZnxsroqBUYZUjvdnyCvICyWpGl5DABmYrQzWrWhtbc6O4JxkLdNU5/wQ+xAZ58pKyTLx7MmFYUMmkg48JL4x8CX/gLXDs7x07pw9unfHrlw4bUvTU/bBjas2NfrEBvq7xSI6e27Y5mbndL5iFl2JPGdltRUL+1ZXnxKjtb0T34dJO33xnCTZrr11zb747Cu7fOmCjY9M2bnTJw2WV6WMpLM2v7RufYNn7NHohL2cX7KWrj5b3dxWE5x8L72zbQP9ffby5aTnUvUNYoJSq7KvAL9so8CBX0IAYh4VEy791NikvQW4tbmlVZKi+JsgZ0o8516Nj40LqMP9I38ivjIYBtzKPcI7gdeGgYAsInGXvhHPj+fF65AnIKPGma26IBjcxwY98YHhMXub8xiwwF6eddet9Ua/g5jB4JXagNeWxG/o1ZHDqHcX5OgEmASUHNYC60SsjBBDYmvHAW4Alw5Vs3BeiNUBM15gzRLlvdSLcYDGUIq1KAleMcaPbGNzI9QwGGZXCCALY4S+Fq/DOcw1sIeU02FoHjzAWKsAPMTwF8vCAbhi0zKMERCuXPeaejKNmTi9ySAPHQ3EI2Ekgm5jDs8zE7g4+FpIGtdnM342JzvePAYJH0fZH//jxzvwP/EdGKqpPr76KN9Dg0fmNjKd9CRSSYAM3diUTE1pnLoZD4yKqOHNhJBNTYAgoDH5JghxOJJoOcXSGRPeEyUJdvS82jrqlLqED4ce14B0TjRn1rQ8RCVRv4J8BtIqPo116ZrYGIs0OR92HOi93aw758mWzD+98QN7gd8lMRG6NNDx6+pSlsk6CrCmtkaJSJwwu2cGCFf3b3AUrAd0DhF+x9HMR2oScVBxIJA0RyQdsgBC23EYBMqkmsMlpWoc0Dzkc0f0cUTl6d6GnwcZGE1oo4QJd5LCIqL2QATSfFNTOOhLywsh4Gw9MQsJeNSW12DglfRW1DuOjSiemxslewONxoybqbsMEdck1C/yMkLQByRwMErmj+6P8coUWxqkAWnIZ4wMDhkNBYkjrbGQ/Ej2JzRiIpoisgJ82BGpgZ5UxYjONbPO4Q9w3TQMaMDAUFGDUGyVI6uqrrAjeRP4AA15D5D48XPXNzVYohRj1rR1dHWrqbEhEysSSGf7aH0HRk80ffMGpB840nsPjAQm8I6EpSgMQzk16A7UIIvMCqH01eR26nYcMrnOPlrTlII0Btq8KRpQrCSEa+sb/lyDUTX3VnJcGu7QQKEIdtQlh7CQF0fEA2dgEAtIbtx4zgeIfr98X4tBEb1JAq2TJppQaNrzjuSiuaR1zT6W3qkzk1xuzDVHj1EDQUIsNs5hRWiNJ5OSY+NeInlVX1urJItEAPSJXuvYVM+bNW0d7TYDgho0RVu71dalrACjorzM1laWrK2lRcZj6EU/GX1pZTTia1O2trklqRZiILGOBEhm1KG5TDzh2fGlxjSIk4BaEVsseFdQiJKUksRFc3rfq359xCCXuCooWSXRJkFCc5jPzxqUSV0wQCSBwqtC0nxiyIA0rNZ6IWGKCGaeLw0K0LvEOqG6qmvU/ORZYy4u9G+QqGPIGOXonM7tEjs8E6EZGawF2j7PMLIl+BxcA1umpcVZRCRyXJ+8UsScYtBaIpkY4h8LmcKRzysT9uCXIcZamcsF+BCOoiUML2DviaGAH4Unu77+OFMOj30tuF58CNjjNGZ4AdCnvT09KohpCLGupe+Mz4vMsz2G0SxhrZG0k5xGuQOtQ14rUH6Ftg9yIy6L4dJAGiwHAzw15dNpyeS4yaUn1Rr6UrAJzeOa9hGtxL0T+y2snZio+mDY9z1nDO/PGcMwPbL02Pdi9sAQIL4Enxqevw8/nQ3C5qZA0TOWXJEDBWh2svb4LsBCMGSWB1HBdfaFoEs6I5OzT0l7zotGYh/IVgom9jKvLw8q9If3D4VQBUnHdXEPeM4YN1eWk+RzLhTsxECf9fb1+tmUKBUCq662Xs1vCiXuJ/eEIpr4zXrm6/AQ0AAyYEghwhJJyc8EmSdMXMurU7a6tW3buzkzUE+HDA+PVMgszi/Y6vKKJOnwnOB8l36t5AG96Y/PAXuBtUjRVZJw+ToNqEKVEZH8B8SmChqEh8EDpk760zL/23e5QuQeOJPkhZQC2QYT5si6u2lYpjWQ5PUZdP/6V7+y6dkZFdE/bNLI/wejRJqBu7uKAWjgw5jQwDv4EYFaozHHPUU+iXwtVevoWK6ffY1MDPcL9LaQxGKE5iWVl2B9iMVY0FCENbK4tGLIcwmQcXikASRxhf3s0kcUn64f7mxY1zOfX5jXgBcAAPGTdVNdDYsgb41BKxrGVDqzZ1PTc5bPFTQEdSNCmAzlatTwfE4Nn7b33ntP5zyIxP/73/8fMX74nOR/rC/2CBItp4eHpVONcfjm+qrNTE/Z6OiIvfvuu0Lrzy8sWSMxI5WS5jJF8/rmhsAt7a2tGnxzVvNF/EI2r7QcWYMSGT3LO4lcM+cebcQGIRExgE26RBlrTQWs9JidOcE18p3BBvuF3FnsU60xmBpJ5aBq8NWmhBSVTKXy6iM1g1kvFNjsRdae6xn7M1NTACk8GDRiewamL7mQDC0xQ8Xc0s97Gi61gIwyO7rHztYoWkt7h3SrMxk8usxy6S2rKEvY229etMTRnrW0tGhYUV3fYIsLq/bFF7dtYGDYRkZe2uDQoO4X5r08c3JPWBFLK8sCOG1s7NjyyqrOaa6R+8tweXtrU7GAmEyjhMEkckzEA/ZLVWCveOxggJWTzCP7iGEBDRPiFJ+5rbVdZwDxj89DjI2xN4H3hqRVnWlTgpwkUj6wdMjPYGNnMnbu1KDt7e7YxXOn7NIbF+2bzz6z0mLBauWBkrCuzlaxIDg7YAElSqtseWXL7tx9bGWVVVZeXWmrK+uKkRgLU3spXyRnSXrD45hxE66B9YC3CzUYMX1malrAi9jEx0gckAZMkP7eTvvVb36l/fjHP/3FZmfnJB2D1CgxgLNUA372e3OjZfNZ29xBsqvS75PAUi6zqplwYHCzlmCeOWDM6x6xX9E5L/OBbj6bVTxjnXHuLy86+hjQCllOFt8YzjVytMKRzM1rqqrlnYWxNUMFhi6sdz0XUNlBKrCoIZ+fa+Wlvl8Uw6ppeldr4ID0EpJ4sOR5X3n2wQ4k10/V2uLKim2lt+1QvkmwAohLZn393Q5cK/DJSm0v5wwiroH6bxemijzmShzghJSahumHdvbUKWusT9k3X31jLU3s74z9H//n/26f/PETS6Wa5Z3y2Rff2NkzQ0Kq//73f7F/ZlBx53vb2dmw/F7ezp0/Y9euvWHffnNHwBhKj+X1dXkQvX39uiVLEvbo4QPdswrJybBWywxstTwGAb0Emd5sJutekHuOwAagBKMier2xJ5RnqtZ3DztnVzlb96hwYFcuv6YG78L8nP4OKR2GaA8ePHxVkwKq4uGrljsS6+78ufMaVFTV1MiInjPUWXTeG4i1Go0+8lT3xXLZSUAo5J3at/FMBVWfxHvG2ai+Xx3opnUR1AkclOgMZ/Uh5N/hkrisE8+NAIY5gpu+B3vZmak+iBNwL+wvEPw93R22trphFbBy21pseWHWhk+22X/56Xu2Nj9pdrgvQNjUxLRY9Rdff03If3xZmhoa7fnz5zY+MSUZtoEzpyyXdqkfOv3Pn45YWXm1jIqXV9esvKJaORyN0e2NNavDu2FrU/FdHnnJcjvYy1s2nbb+gV6rqKmykbFR5UPkvc0tbZIjnpiatmz+0PYBkVXVyEvLPe7ctBt0O3ktOSLnPOcTTOXR0VGt9ba2duWpMKGpd8SsLknYwuKSjY9PaDhBTHOmqcvEkofx7Hg2ACQ4y2L8khRWqMc9lw1gNnly45cD8476xeOJ53BId7r0KQEIYAFyTtRNPFfOntraetva2tTrMbQkH6X24zteko3NTcrvtzZhawR2uWTFyu382dP29ME9u3LhjC3NvLSb775lz+7dluk9/n2Xr5xTvllTE6RgK5BShYUFCwRW6Yp1dbXak2djdu3t1216Zlr38M7tu3bm1Cl7+nDCLl86bQuLyxqK0qda28pYW/cJe/BszCbnV6y1t9+W1jYUk8ipAbIyXGCgwF6DDYc0nfoUYSDLd/nlhRqCgfL0zJyeGWcj5ztm2gy8h4eHwvOtVm0H6559FhlEAscFSU6XVk44qFFsbnwjnDHFeUsfgxjjHg9u4uwycZ4Tq18ntkGVck/VZBpM7Ckv1HAhSG87O79EuYxANZIP8zUhWVfULULdxDpgWBN9XVUv/nBQEekEQaVEcaqlReuJ15WEJObzWbz8nH1FHCEONDTUKe5y3QDINmE0hdwJ6TryZzHZ2UeVFfI+4nyN/RYNQCTN62sW+VXqRPeRdD8j7jHrG1APn1lm3ykfCCHxxXWI3RGGD69GMA7s9FanA41c9tZ9ufT3AdgdhxM/Dir+J27I/3jp//934FxjozZTPJgJQJJkCLSkiDJiR0SzYpJ3DjUKPPZIZiftkk4kjASwkBRQvFOQgQpTASoXew9EfMXkkwaDdLeRBlAQc4kXbWghJpziJIbFgTeeY9OGzUmxz5cQnCom8sdIVzWpFdBdP47GoppohcgsOLJkKchBbwQ626NcDU41QctKdfAWzafNHDTQ6PisagAFY28OfwVaNaZdMztVl1KCHtEBESWnxEvNjZwSeZJokL8cCEx6+RwEdqHiqqs1PY8yUVEqhIRBbIOAiI80bE3Hg0+Fkk6ZufoggMqaex3ZFKJw03iMXiOBcRKTNa5DQk4MkoTypMngGsueGAbdUDXj3McCjX9HpUTtQEdP6yDS+yXEYDj2npBGNfIRr5JNGpyRbQOtXKVQaNa5lI37bkSEfUwsHVXPUMARxJ5o0zh3pUP93PH/C3IQar1S/Pt1Sac0SPRw2DpCtlSNbg5xIUAxvRXimWYwngJHShZ3MmlJQCB1wHoBz8V6pcHBM+Bg1B4R8tElUEjO+RK9kqFfQLzquQQ5LPeeoJhD2sOTAZnCB4RQHCzEg1PJt2TLfFDG+7JPQZ3IiDx4U0jzmoM06N1rGBY08OPrRw8K1o2kt9Rgdy1afp+fI5F0c2FQrd441TCNxmgwA48NUZ6EN7zdi8RlXny4SOaLdAUJp2ia+OOEhrSvVZ5ZQlRYGj+sQ+KQN7qdCUCtRHMLVM35s2cle6A1UFJiE2PP1SSfm5/TPaHxjezDfs7lZtAc7emGVbCtgcVeBuRitc3NL1oGjf5Ure3x3IIsHglYNDAXwpznuI1RbkHIFbGiRIsP8iNBjkPSNEIjugE1a47YyE9pUKb9yrDW/577KEYDCSFyDPK5MMUIHwYhd8Ua8SYWSBFf/47i0DAq54mfUEYMSUV737PVtVUvHvVcyo69DWiS4FUh42MSRIa/xM4gw0EDTB4W8oKgMPXYDkI+onCUHAY0MwUSMhYb65thfXBeeMPnFdXeh5UqmIOGrWJp2MuRRSVNWwZAAeHPs9dnTfq6I27RbKPpU11TpSSQvUbhRwEP64Ezir9DqsgTQM43Ghp1KqK5wdC61SQ5OBDCjD/DiCI+OWqwUkUEX3hpxIaKNJeDx0S85sjyIjkVO0tIMtdnjUizKMGivRESfy8CHVHGvXJjOD8Dtd9BVYdhuKOaGMi0KFFmXzDA8/3oMTnuN+4ZAwIGMjBOaKBT6EoehjMc6cCAMKT5BypbTC4avsQvIZB86MvaQtOeooLiRFItSIBVohHv3glQ3uPvMbxVAr+Xt/LKsL73HP0OK6lwuK/hRE9Ph42NPpOfgA8DnaUJ6hLJGZpt7ufhTBKuHUkfmeUxRC09tOwuUksY8R1aW1uz9kmSOEzhnc7Z2s6uHSXKrKSswtK7eQOZBnuC3TMzOS0qOPkNEg00FcgF2lqRmQH9uam4g3Y4FHHit8v3OUM0ykt44ZXT2uOF2TfomVMEYfa8E3TvKZJoMks67ODQtja3hArDzFJm0KDQkKgMEjj9JwbEfFheWpY/GEMUzkeBQfRc8s5maGsNTMcjq6x2ND/XSdFFnCWNWFlbFnL49OkhOzk0pGeGETFDJS6aZ7extalGL3IWlclysbq4HpDSYp2mM86uDQNKGsRd3d3Km8i3GOzy725O6d5TrFNJWxZ9SEicY52DYMWkcWNzTbkUw46hwTM2+nzCHjx+JuNQBi0wBhubyJ/SdnRIs7NDBSpNJc4szCTliRWeAUGWwSlo12tvvKHid2Z60tpbW9TwfzE+blevXpbJ6JNnz62T669Dozgv4+aVtTWxe1qbmyX/V9g/VMznWW/vpK2i2u8bcicC4xR9cM/9pPkZzwuXfPSi06VuQAU7I9C11I+EkKUpzb7g3imvs8TxEEv5qfJUBnwOHnI5Uh/4R0NTQAseYxkehxwiGD4KWBNYxzzLmEOwpp0JtWI/+fAdO9Hfa3OzM4pzIHbLdTajW71puVzWypMJy2xvmh3m7eOfvmuVhgcXjI2kJWC2ZQ/s3v0nVlffatPTi9bS2qbhHkMyMU328kJ8q8Av4h2QVWMEE2jOGAYisGC0j4L83OzcvPY/z5rXEwoTU+pUjTwNaPggo9HV0REYUDk1RbiP6PXToBezGaNZeWQ5Y5WvTBbEf0LncaqaOMbAl/y5QjI7AkWUJa22usLKS83aWxrtzTevqCaaHB+zhblp6ZxjMl6bqtLAhSZjeidvs7Mr9vjRmO0fFe3Slcv2zbffWUNDkzz8YJ+wzwEhwPaDYUhzSR4VnAEVmIHuijUkc9rDI9vb3bXyCpeJpWm+u7crn639XNZ6ezrt5z//uV7397//gy0scU65Fx7DGfYF64XnzQAyu5+13TxSv+LYaW2Sn6sewVMq5ArEfiSGoiegJ/xHQUrNdcJhHrmcUpmtr66pFmpuahLIJZ1Dgsksz1CV+i54VuFU7b58jqg9Svj55qa7UdicvCPI9UqyBNS8n/0MJRhy0DgmbxKTsqJSQxV5V4F2RQqSoTgeMdvIOxbsQKwRapCEzglqMmTOIBpvb8O29yqC8zPNwC4MKjxXK1g9zeTttL197bL193bZrc+/0DPgs/wv//pP9uWXt62+vl0x6a+ff2lnzgxpkPunP39m//TbX9u972GebQvERhPsF//wM/vq1jeSc8nm9qExiznB0IDm6v379/RMS7gPh0XbzR0IqEIOxJlOboLqwYvn42r6cZ2nTp3SmUPTXJhAahhkjQ/JH0M9F7wF2Ud8VnLJt9+6JvYeNQp1OLlt/8CA3b79nfauQBYCVgRDddg2GBWfO2fzCwvaM1OT0w4mQX5rd0+5hdfOiSDf6N4S5BlcV6yDYq0sD43gRyaQZNinxEn6BpLhDJ6a7G/V2oHlSk1OXFUNDbDl4MD9bvhdajmZzyMbGOrk0PQUiC9hlqqmwVstaUfiZ2tLk2W21+218yfs5ntv2MrMhB0d5Kw+VW8vJ6Zsf79gV997S89hLw1Tot5Gnjy1sRcv7a13rktukgG1JI/Kyu3p46dWOEpadv/IXk4uWrIMJhFyijVGtXZq6KQ11qXk85U/KFh3T58tzc9bW3OT9fb3iB06uzAvUCNDCvbtytqmjU1MWllVjdU1t6hu4fPzfqwRGZgHnynuB6h9zmFnSB9K2nt6ZkYSiN09Xcr9R0dGbODECUkc3v7ujvZgLg8rApY+tYMDiATeCPmpei2hH+E5rbNUFHeCoTEXxp8FemG4yTBD0sxBWSP4VLCX29qalHdRm/PvXB9STNEwmXVDLtRY3xgkAvEgq9SAW0yKHK/PUIW6o8xODw/ayKMH9vrFs7Y8O2kfvfeWTY48tsETPTYxMWUXL50Wg7C5qUXgvvpamKKl7plTONAAoqmp1p48Hrd33r9qE5NTdubcaXv88LGdHhqyibEpu3ThvI2Ojltza5ttbm/Z6mbWTpw+a3dlpr1h7X39Nre4Yg0tzWKOcW4xlEeiqbenT4ADmutIl6oul3IEQDGksxyoxzB1dnbe2jo6dC+Q+IYFMzU1LaYuMlbkzNSTU5NTnn+FXJ5YQbuA/SPGZuiZ8Wfk2qidyUMl71ZwMBRsSOVUfI+S8QGoxV4UMA35v9BUZ28TE3wg6YNC6g7vzfl+J/cQK7y8wv1uAZbQV5ME/KGG2KxNfb6g8qJj6hWZwD1yQr8FZr7UYnI5DelY2/JKRNIpt6d8k5qYfx8aHFIuzNojL+C6qSMEEsz7oEWDUAasRQcLcS5HgJXWsPo3zuLTYCUMy5AQjJ+fwbHYy/K/rFUchL0hxRjAAKG2P26fUdeG4amAuoFxwvXHvaRY+gNL7R8HFb4mfvz6G7oDlzSx9aKExg8HBQUExSyT5Ihsr8cQjWQPI8T1AAAgAElEQVQSFNv+vhC9bFSSexkjBjQWhx0HlhI4gmiQqyDhESUKlCBJTZAGclkovBJA8nsyoukjhZ4SBd/0r1gE3sSKf69p/ZEjO3lNIdcqXUebwkVDAnT5g6EPAZ/PAAMESiaJFChKClZek4Oc5j+mqwQQKNFK2PYo4qCi0WA9VFPaEQOhIaEGvKN9eQ+SX4p8xxs56oBrQX8SCi1JuAYu3HeYJyA9KhzBrsOCRhqBjwHRHs0Cb144G4LiD2kLR+uK0UHyFhL6KKV0LHkVmAC8Fpr3FBeR2k9DPN5bl1ByXcho7OyIUGe66LtkmV7Rdn3aGw2tHYET0RIuJ+WICgoNNfeZlFO8QKMFhatGqh+2/rMYKR3qGl2D75hA46XQkd+HiMr2IZubi0eEjqTBQsKtgB/0VUVRjSebDgAfPnBdVTCIrCj0HH/P+RfR0RyQajxhhKvEFqkFtCKD4d7RoZWW80zLpb1YVlElqjgDi+0dtE+ZxpO8V0hWIR6ksbHprAqflsemLQWo6LKggA4xlyu4eWtJQkkjX9JvDcZxcTgQG5wyWJYRNjIuKaFPeH2KDZBrJKpC5IcCz5kVbvCtgz8UESoCZfJeZklo5khNcR+UNDkCKRoeiqZN4oGmsNDVjuT3zxvYP8Ew3RHxXhhwDSA1aUhEMzxen6RAzxuUBXszaL+zx9nPQn6COFVzH+kkmC8wkaIMgGt+Li8uSppma3PHyiqS1tzSLJYD0hGLS5tK+GEx0PiCUt3e2mg//clHetYgwZ48HbUkMZLkZW9PjVkQg3xeYggNFQp/inAQmnwuYhgyJt6IclrzztaW7i/XjqQGnzcaB3N/XNvVhwbcH16DZwYKQw1vIdxrhAziv4lRNBtpvJH0kDxSANGclLyL5M+csioWRSjuuCaSL6S4iJkxzrJ2hBgPBmgaroGITtUqcWRPsRZhoHC9FAl8NphpoE5I7Gjo83qcIdCd5WWQz8urB38KNeQ06AzoOeRvuruDvwcGqjTi3ZdI7BKtJY/3jposVYOdYpkvmrFIX8QhS9xTGlbg81Pueq3cc5574qgoGQjuMYhmEnC+WAvO0PJBjwqnVMplCSsrhSjkPRlWsGZ5Pa4lsiHEGvtBHNTaJOaH4jdK8/F63A8+l6OgX+17Pl88C/gcDZJI2pHWNPfi8ePHel/tMw3uPXHlOYmyHIYb/Bt7lKE8zySaWJOQH/tlwJRRE+pIMiugQTu7Om1qZt66u9rVjCHOIDXGOpQOdPDLiKjjOOAgEW9sbFHSLe+JsgoNS6CqE3NlVnlwYJtb3Hf3momDdW/mE5e9OYXkRGNjnZ0c6LNrV1+3b766ZS3NDY7IZ96YLBXrh4EXbKeTJ04K9YqMGfJBnKEUpfSHK5Jm3R011tnZal09ndbd321lFWW2h+TbYdEWVjcsu1+0QqLcDoulMkOmaEL2Sb5SFY5k28/mbXx0TPtoT4wl2Bn1ikkvJ18qPrIOHBgAE49hvhfrnHHS3pYxn6NAXWc+rcaC/IQwnKWBt5+3jvYO5V433n1PudXdu98pNxk4MSB5EvYXr/Fv//Zv3ngIflfsQ1CGyBXAAKQgHh4eti+/+FrSZa9dOm+PHz9SnIgynVevXbPHD5/Y6vqyNTal7L33P5AWL+cCEjwgQyU1gywGZwlsoN20jT17bsliiZroPG/lhiDxZfyLjKIPATVMlqTlke47Q4U4uBO7I+QycYjPvmJwByuOgfHw8Emhq5HxIOb29Q/aYSFhf/rLX4VSQxpqd49GEGw4L2TrauskbYfROPGGe480X19fj86jjfU1eeDArFqaX7T//rvf2YP738uXiLzt5cSEnT49rHiJOWVNba1QtDvprDSkZ+cXJPnDkIL3o6EAq4XClftFI5nvrHexMosF9x7TsA8GC95hbhrLF39PrCQmSodbMQN/tUoHawTTYp65JFVzzq5gj7/xxhta8xTt/Jl7541T03XJM07sX/ep8Hjq/m2c9bwHz5RnyN9zvTwz3offFQOkcCCU6dWrr9n8zKzd+vyWra9nbOjMEGNq6z9xwv2QshnLZ9OW3l6zc8O91j/QoYG/0JWpWht9PmXffPPQOru77P6DSXv/vbdsO7Mj9CcNAuoAmvXEP8Ae+4fIRaUtVVenc5R1hGk1+Ud9XZ2QsjAbaSaRE2EuC/OHoRF5AMMFwAqZ9LbQw6AOOWu5vwxTGXZzNrAe8edhfXEWAo5YXFyyIgzMMtfax6gACRzWUp7cRzr5lZbNpq21scE62pqsrane+jpalH/0nT1j6ZVFu3Xrr1ZbV22NDXW6ps6ObqsoT9nE+KyNPHth6Vze2rq67SVN3Opqq6yq1v0v0dkIG9kRtMRFGhM0k3m2xAeGNYAsOE8YBMa4R9zCs4dBKAMkGuj/+I//1XYze/af/+MPyk9raxtkVO4ebt4gAmjA89473LftTNpBOOQMsDP38ZNxoAgMM5pkyudhBIc8jdpDfm2lCeXSOp8Cg519wl6kAcQwlqFUEbm1QsG2QLxKThLGsDeUYUWwn2C5IqlKfs/n5N+jhBugG+XLpaXBM67RzxCGVVxfAgY7w2HYeTSdnFUGcIg8gLUFs47rz2R3LR9AIRUV+IildU/xQnKcDYOXpBrCGPnGJj+oGGRLGVTUVFfa7s6e3Xj7Nfv445uW3tqwr259bpMTs/ab3/zc7t59aK2tPfK5+eunt2z4zJB1d3Xbnz+9Zb/9b79UbF6YmxPIBgmtDz/8wO59f99m5uZsK7NvR+aNL4bW199+2z795C82PbNouX1XPDhwmXoHDpUmdU68de2a/eXPf9Gz5My9+vob+nd5VNBQlqO6D0yJW5znNHEFiBKjB+nDvN28+ZFNvBgTwIPn3tLSZj09vXbv/r0A2sETqMwOlIfTaETSM2mDJ0/4kMfwTBgXYNGZj25ay2txdu7lsgIfEOedoYtkrdfvkZ3P2aD9ieyqgGslxwM8eg/EK+KX5L1yfibBqlbDvMR/NnoEscdpdCPbI7BPAE4pbwoekhG4Sf3e29Ot611cWFLuRZOaHOGda6fsg+uv2dLMhBUP81ZbXWfPR1+IBfPex+86aDGXs4amFpscG9PQ6fIbb1htY6PtoIVP7VRWrjM4X0hYQ2unPX323Da3kdThd/eN8dzpoX7r7+60hYUFAdbw7dlBkq+vW/5BsIJYm4sw+Tc3lSclkxVWUV1rC2trtpvft/3DgsyVnz4ZUX57+fIl5Sr3H9y3vVzBPr75nk28nLLJqRnr6WqzS5cu2Z27dyV3d+PGm8p3PvnkMzs5NKDm+WdffOWsZlgVkrahf+RMcnor3D/FW+ozzqzApFAPIQDO3OvMcz/WD4whnpEDzoh/vr/Z5xqSyoenUexJB60CejhQfhsBDuTBDhADnFKwUnpJ8grIW2ZnxzKZPatvqNWAl3MOZuXzJ4/s6qVztjgzYR/eeNMWXo7a6eEBe/58zC5eOmtPnjyzjrZOe/78pbVocM7+qlfMXd3e0lkzPTFpQ2dO29OREZ2V392+Z6+/dsGmJ2ftwrlzNv7ipTV3dNrU5KRlcoc2MHTObt9/bEubGWvvG7DJ2XnrwHx+N6PzEOYI/bfunh6XRUOdQ+DGUg3jY1M75lMMjGC0dgT5Xu6d8vmpaevt7bHpqenjof8C3mL+FI5BtMR0H+Z5bKeu4j1dNjgh8AUhpquzQ3+m1mRQQ21FfHZvT2cKeM1P/6RasWB5ecXa2tukWqHaM4BweT9k9xiokA/70NCfN/VmCecJQw9AHVKDQAbTJd15xv8fRoV/nKDW4twCcrTY5GfVAdoCLMSaIQfwPMpZ0q3NLQJh0NfkrOIDSKlhY0MyelKyoD6MbNdUSqAdWNDIApP/qlYMUr0O5Aqev+QL5eXKvWFrSDbczOqU/+e9BtAACG8zV5gJ0jKKdd5P81yA1ySHIcaJ5RHYKZJ+jk/1R+mnVzfjx//627gDVzra1WTjgCCIaMOF4QNotNg44aBwCphvvsb6BhUMJHQkBLExgqZsGRIHNKnVxKe5WmqrKytqqnnTErQfxW9s4PskV8hSmZKC5AkBLVAEY1CNDIZomi3qW0BluIyGy0XR3I86iQQ1ClMGMby/TCfVOHbDRSi+boidVNOAoiLq8IOy8eCac7R5MBqO+u0RaSq5HtCdAUFAYU6AcaS869zx5R4D3oSLjWkh6kDTRQPx0FBUoIPCKvSWa5VzKkjageZ1kAvhdcUm2HefgmO2yQ+knAj23DMQaSCg4/WI3hwCYKTTRsaLhiuByuv3DcI26CVvcLrckwdWyQYpGQHt5GagkUmiYRfNCoyvgla6CqRozgfaLzBmfDDihxUJrij5AQnI5+T9aVLEIj6aqnGokJyQzLg0gZtzi+576EWoEDIBmeUNPjwWYBsUj9kS0JdZTwwsSGh5piTfuscMqkAZIA+jA2bP0Y+YowZ6JMMKkkKkU9CW5VDmvfz6HJntB4ybmceGMoVZ9FDxgU1EHEUTbV8v8dmwRyN6QAOvgEYI57XOOT4qr0mio4EAjJdAu1ZCSCMxDKB8IOQHvNZ2QDjw80I7BFq1s1l8WMgTishYmq9x2ESDP5rBxiGaXg8ztR9eJ68dmDE6nANyhteJAzvJaFAEyQcnsGiErPJGC3tZvhml7s9SiTYt2tiSkzkIezpnV69dVeL8fGzMkuhygsTcWBdFujThXgZ1DcgwuZdFV3un0IGYP965e0+GdJWplL7TmCUxlpePhiYpNYD5b5CvNKD54s8+bIm0WJqxLgOkIVRgWgDXI8bEz80+pvGoARr02eBxEe+1Gs80KwKaUAw2pL4kQcfAzIdqWkNIewTjVl9rLoEiA7bQfDweIoX7z79HlCXf19bXFOcp7vicky8n9d+nTp22ly9fCuEEE6yvt0808ampKSX0p06fsbvf39PwBNM0mlEM7sT6oiCUvETCWpqbNexhL4vVFoxi1cxGN1xSF+77wD7mg7E32VsxdvlAw+NObMjFZiGrWgMhEHflFWp8sa5p5umeiJ7r68nXreuQqsFOQixmmTPE/Nzyc8bjne9PN0F35pcKrzAo4tnwWSn0aFRyjvig3hGLxMHoHRL3Comr05OD6Xw0bA+DTOKHhkYHLisYxexEPQ4eQDoDAuvqmJ3xA7+LSNHn3Lt69Q3dC7w+eG5ff/tN2H801V2CSJ4cJW4MHgetxzJ+paVqtO9gOA+9/eBQ/2P4QUNWvhcqFNZ0BjN8gdHkMlQ0UT3GsF9pPnOGbEsyocpqqirs3NnT0hnfQToxsyuGIc9+fXVD6G6MKH0Qi9QXBq95q6urstrKUrt49pR05S1Jw29fKK0DmuqFI1tY27aCIZlRbolkhZWWIdvjSLADmauWWzadcZTg3r7Q8xgKw7RiKMkzfvzkkftwBHq2FxO+v1lYNFjJDdjb+rw0hmAPMuRSbhRZKqB3CzY4OHjMQuF1YBTsZnbch0qm5qxJ1+OWxBaGvqDdAtoUBhGSSayzvv5eMYYESsCcHEPbjQ1n2qyt6exC7gnmHffs6ptvyjsA5DYyWBSn7D/QeSrsVFhu2vzMnOUyrsvLZ/C45PJX5G3REPqAYQISOAxyCs6kcPRtUShaPhNxBdQ+jUf+XYCSXF6Mir0whCBm8rogi5eW1uzs2YtWVlaJQKi1tjbZTmbbZmdndK95bZgI6B7js8LnRvKN+E4DZfDkSTVUQHePjz5XQ25ne8sunT9nudyu5E2IY/jY7OUPVIgCCFleWZcMFCaiKytrNniyX3Gkr69XjdLV1Q3FJOK/pHVADCbJjfBPcDk3Hzx7PsMXf07vMGip09pw02tkT3iNSj0vnpX8LCQJ4Hkya4nzu3+gX7EXeSCYODRyiSsgf+XnFmQ5Of/lZZV3ZlkBNh7goiAFRozv6OxQI1LDCxqUgUELS+IffvaRDZ7oVe6ztrIqA2tLJK29s9cqa1LKT2cmJ+wgv2s1FUk7c7bf9tNrVp0iZh8KuJHO5Oz+gxFraGy3dJpBREHIdrEuhEQsqrk4PTMrZgU5KrJRnBHK+S3hEg2wqhjWHrIWtyzLn2vrbHUVOZB6NZGQQULuCnPjb775xr3kAusXTWwNwY8KkslYWV7RPmDYTrOkr7/Pvv/+niXLKyWnw/pAQormP4Nr5Ux4mom1t2sVZSUgl+z9G9fszIl+sTbR86+pQ17x0B4+vGttrR4rGuoaraayzp6PTNrLl3N2mEjaVtbPNj4HUkdibBwWlDfspHeC0WzIN8rccJszlHsSB51uXA3jjnUB+4sBNLI4RRs60WG/+uUvbX1907786ltbW99S/gwggPulswZ/goRpDaVhYhQwL/ezxCVCQNa615/QtsGfggGqQCs0SwRy4EzOWlU4Z4j/rGvuOcNlBssD/f2KAdu7GdtjSAC7q4xmpnsdUFfKeFWFQFGALIYExBm+eL6RzRjzJM4asU73slYrb6UdNc6QoUP6ieYl8lDOjnY5EwY9vAf7lXtfBERVwNOgoME477GfPzA7on7wukEs7qSDtsj3ZcSdRP6Jfr+bdZw5NaS90txYr3xyavy5Gt3/8R9/sN6+Ya2DL259Y4NDA9bW3mGff/md/ctvf22ff35LPiScNTAbf/p3N+3OnTs2Ojah+4vXHTr5nV0d9sH779qtLz63qak5gbqKDI+Q5yoxy+HLUl0jZuhrFy/ZH//wJ4HteM4XL17Sfnzy9IkDCDWo8OG8hkFCsCN/Re6h268hwo3r1xVfOftYC/gn0GR7+mxUdaQYn5JYPVDOjPQXMqrDQ0Oqf5HBgx3IcyTu0NaWvxN5vvYR/mfODNPZBoDiWDrxVUx02WFvrhITHbhELRy8rIJsFfGUBqrWIj4XrDHOYwHxaALCQHNZKQ1jj4pis0TpadWMkuCjP8DZV2HdXZ0aoNJMbG5osOWFBbv5/iV76+p5W5+btEMQ2qXl9uzZuOUODuyjn32kz5XPMqhospWFBfkC9Q8OWmVDo20uLwtAlt/N2sOHj62sut6S1bX2+Nmo7eUAaSExdCAUfWdLi2qazY0d6+nttIb6JistKdqJ3i5raWu1rfSOvJGIkg4OStr2zq41trbaHz79zBZXN2xw+KQNDpywb76+Le/ED967rjPhu9t3dB9vfvShjY4+FwORwf9rl16z75AjS6ftxo23dZ8++/yWdXV12Nmz5+yrr79VriDWvEq3hGIWccdzAheKE2gzoMX58zHwMbB12bvEZ8lmK9+OdZ3XxpxD5BMMFwWCIZcrukxx7E3RDGfQ5TJf7kXqsqP7YkEi3Yg8KCxbLXSGIIUjMfMHents/Nlju3b5vM1PvrD3r1+1scf37LULXttcef2SfKvaO7ptfOSFtbS02kG+qGFHSWlReVRLS6NiW9fwkE2Nj9u5C6ftL3+8bVffGLbJFzN29cplgR5aO7tsZnbWLFlhtU0d9u29R7a2s2cdfSdsYmbOenr7NKhwqbEusZBcrgsGuQNY+a6qIKigiLGAafz+gS0uLFtPb69twVA1E0sGDxIAK0iv1tcDcjnUWUnOpsGEWNYOEGVv0fcgl5YnYmAHEOPVG2NorPylKO8wAXGCbw33OnqoRlAkeR/vIw/OnLP/WfP0TVgIvG/8Pa9lABh7rUytiCn1kUCHziZ32Ul6NQ6W9H5Q7Fq8UvWOoIsoEc36kHcJjNYAlCJuER+4JvqSDAx5XQeXeD9NPjYNjZJmir5xOhODtPvqypoY+2LqSao4MoU8v3PPRj6r1zcM7BlC0Tflz/IRzO0p9jiTDBCeqxeopgv1uGo57kuQwXbjcQdnxq4NzMPjIeCPg4q/jeb8j5/i1R04SXDA0Cxo35MwoPcKWpaApiIzTDPdl8A9DOpStWqAkjgj9cEmBaUEoslRYTRgfFJO8IGd4AVJdKoPUjwhIXGdvGiIDBobXU3X9ZUueEA9RAS/pGAC0pY62enzNI8cmakJrH7Hm/sU2kp0odAVveiLwxAaCQQKXWvwWgB9Q4MbHULeEwSnzEb1GbdcFsPbV66BCTMiFOm8tt5HjVzxPxRO1cAJSBV+Xv4NJclg+OPNXX4+ItElQxQb8EGDU0nU/r6CKMkrrytEbQiKknEJNAShfNX9dTYEuZoa3KE54kyWoMmpT/TqmUhDPgyJXlHPKF7c30INh2BkLkkaCmM1U/xAVYKCTFfQUvRAXrQKtH8peAzkFablXowcSw0FmRJPPsuE/IpJK1dIYSEDuJBskJwwlabxFYddQpyFRMWv0Vt5FF80qF3znqaBD6cc1fFKHMpNtZng+wHO4SpJFCXiaEbv6fecjn6kaThoN96fYrM0Wa61QeLvSk38Ls19ZIkaj4cBcU3zTKLWvdgn3AMVRz6oiugJDkkd5MGbJaIpfvh89Gy99gjyWAklLI7mxbj6UHRtmiwRLUtjwjUYff1pGCZvZr8vLg3kRaLWdZAmkk8ImucBoamkJ6I9wr6j6CB51FoLFEbQCcfyPoFp4g0sf/+YrMinwFy2Q4lSMAznfSiMJJ9FfAqFiBDs+znr6WyXHiRMCoZh6FQPDZ+SJEhZZbkaUAvLy0I4edPP5aYqa6pEu60oT1qWRlyyzFqammx5dVXNiYKVWB7TsSSD2MAGCTJXDKiIQcRC5I7kdxLoqa6Q4yha/rO3D5QMGtOlQpywQjS0pLkdWEjIDshPQSbWvt9iMcda4V7yeYnTLnXmzXgaFbGRie41z1w68zU10roHXbyyCqq40QZODghtCsWb+Hjq1LAYJKwN0EJXLl9W4ULCDrofTWUQOjQBQavw85hZ8/s0btmDNLVdQgTmSouSQ14PFgSfHc1rxSf1/WlSMfjxwZQk/0o9vhCb+cygVmInnuTSC0gYKmh6YyqHbq7L0fG6Ml7FkwOfmcBUi2eFGCUMyYNBOc/AvR2cseQNQ+IjuufIHHjclHBckBukKceaJFGkUaIENlw/7yNZnRLXeWadx70jRh7arzU1YjqoWbMNirAsDF/dqyaeb3HI64WE3ye+eP04xNP7UEzDdgjGpuwFR6gH4+nAGDseLgavHJd48vfr7+8TisglE91Dgrmhzn3Jt3mBEIeUrktL0yAguxIm/V15q2C8FxpHFAVqIkneq0R61f7lkoSSCYJJVU4sdQADRStIXM7v6mo3Zz1/9oy1d7bb2PikzS/Mib15+tSwPXn01IpHCTt5YljxEjZBbi9jVTUlNtDfZSe6O6yxoVafh32fzmbEjNorHNn6Tsb2Ds1yhwkrlpRLH5pP6c/XrATmHYCAnGuclyeSYlPM4o+RqtP5hffPi8kJNS9c+o5ChwFC2PvBSwtZBIaWQpzh5yRPn3i2R8NP8p09FeQMPpF0omghHiHB5kgyJC04P31doiPMdxgU9XX4axFXWZOgv5yBxTMmr0FmhDXJELGnp1vNTpDkoBhpuj9+/EDnFuyBVG29HGX3so70Ei2dBkQAU3AGLs0vO/IuyHvCVKRgBjHNEIDPQFOXJiHXQmFLU91Znn4PdLaEpjhxkOYS+14SgOVl1tzcaLtZR2e2t3fY0vKaLS+v2Y13b1p9Q6ONvRgzjBAHBvrs4DAn9C77gJzK96uvUWLKYZBVEtKb/O+wYItzCzY5MWGb62v25rU3NBCafDlhb7zxugY9z8fHrb2jUwUkcSsHwvfI5H0BC8xp+kjTwFBgCAPri58p6gxggJRJb+n+RS8mroc14nuvVENchjWSYTlEgtCb6C4N5R5A7F2uxwvhwC7TEL5MA2Oak/IcEfNOwhDHchvsQc5IPjNrg4a8M2qcyerxzuUaiSNC7AXJRhX3Wxv2kw/ftrOnh9T8RwJtcmrW0qD5aeKG55hjbyH7eZizKxcHrT6VVP5eQnO9otompubs0WPOkSabeLmkxtns/JxkKYi1sCMYVCAlhXY7cdWZisiKYDC6Y50d7TLopEnqUn15rWMBYDB+RQ6kANvNGbA0Xcaej7nJL/4CNTXOWC0eGbIQqVSdLS4sKPeHJcgXcZN1uLWza3t5R5gSg5iPw6bQGS2gAc/nwGrwRwGhfPGMDFnzu7syVydO95zss2R5iT17eM/q6mutv2fAKspr7NmjMVtYWLOSylo7Kk3a+uaWrWMiX15hTS0tNr+4qOtl/RM3OJdo4JFb0DD1plOdztT1dVDh+1ZTzYD3yHq6um3wRJ+uWf6ahUMNofGccg8MBiAZezYyYplMNphgO4BsEKmSqSlbF/OzPOT0LgnpADGXexLQ66hg1WL9EL/L1FiCDUejrb7WmfYCoQSTbGICA2qxGvBSIq8vK7Hd3L5MxZ30jVyUN3yUgZbSvHQdbmFMQ72ngbwQpoENrhrTaytiIvfO17APzCvLkTYJABv9aqgfgoyp8oIScjCaZWWSfgK9LLafJS2dQXbTa9rSMvxknCVGvMYcW/Q98o2ypHxv6lJl9uTxc3v/xhUbHh4UKvje7btWUsqQPm0PHz+1gYEBq0nV2t17T+1/+19/Z3/506eW3tnS3iVP/eCDG2JQvpicsj28IQ8KBgu4q6vTblx/27795hubmp62wlHCDosAVZAkObTDowMN2BlQc0Z+/tfPj5vFZ8+e13McGR1xj0U1t4kFPjCgKlMiGcykyQU4fz54730bG3vuJsUHh9bV1W2NTY326OFjMW4FoEq4v1gdeWZXp2Uzaevq7pLXD5KQ83MLkusDaBAbdxFQIs8JyTB5HoMUGHXKMdtXMp0+KIsMcpeZcganJVy6k2fuoL8D5dXyiCT/oVmq+tmboxFYAgMwym2yfsVeCuxt9370Gpf1xpCU2E5juK6m2taWFu3tq8P2zpuXLLOxbGUJ8qmEff/dAz3v9z56V88TVmmqqkY5+MbWtp2/eNEqGKTgK4TXxH7eHt5/ZMWKGktW19n3D55IUg9WCTkRA7YSzgOtb1cyYG/ClLpy6Zz19PeJXQYAg/jEEDK9gw9c0YZPn7H/+P0fbW55xZOFkVkAACAASURBVE6dGbaTff325Zdfaa++fuWynhvyQuyjq1evKj9j0EHty/oUc1v5Z0K5PPuKewfY5PvvH0j2yHP3IP8awEBxUMHr8j/2pZrK0R04ZIECEwrBj2+E5/byotrZUQyGtcOaA1xB/cH7V1dTF8CucilaYlhDXa1ekZhE/hBNnJUH1+CLgAeJA6EAJYhJV+KDjhP9fTb27JG9deWizb0csw9uvGlP7nxrr106bZOTs3bl8lkbG39hnZ3dNjkxbb09/WLmNzU1SFYQ36zGxhrJX548d9Zmp1/Ko+L7O/ft7Olhe/xwzN55+w178PCJ9Q4M2OLyshWTFZZqarfb3z+yjUzeOvpP2uTsnHX19FpmBxnJA8kVcnZxP+g5kX95fsBgNAKnPCaqF3RwKDbMycFBW8eovbRE7FL8v/r6+m12dlZ+JNwTmDmSTKV/JHYgssUO3IwAX95DAJdQ2xAXUKYgdxArO/QIkmXOnvV6wOsegCaco2L3CVzjkpPkQNS0UQGB2ogckecAyETgVIH6gu/k5oYlkN0uccafgGFi3u279BMpevDfk18R6hKhXyYZWckjei8wyuZSW5IrcK5KujiJXK3X2YBS1UeTj8UryXlqTXLxufl5fxYhPkYzc7FhQ1+O/cJaVg6cwifFa2GuW2xR1qF6heVSY6A2AaTK4Fv3mM8DJUo9HI9x6sHKO8QHHnqdXeQZg38nsvaK44C+Sn80037V3v7xv/5W7kA3qP9N/CNAPzn678SJEwp2TIs5/AlYFKAy1jaTDIOo6EwqZdZ3oI1OgcCEUAWspHs42EHNmhpOQqIHHW1elw0X/46igw2eTu86ta6pWXIbldJJdySYJrw0MkkmhLRx/TY2qALkPhR6Nrz3tsRcAFUWgq3LHrhJN4kI7wedU1qtwQ+Czc97gU5yMy6njkKzpkECXZgEmNclaMs/Q3I3JrRubCgR2CgwkRShidLS0qQmO8Z/JPRc73ETSr4AzpKIXy4dgqSGSz1AL2OiLKmkaN5KwSmzW5dRcQM0R/QSkLmnx8he1QHB+yMkDxH16cMZUPneSI0JpNDLDiR+NcYIhbAPQBwxEQsGDhJkrUDLgNiVlFRAkGtIEEw0SdDcdM2bFpqKM8RAvkRIMOSYSoVYku4wjY2CM1s4CJxKGjQN0bJF2kva265NyjpmcMD10FClkYQ+vibWILFzeR1wFPocVJqyM0BDMkpNJNfEZd1QvEhje/9AMiA8NxBLoB44kDlMWCsk4xzKMu8DzS4qbJWjtcLn5D7REAZdKvNlNWV9CEBRL9Nj0WGj1j7DOF/H7iPhjVyekeSthKB2gzmX5SkI2Yb0BAkN6GJQYaw9yfugb83QJUjd8F2Gv9LUd7SGsxYoXPDXCMiYgDBwKqPTcKNEFL8ng+3gmyHmRDBi1x6XMR8IYqcsspe515EWGQdpsRHPgewoJ0/KPWlxszukV/g5YgjyAs7W8mGOJwcZNpENDfRYc1ODqL40qGB8gcgGadvW0WUt7e129/4DIZ/2949UPIJCaWhuVGJMy7y5od72MlnpsIPcTIOkpGigsYbfR0D+xsFRlOAhOXOEiqPx9fkkV+bG2iRYbW2t1tzYpOaRvHvKy4XW5HOvy5zUGzTordMUY53RwKSAnZmZsZXlZWtrb7e2llY1ahgEoKELspSfh0oLyoNEFQQHhUx5WYXiOsUt9OPq2hrJyTD0AOnOs8F/AaO1uOkZPkDBjVRqmo5V1W6QTLzIYMhZ5s1qvoiPknqJTKFEqYYXfDkFHKQ3LAiemaPa2GO8N82UpaVFN1PGTFfJM94trpsrqaQwfOTMaW5u8tfLuXa7GkoBNReZFjR+QKtwX1mvQu/QJJfuqSPShcISLbdO7yfJAa1p9xrid0mmXTfZG5wkqhGZTozmGUbEtOSpZFjspsgaRhaLarrRdOR/IGp4bhRkDFMiYjo2DKO8E+ePCvGAvnaNZopw17WP18izcJSN68Zy//357KpRrIYDeyYYjguZpuGB6zWzHjHZ5DXYZ9KBr6zSGaLhiaxkfdjqhniOThQLInjQcN7tH7huuySJhMoKsmIheV9cXrJ0Oiu2WaraPUO4HxFFzn0ADS1TxUxaDAv2+NDQSVHHkXjKZDM6Y/r6e6QDnN8rmB0BrqizJ48fWVd3q11986Id5Heso7lJQw+xGIjTNSnbwNTWSmxmec1KyiutYKV2lPDBsoxWdf54w5bCZWt9Q8MXZECQa0C6kPMLGTfuHfGeIoPhEwUYMYi1pP0vf5ZSPeuO9k47e+aszc7NqSHA3j9mq8H2Ozpy5lvRKeEUljwP+c2o48jf10s2RXr6x9KA3jDVeVo8svqGOsU+GhC+ph3Bjz45rAXiCqwN9tKf/vhH/R4/Mz4+JlZMRSXnk5tVc17yOx1dHZYA5QbdvHCgPGd5edVZuLDK8FlBCiawgOJeoLnP/uLMy+WzWm80IMi9aFh6oeymp+wjBnf8vVhSZtbT02XTM1PW39evYnp1bdOejYzb9evv2WtXXrexsTGZaQ+fHrJ8PuvN/HA20tSJkqGSRBIb4UBrlL1AIwxpjcw2UnmbdvOD9yVzNDY6Ii8E9vzE5KR1dvfIX4UmLyyAtbUNy+/DYmmU9wdxwI1YYc+gfZ7S+ZvezlhLa5OMP/lZ9iuygJwNNPckKRQ8ABzttxM82pCRcfYYP8swFSkuinzyafd1cpCO8qyqCme/VYG6dNQ3PkZRJtEH/zCbaNa5fwrnMeuT64rSJ9wr/sefPdc+EptjY33V/v6jG3b2FPcYNkPKbn35tb2YmLKjBEAYH6zYEehfzuVK+9Uv3rGaKkfPkl/UNrbYwsKKPXo0Zqm6ZjsouGEuOdrqyrK+s4+IB8geEbcZptNk6WzvUKwG0X3h7DlbWl7UUJxhIM8IaQyQsTwHciE+38SLca19EP8vxl/o8zPMiP4crNehwUE1HVwO70BDO2Ib5xCNCkqdpZV1xcCaau6xS1HyLKQSXkLjIWnpzQ2rqii14RO91t/ZpoY1e0QoYivY4PAJo5nz8N73Vl5WZScHhu3J41GbmV62LP2eskrpx2fkW1RmQ6fP2LORZ8pzhwZPygw1xeAlmVSTjb1NjnD6zCmtT2/KeqOe4d5//c0/WFNDne3tZsSg0YAMRvsaMhUdtpPetepUvaTy/vjHP9nOThZlK6upTtrrV6/ZwtKSTc/O6X6JoWj4BjVJFiN6VAD80esGnzLWPF+wz2l0IYNE4kYTln1NfsP9JR6yphiACgFeWiJGhfO0ncWj7LaYcA8IGjUM04KHVGwwR/Ytf4769xFYJaYgkjkB2EZAVfM6GJQLxCApYfJdz73FvBabiSZQqeWy1H0Ae1hSDO68liEHKBRppLkPo9gHMFkP99Vc4hrevf66zLQ/+cvnWHfb0GCb/fznPxVbjzrw008/s+djL+zEiUG9xvPnE/av//rf7c9/+ovr8x8daX3f/PADu3vnjhqYDCrIVWEXMSB95/pb9u03X9n09KzOsoMCRQJs2SMNKnjesIVODQ3aF599rjyEz3zhwgXtj9Gx58eDSs3jw2fjGbBHXnk+KZrajevv2NjzUeU5nA0MKsinGaQI6QxDQWoGnI1ldv7cactmHby4ub0tOcHxsQlncJXCtngFriNera4ue5MtyFABJuO/ozQmz5jX1hA35Daxrj9mtAeABnFP0r1BioXf5fzmvRlIcjZFNQbVQ7UMPamvN/Qznt95Phsb7eRwMHQYspDDw5bJbq/bO29dsKtXztjG/LRVsQcPzT795FtrbGm0j/7Lh7a7vWm76V2rT6VkYs8A8sLFS9aAZ0R2zz3fcnl7cO+BlVSlrLa13e49eGrpLAbqRaupqnEjaepmZkhCWLtENtJuHW2N1oL0086OrW1uKt+DcVldlVKO1QpLdm7WEvhSlCWtq71D8U5AyINDMbI4A7xxndQzhX344MED5WWwBzh/no08VZMbvymGpJyHyCG9nJpxtYgKPJUcac72Za3FgXoEnnE/43nsLGQ+i9d45KicO3hNqMkeWK2Rea4dKtnbaoEtBTz0R6T7SM5IvQObV1Kz++79KVlxO7LalINo8KfgzGewKr+z2gY7c+qkPbl/z95+/YLNTY3ZB+9gpv2dXb50zl68mLA3r71m33131/qRZ3o5Y4NDw7a5vmXt7a22ve33HEUG2HgDQ0PyCrlw6YyeKZJPTx+P2Buvv263b9+1weFhGxkft2RljbX1nLCv7ty3zcyBtff329TMgvywGPSSs/Ic8MuCvcQzIM8htxZIUPWVe+dFo2gG/Msra/KOIb+MYK6VlWWpAgA2w/OIL3JLH3o5AEus/cD0jQA59g2MTupqalbyPB8Yew8JbxueoZjTAjE6mCp+dznnOEx2GTcNE9Q7Q4LcmVgsmON97bvuWNpSEnRB8lkxXPUNr0uPw3NH1pz6RUkG0QxMX0mnI4kcB5j8PT1Iaj56mfQ8+fzEO2pJPi+SnuQS5NaSIJT0b0GgExRSBBgIcmP8Hiwd8mhiAnUysUhgD/Iwnk0AXysPTiY12OfnABlw0yTXnMu5bOgPBhVqrQV2vvo/gEgYpEqNAtY5dQGyujF2c1iiUOn76UePinCs//jtb+cOtAcZJpIDR7eiFdik4poGEdPEWHjSIHXdbyjrO5oIyoiHoimXU3HEocnfiUaWd5Qo9G7pBQtxSoPWCy1R/2trrbur69jgCkTuzOycAhnIH5rAEVUutLhoUO7V4DRCR4NFuqYSGQVEn86qAZpwSpUbCRclkyKkfKpWn5EiFDQkwYXPKr8LEOlqkvv0kyKYph7NTJIaJtgUFkJuSePXrLa6RoOZKKVCQSzkuOQgXJ7HG6uuVe0JsptJK1Du7Yl2yc+o6QSVNZiEEqho3tHwQvoFuhoBlINLxWWyTAWz6JUcQIEuRmNapj1C0HrThiAnqpl071+ZmpHQ8uXX5gFSmJtggkWCJ0QZeC3Q+eHnhMIPxr3+s9Ew3SdG3hDzIYbMtNX42Xd5AQYF3vfyQiDIgfA+JFU8G+nmx6YGEgqV6LGjUenJq1+TDzWOi/g9DKk61Lh58fKlbWxs6b0EntJ3DmkfEEk+SHqYjgDheihMvfhHixs0bMIaMT3PQI30RE/yLEHOi9ckMRKNOrApYhNSRl/h4OGw09SfQxrDQWkyBupxlJHRQecm4qwNIcnEZPLDKMqOeTLoCX5sFrP+NLhK4qviRlLoxXOvRW0kaZXW+K7e3zWvnR8k+RqqVrGA/JmArNAQSXJG3qyUGWO5I8EZsHhi6qbOkh4KUjVC06pgOND78sX+opjl4I5I8Yhq0mcQ4jUgmQILhGfyQ48HnhOFC4wcZ0J5jBAN/6hg/V3t1tnepmKdpv72Jk2ISjXf+gZOWmdfrz0dGdPgYXZ+0UqS5SpA+UwUuuyfrY0NJRZdHZ1iloFYqmtosDWYYUk3pCMmSDoMamt2T40+BgnSz62p8b2vRgHPORo807irsob6OiX+jx4+UgMQ8zoGDCurK2pEUChQHIDEIkax53l97h0yCqnalBIhYpYQhKCGNRRM6vmDuOjs6rJcdk+DCKdde0ObATDDKSQeoqSRBruB8Rab3ewr7iuNCBqmkg8LpsbEbZqYcUil9RO0NIlNNALLqyp1/9001hvrkpQIbB32ooYEqdRxwUtizfnD56doIS5GxoP0Twsu18bejIbOcfAhdDNnAz4T6LPnnH3ViLF58HXobGvXz8h/gmalEPQJeWxoaHIsO0ah44ZvknyA0RAaYQw6oC87GtkTdC+m3e9GHkiZjNU3NOh5RekprklxVfHwUJ9D0hliD7ieb2SDsSfktyRjXT8fjr1ggpZrZHlEZhbvydkVZRwVv0HVB1kZmjW8htg7Yk4wwCqXfwtGwlG+kYYJ5rH+ukXJJwidKFlDL0x0Bkg9zJs1FL005pxd6HGNdU/jkp+qq3VvDR/sekwH7QsAgM/R2t6hZjQ0e2SyYO9wTxhA76Z3JI+Ab4MlzbY3V2W4TWxKllRadnfftja27esvb9mZcyfs+odX7en92zY40Kuzj7i8Dxq9vNLmV9eFaFta37BiaZkkn9DIo/BBWkOD9wQMynU12DET3N/bU4Fb2D+wqReTtrOxpWYy97Wzs8da2lrs/r17QtDTnBOjUOvImaHsG+5lXW2D8iMGIo7URC6lRogp1h/yaQwdOZRhoFIo0mCgQ+FMokor7DtqkKYX+7y+LmVNDQ02Oz+jcwpd8MGhQXv08IHMH5GF4f4SWxhUomGN/BF7lf396OFDxfy5uVlpa0vxRbHcEQr+HEusWHCU37Wrb9j3d++KGUSjXFJZezkVbDSOGYiy/4nvDBnZ3zTmkTVhv7LXI9OMz9Tb494RrHX2k8y68VVBKg0zWis4C1HsqzKbnJqzlpZOa2hs0sCBAQg/w3BXnlPkHxSaRy7nST7Cwcla5DxlqCPGAush+IrRwHjrzau2vblhoyNj9vc/vWnrG2s2Ne0yRMQXmlT1jU3yviB2wkThnEIqbW5+Tp+fHBJEqzMbSsVKY0BNzHWZUUdiE3c4s4UgDwak3MtjLWrQsfm8PAKiRCd5Mesk5hLkEVFqDkkrzn0Kdhr+5Kv8rufN3pCIgw6ajcQ+PTsxEz0njmxfMTiCVIcQ5Imi/fSjd2U6ijkw59BfP/3cHj56pkHFXt5zuPraSisrKYpV8bOP37bKMqQ1anXmIoX1dPSFTU5hFFtj2b2CdNvnkBlpqPMaIVkmyRsQp+xDvIA0GK1JKc8HvdrahBko5sgV2o/kTUifyHiZnKTCdaAX5ufVjOHsW1xatQZ8Eag7ks460JqsqtTeE8CqukZnLLEJ9inrCgYcjSwYSI0MTzHdJN+E6UdzGAYqTYPyUrFILp49bV1tDba7vaW1B+MTRPXJwX6ra663zNa2Pfj+vl28dMVGR17a4qIzKjL5A9sN3kHcq86ubg0+yW8YZpFHVMEGw2S8UBBbgRuC7Be5AoMMrfWDQ7HIfv73H5kVDrRfYZjBYuBc53tza7ua+DBK5dlQ36jcYGF+QUO3X/zDL8WAvHvne91/EP/z80s6RzmTI2NdDaKQIwopG0FRmLYDkBEDlBa656udnZ22sbqma+jqdH80IcALh7YLoE04L2cCaUQJCEcHpbN+tG9ZiyGH0boPjeTIvo31hwBa1EU0zwCDCbHtGt+cJdqbocOjRnGQDhUaWzJkZlWVZQK5KOaUEMcYyFZqaCI5qhJnF7OXGeCC6K+pKredzR27+dENu3LpvC3Oz9iTh09sdmbBfvvbn9vCwqKkMj/55FN7Oblkp8+cVDP5xYtp+5d/+Wf7w+8/sf39rPZ0e2ur3bx5027dumULS8uWZVABCKusXM/92tUr9u3XX9vMzJwdJZJW0GAH/0TuE8zShHV3dtqJgQH78osvA7v90C5dvqz4wYBXOX5oTnJviNfUWhpOAUDg78Ig6FrwwkGKTB5lHZ2Kyc+ejSjGyZMuGJrjUdLf263GPjkoQxYGkTBxYdhLHsi8NqFWIMYQcxjOE/eJewDU+IqymA6289pDOdAPmBX8vPTjpURALeQ5D+tAoC/OMoZI5CKVVT+Qng1a/Lyf2ILEEGetRg8nsT1LS8VA5JkvLa24N1xNle1ub9tPP7xil88P2urCtFUBwjwoalBxYnDA3r55zbI7W5be2rGG2jqbnJy0hcUlu3j5ijyjGNxRmxO3FqZmLFFVbd1nztv6yrptbGctm6P+dG+CsjCY4LOo1mZAzDXndtWA383vKc4eHngTW76T1HtHRevo7bX6lmZ78WLciodHqgV5hpyzvBa5Fqw+5YqBaUSOwLCMng1xoqW1WfFxCfnuinJJuk5Nz9jIs1GtSYATcVABEIBznTPdAZTOdnamsdfX6v2Es0nMYQCgDISDmbaGgGLMIZscfBvDGcF5xppT/hJqSDfJdilD7itnAK9FT2R5dcWZFwCu8m6ITH1A7s2a7+/pttEnj+y9t6/YzMSo3bh2xR59d8feefuKjYyM2vX33rKvP/9SDJOnTybs7Llh21jdkon59va6GKfUOge5fWvt7LS5xSU7Mdhjd757Zm9du2Avx1/albev28Pv7ljv4KDd+e6u1Ta1WHNnr315+55tZQvW1tNnMwuL8h4BoJMo+rAS/6n2ji6d+0jSuZIFAM+CDw4CwJL4i6fYxsa2pJ8YQpNzULMT38n9kOvt7evTs5nBe5b8R+AHN74n54Ux4X6FCmnHfTQN/niOQX7ZvQ0d4BnZMhEwKMl31mlgGGjUG5gW7C2GSLwX996H7AxCvAbzXMR/XqoBsCnKYMQ6yy6fxcPx1bCS9wAUGnsVis2qRxw8K4WD4F3D8yYe+eDekT+8LnU/cYF9VFVRpWvAw9Dvs6uMKNfdZ3hNDeisESm2BEAHPRb+zmWWc4GF5LEkTIGVb4m5gYxuUBegPqR354MK7xPG3gvPQTliOPPcU9YBu3FQcUxQ4tfEKHH57B8HFX87/fkfP0m4A72lSDvBiED/zyWMOjq7hEKmUaSEIaCb1ZzQhDqlv4Nmy+bTRJzfr6yQ+QzoVU3tA0qdBGB9A3SSN2KcVoXpVoUKBQ4WkpU4cAC15shuP+T8UHJ2BMlIbKJHaiYsEIo0EpZouqXmP5NgmmaHhWPjbzW4CjT3XNtWaNg8h7upoPb8mITVZZAoOPjHzY0tXXd1Cg1l19iNeukKHgS5gI5Xo6KcBoPrXRNAxDw5OPCCKMg7+eDFDXJEOy3QvPKpLI0M+SOI4ZFUg5wA29Tc7LIA0oJ0aitIcQozT+6iOakj5jg0oiYyRTyHEYe5J3EMfbwR7tRuP5AkwROMnEW9VsPcpWvcm8KDaETmxc2kxBOaXZkXdRoSBXNmMbnxN5FXgje/ORSY0QugG6jlEWXqlLdyFaogLflirUnfO6Cjub/SaKQZE4ZBPvFIqGkUafwM3dDo1WcTVItrd6qcxjok2ip8vEGvZj1YwSBLwxqQzn+Q6RGyhfVfhVSQe5fwni5NlVMi5AYRpgZYbFiTAIAY5XUZSnFvhFo+OtIziVQ+N0YPsl7hNHINfm8m+wHmU3eXz3ATdt8P6O3ngkcM6OYjIQGUgBQdvcA9gyUgM6kwaPE97myioHnjhUTQjIwJpuSfuB9quhRkesmOFIoAlBryJsEo1VEYPjSTTjfNkR8wQYSED2vP10RA5Qd5H9dl1CdVQcl+ADmBqSbN58WFeTWCfVhkdvX112xmfNSaUpiqptQ05NqWFpZsbW3HkuWl1tHdLUTL/lHRVtY3bSeDSWq1lZZTaIC2zanQTkFjPji0lqZmoaHkmCJUaqlo9nwuEmkSYvYDz1gydTs7zpoJQ0+unsdFAefrzwskNXdTKTEgWAN8UTTwWYXQPda7RK4M/w1QLCSoTpGWbEdAs8O0iuw0kn4azaxv1gxIc4bLFNpCYaj5CAMoIXQHDeZYWPB8nBLsCFQuwnVhnTXniBlvbEXaMGdHpNuLzYS/Bh5FsHrKvekbKfzcu83NLa0pl65yXw6tPQZUMi7skT68M6MwLqyVCZqz4wpiI5DkEu+4X8QQdEQZEJHAcT0ugZU5Nm1WwopRWdGsubExSICUKWaAhDoeBGIOGu5BHCzyepXVjryNcZIhtdgyiht+HvH8+RzyyAHVExA1+qxB89jlCR2pE3W4OTv53Ayi2XuRAcdr8rziEMIR1t5wiejRV6ibhM7QOLSOww6enVA+okk7a5Dt5JJpLl0ninhdnYZXfD7eH63x6gpo257sw3zh7KD5qTWgQaX/Pc9a7MQq17Znz9NQUimAUR3ocDHdGM44w4j/I4aC+E1v76jQpWlG0fs//vAHrdUb779ve5mMrmdrc8M+/+wL++ijj80S0NzR8d1VDGAIub+HbMShzUxNWmtbyn7yi/dtbmrEerrb1PSAxVHb2GrLG9tWXtNgC6vrtn9klqeBAXoTpPmha+Tu5zBHdbN0iiWeI8OW/G5OLJGXYy8MD57MdtqH22V+/sjoDwlKnU15Ndqh7c/OzGrfg5Cj+UN+RMM95gWOInWJrRiDOe/QvgUVy7UxOae5hCQn+tPra5uWqk5prVJz0QxHopLhDdeNDjxDg7GxcTU6ySeIG729vZZO71h//4AatYAelhaXdFaDpAasgh47awS5Hkk+BUmTMsAou2n76U8+NoaJ7F+aLxHYISBBOAfcC4qcwmOa4k+l09fFfA3MB9YSLDGaCEg7cLaNjo7quRLXQe6CoGe9IA2EwejC4qqVluIJUia5FiEl97MqttlrLinlMjKRWkv9pmE+O02DeIaqIPPCuW9Fe/edtyT9NDszZaeGhsTUmptfFJAGQ2c8Uxgw0QRgXw0NDdn8woIMK4mjNEAdwOEeWuwVhjMg8VjDcTAgKZKA9tbAU9IAyBF4Hp5Jc35U6TnyuhTJYlyQA0nG0GUPvFBOah/CspF/AoW4TI6d1aq8uRSgjevRRzkw9imxhTj0Q7AJ649nxO/x/mJlpbftJzfftaGT/ZaXcXq9vXw5ZePjk5bepaHmA5YEXhysxXzWfvZ379jG8oz19vfqvlTTqJtetCdPJqyius7W1tNiqjBIo7lKPOF9ieMwjgAQkUft7GQkf0T85/w80d+vz09Mwy+G3LS1rV0eHQzuqTGUvyfZI+tCua8h2UrelEzab/7bP9rXX35t09OTWg9ITQmhWFEptK6zdl2CTB4oauaYZTM77qlUXmH7YjG71xbxrL6m2vazaTs9fMJ6OpttdwcD74zYHC1NDZZKwZ7JWX1nu9299ZUNDp+xsbEp297J2mZ6z3bxGADAwRBfTe8Sa25ttqbGZunBb29sCLHr2uEeN6TvnSy1ltZWB6+AbrUjqygvtXNnTtnRft62NtaFoq2srBbzUR5yR0ogXeqH4cVOWmuG5jH77cL585Lmcu+oEl3TzOy8ffb5FxrEReZzBFmxkv0BmgAAIABJREFU0bSPzL2biCkSEEo4SpqGGzGUhvny0rLOWhpwnHUHyIyQI4HKPUKmFJ6KA5nUiOZelPpw0VVE43jc8/XYAIu9oIgO5vflmRFkNMR6QEc9AosEzgqm28EvzRHB5D146iD32aC6j3tXhlRWZtcy6awzsYougcckhDUEW4R9XlWBTFLWLl88a2fPDAtwVl6asBfjo3ZioN/+/f/6d7vyBvI6CzYyMmeXXz+jAd7d75/Zr3/1M/vzn76wQsHzY/xibty4YV98cctWaRZnc/LzEONmaMhev3zJvv7qS5udnTdL4LFUEthNBck/EQd7unrkjfHt198qJ2F/vf76VeUd4y9eOKgIwFa4l9wvRrcBK3Sck3LWvXP9uk1PT8lnkryxvbPTalO1YmYQq6j5VJJIJrfKWpsaNajgPTlj+R9DFWd+MxRxzXh5CpGP0NwWY8mHuTwLziRqBjUMwzoTU5fmdDgriU/sX6G3w+cQazSA9IiTDprwmoU3Iy5GmTBqS87quLa4HoH3Qu0nBHmhIB8nBzwghVMm4+zNtQ37zS+u2/mhXltbnLVKNRET9uc/f231jfX2s19/bPm9jJqrqdoGG3/2zJZXVu2Na9esqrbWttY3lSshMbkwN2/bubxdevMtSyQrbXl9y9a3dq26ulb7Sh6PwaNIihCky9ReOZeM4V4RL0HD8xnKUcXoH9De3t7bFWMJthhnEtKV3IMLF85reDY/N6d4io/B+Pi4pPd6e7slFXn72zuKwR+8/468qZ6NPNd59LOf/UwMrc8++1zDEBQAiJU8U7IH6qJ4prH/+HMcLLBfyQ9iPes1kftRcLYgK0stqJyZtRAkv/jcYoSWe7M2esJxnsqrL3zFOkGDKnLt2lqtJ9gPnIMCkiiHdqncrs52mxofsWuXL9jMi+f24Y1r9s2nt+3mh5c1iHvv4/fs9q0v7eTJk/bg3qhdvHjGFuaXbWCgxxaWZt3fB5aLJayxpcUWV5atvbPN7nw7ateunraRp8/tvQ/et4cPHlj/qdP2/Xd3rav/hCUqasWoyOQLGlrML69qSJ3e2dazbairU25GDiTwVKkDRr2H4iBR7gFxmbOcXA0fLXI82NH0ttjbG2vrkmB7+XJSwxZyCp47zyf2D7gPAseSn+sMrNR39S80dKI+ddApsZU6nzMIplIES0T/RK5PwDTktQLYURLbIb9R/ybIZFM/xMED/80zA3jIfpX0Lv8H+IH9GzxQYw8RwAS5DyxV1giS27rEwLQh1sCoIN5F4JCAD0ECXkMBPlVpQgoxxJ3dtDNX6fVImUX+GIAYGdy6NB15qgDMIQ6Rg0cGf/TmiEMSnokDjMrV75EENsyS4ClL3eWMiox6ebp+gYIA+9J/Cqy9Uu+3CGjLvdXQBdBblH5y9mo8C38cVByHgx//42/lDvSUkPyCqn5l8gy6l6kiG9M3GklcQGayeUEeByNqklOkANg4ceMhgyMpGhC7AZUHMphiQslAYDwQtGjq8TNsWCh8sckmOlfQzSXppRgimaHwYkPHQBuHKByoOtBDQiuEQGjkkWwRjAiekpoiMQJVG+RbKiocMQqigwYxRS+Iz2hqKukZEBApjAOdVkywzmbd9JR7hw4qQSg2jzhQXTIEXT5HqTm7xKUxomyGEjeKB9CAfD4ZKQdN9GA8ThEBJY0CnoANtU/6fyDnqqqFIOO9YlOL6TEHKIgNDitnhnCdBauodpkBDjfuF2hT9wJwFQiCbPzimuLBo4FRkJmKiBYOaDUAhHBxaSEKSIZD8jPRJN4btD7UcM8S0T55VtI6R/uwqGtxc1ZnEWA0RALCwcQ16aAL9z6bzwYmjBvkcQ0R0c/PcR9ILCMdj4OZBjJIHn4OVBmyTF5wOQPFh9k0Glzvn8aPrj0UThQhSD5xHrA+aBRwoGlYkXeDXaEEQP3IeLSoSbl6JmFNcp1R8oKfc3QRGteHSh4dzeDDBPf3cG8GkMZIhbD+OUB9ck4xF5gQMgwPrJBgxK1rL/WGKc1qN0F0lBL3Bp8VhiiR8eBm5k6H96GHS36JoRT8So69PALTh/ckuYn8i1cN6HJPwoOmYqTwiprI84LdE7RfvTFKEyqvQoXGRmTQgCJlz0UvEYofXpNBBfeShgOGc9xf0HJIJazMTFp5SVGMnWSiVGhI1hVJ3PrGlgYUBUtaZ2+/0C+HNExBrKs5X2bNLU1aZ2jsFvIHao4w1NnNZSWPh4wSpq4yAy7gBYCmpcdP0EogMGloxMEON53mJYgfx2cUj4seNa2gTksX003MJJ+3R2Mh0HwlSF9yjDoiJol5FFD+ai5pOOg60RoQBMkd9jtJEl/SkAbpXOKxi+YlrCHurwKqTMYcKRmHyS7F5qgyBnygy1X8lZTotXhtmox8LhqzFDEMDBz5Vm619bVuEitjZwbHPhB3jdIja2nmOZYoKeU6NMirc/kqvqNpz9pnCM6/yawWZoeKIu6x62Vz9oBOYey4kwF5TPMge7wf+WxRgonr7OzolCFzbMrxeblvrD++fAjhg9KYnFNs8f7EMIZALt3iUiPe4ILlFQ3vXTf2h4bYzl5zg9todq5iLOinavBTLAqxzHf2g9CFYfAcUUJcm5+pwdeDfQvLJPheRE+TOMCNvx9jPL/vrAofxvK58agAmcv18G+//sdfW20lhuLpY6Q1QzIxhVK1ilsuz+BFCU1dzFDVUJIp9qHkCkjiuQc0ONlboN6lsUpcp8kAGjK/b3UNjba1lbZiokR7a2ZmVqg9mo3EB5pbDx88tJMnB213d9t20uu2n9+Vznx1Ra1trG1LQ7x4dGA1qRL76Bfv2/LsiNU1VDtrrabR1lc2bGv3wCrrmm1je9cSSPkU8BTKayDDILK6MmX5LPKJbl4nRhkDZzXREJ4qsZXFJVuYmbXG+kZbWV7VzypeAkbAtNd4dshpNcukHPr+0uKyhg6c4ciqQNGXUW5kluqelEsfOlXtUpk0nmkWMOzL5nNC8p85dUYN+nt3HwhR7i0VNyFHbiWZTCiWnh4+pYLvxfiE5fIuAcdaZk/xjFhXsGEZ3snDZn3d1re3raenz8orq2xhcdEKh45gTYH+4lwQarZgTfX18qaZnZ3WGV1TixwfPgjlKrjq6xoMLXX3rSrK4wZJN0AgeOQQ6zraOyQls7mxEUydy/SekmkhpmhQWxSjbHZuNkg+oKleYotLK1ZWXqMhp5C0paD0iJfe2FABqiEF51dgsPrkIujd+9nJM4ORR+OCJviV1y4q5k9PvZTsCvI7sDDxwiBToYFLDsHQmrWMHE5bZ7s8fhwd6LrZnPsMDsSmQV6uygdZMX+SdBPMrcCkdB8NB+QQs1wSwQ3KiaHSb+bMD/rN/DyfheKYc4aYld1ziU+haAXAQI6D88l1oTkrDw6dQUFuJmnM4EsREXrkKs7Y8jpAg1ENnnP2wY237PTwSd1fmv8wCcdfTMpfgN+j0bWX2bbO9lbLptft8sUh21iZtTPnznjdUEzYdnrPnjx9YaVlNVY4AsSEpI/79NQ11DubCV+6nAM91IgJiGu1UBNFNYW59v+Xvfd+jjM78/2ebnQ3GmjkSAAEATCBmUMO8wxnJI00o1lppZXulnevb5XL/su8W3XtKv/gdXmvXddeSRNIDicwZxJMAAEQOYeOaLg+3+cccLbK/8BVDVQUOSTQ/fb7nvOcJ3wDZ1lhA0m8hC0uL8njRoPioHNPLORsRWqN+Hb71m2dYz19vVr3DP3cHy6ps5if5UwiDpIb6/PkkcqrFytTpujVLZnQ1uUaZHQrZuB21fJrq2J8XTj3nvX3tdsSHhq5BpufnrH6bK0dGt6n79tKbNvDBw9taN9BW17ZsNX1gs0trtjo+ITY2fi0rW6UrL+/x06dcuT7q5cvbA1WEsPPwNhERoJzliY+eylbD9iLBotZNl1j7508Jt+MteVlez7yXICZRJLcHwk4wYJkbsxgl4Ydutt7dveLFQQ7qK+nzybGJ8Q+oQmahoU2NSUJnzhEd+CTszi8aexZNMNIYj3Xy6CGISc56q6ubhsbHVUeBqMiv7FhRczQQTnzSkJZI/2kDH2HVSsQCxMBNY+9cebNGGdlaoYROzQBaKQmqBpQwdw5zR50oIWfnV576SwGpMUcODRaHaRDXZi1Q8PDanCWS1ti1szOztvrN6P+uZEOhnlQqVqpXJCZdltzo5VLeTt+9JBtlQu2MDtjlz+8YL39vWIl/eXf/iSZnqkpBhUzdvGDY3bk6HGbmpox6s+vvvrWKuW85OOIwxcvnbOrV6/b0uqa/GA0qEil7fDhQ/beieN27dpVNf8xtZd8oZgELjeG4kD/7n7bhcTpDzf03NgzZ8+ek4ckAyyt/1RgsAcENNJPMRck32PN0/j76PJle/rksQaB7LHBvUNq8sJ+dKAO50+dGH3M1TEoVg5fqdjs4rIlUimbnsKfyuMyptRCJ4cvanuuJ8rf0rQjZnnM+xF4CkCImI8MpZHojY06l1mNDG3/GWe4844RCMT7k6/LkF35m/88sZb39jPDdfgj6ER5G2dRd6ck9dRE367Y2uKC/f5vLtuBgW6bnhi1HEzsRMa+/fa25Rob7eJH7wtMAZujqa3DHt66JdnAix9+aOm6Oluam1eMBgz16sUrW95Yt3OXP5IU3J17T+z+4+e+B2Hpyx8RX02/H2KySoXAvR+Io4AtiVOJrao1NzTascNHpTzww61bGrQdOX5Y+RKADz7b3/7tb+358xf25CmG6Bn75Bef2O3bt23i7YwNDey24eFhu3rlmlD0lz+8pPr01u1bAgx8+ulnqtP+8sVXkoHSALdY1vvF2iI+iwjSUX0R8t/IBPahkPcBxO5oaZZUVmTOwEAmf/Q611RTRllCoeEFCIUB7w11/o06iH4J9T1Nf1jwDDiWlxbkn1efzSg2eA2Ttd293Tb2csSOHthnsxPj9rMPT9sPX31vH1w6bo8fPbGPf3nZvvn6iu4HMk4nThxXDjAwtMeeP3ui86NUqAjEgnn59Nys7e7vtTt3HtmJY8N2784j+9nPLtu33/1gBw4fsbv37tvA/gNWSdbZd7fu23p5y1o7e+3tLAOFPuXI3JW60ITv7enTeifOSHYzSLlqaBE8CXhGrGfYbwcOHpS8L0N/ahak1Pv6euz161EbGhwSOGVuDmmojA+9zZTTs99KlZKYIWKHSva8JuQPDtZVr02Aj3d9AWKohlDplHI3cgh5FNLzkfy7514uuY3sq/fAeG9yKKQU6ffw9+STqtXSaQGneE9ycwHJWD9B9pLcJ6qToNrCUNmlAn1N+BmxLYklchXJwSWpZzbk3RNZ8wywxZZFXhWgcjYr4Ah1CzkQ+bEMvrerWu8Chsh0mzzP5cHleyUFAxQHPG44Q9QZRfyZ8x0ghOpY1RQuIQJIkHvFzwIKcMCc1x76nuBXwRqnx+T3gXPWAd7eVvK9o0rADVF/YlTsnCw//eGv5g4MZettZXXFEy+ZWdZpYDAFLbu5eUeHn2BEU5zDiGTLJ8nbajBJ/kimj45klfxO0PT2KWHCpianrXtXl0tmqPnlOvgkHBwy0UyJw9tHi57UyOyUxhqoRVFzXf+b5MIbQxRnFBFrwRjZzc4IIhFxQTBhSEGA42doRtKopWiZmZlVAsBh6wa5HpDR9SfRFhqFhmzRkVy8/+TklJKF+hz0Om+ucm/ioEADjkxKRocMEAiWBGHehwZFRP6BNuU1XRLF30uNvZjERW+AZNK6Ojt17chOYUDIQAeKM009PqekBUJiRtMOfXs092ITDapnoVxSssw1wJgRSjvIxezQCIO/QKRm+mHhEjDcc4Kjo3sZqHhi5434QLHWYeLNUH7XswAxiGxB3vUx+SIQO82YgwV0D+hrN3xmIEPDjhpFJkhiKdQIiUnRsboBnb1GDBbQdEzJ5xcXhHzdM7BHz5kDWbIKCTfGpYHJM8TQjedBkQbbxAcJjqyMUicyScTzAsRXaPBSlNWm03oPElAltdK7T2stkzSTbFNCUQTy3zBdaFyAxHKkUI2kBRg48CxICDj0ZI6OTEXQ4nXJJF//aihLZst9UURlr3HZpPh3UUs+Io8keSZ2hDczo8QBCUGkWkbJNApuin81sZGeEQPIE0P5CETTvaD/6Il8kAYTJdsZHKJJg0IL0lM0RmmcRLQ81ybd7HDfSQpoQsdGNjEEirjMvLK1Qn1gSsbeQHOaayFZRrec5wASikRWbJpQYOzq7rD80oJlk8jVZCwBKgGkS0uzhgyz80u2XihZsbJt6fqcrW7kbWll1WpzOathSFLCIJnCoGrdHR0adLC/8XSA/ZJMe9MQJBbNFJr0zsJy9C5sqLmFeSXGkQlGY4F1jSEuzU556ySc2ooWP7FCBqsBcSI2EqifsH9ijFQsC8mREJiloqMcA9NJA7R0xuob6kPRRqKUsnKxYo05mstOxccnoKEJP4xaXScDZOI+yGvQRyAfeWYUDfzOgJbfifMgwdlLFKnsMZJ01/10hgkFAJKA0cgQ2T7XuvYBIEmpUq0EjU3/7Fzz7v7dNjszK0o3hTsoJ9cdrdF6kDZw8DsR+jGw6qK3jidunsiBGpPRdaApx4acpAjzeTtx/ISumdcGpUwyyVmVq0cHtuxSXjSKc7BjQDdty4iZv6R5xTpAxg40Nes5k6pVY0ADDKE2oUV7ESRWTTFIAUmfGUk/l/TgczhbAWS46ZxlH3e2dQi95o3fDcXNSLmW3BBNrbA/KejZczIgNlOTTWj0QkF7hcEZZpbuKYUguumchmkHUo+GKIU7ptBPnz3TZ+eZ/vEPv7Pl5Vl7/eqFGodIsuzdO6TiD8Qb1wzLxLWvt9Rs5BrZY8hFCIlVKtrbiQk1MXj2rJnVtRWtjT2DA5bDHyRh8qKiynj05Km9fTtj9Q2NNjo6Ln1lpAzY44NDQyqqWWdIuDGkyGQc4ZXcMsuvFay9rcOaGutsM79kZ88fs6WVGWttb7REKmkrawXbsrRVa7K2Xqza/NKq5Utb1tLepuLPCyfMZrOW2KY56+wY3o99SrxhSFHCKyuVth++/c76e3fbGBT6qlPWkU5BnoZ1gIFmfbbePvnkF/bt9etWL2PpDSGZJ6emRdNnaCADZkmrwcBiwI8pYdIWlxYEzOCe7xka1ECZ4Q3XR56BgTgDcvaS5xAZ+/Of/2QFCsFK2fbt3SckGENDnhlIRTdEN4ExNDxCPz7jvhCZhpztP3TI9gwMSvaJpiTyAKOvXtvK4pKkK7ZpnleROCjYR5c/sJmZKQ2sALXwWcij2Fes2Wha3NraLuNW9h1nG+cMBdZnn36mPBHJCdYjuQzXApNmcnJSGsIaprS1amirRnKhaI1Nrba56ehRmq8ATiRbhEcHOYSQs87ict6RI9Qiss9BGBR2Xsjqv5CptKrtGxqwSqloM9NTkvpg3WJw3NW9S34cGWkRp9Sgr6t39Cd5MjkGMjnkKCzI2kydG3ouLTrbuJ41ydrCZNI9NPg+8hiekYwmYcipgbeuPKcRCQyKcRnceq4Uaf7xXOG5s+d4LWIFxS4IcO4jklvR+4V96MxQWBaeRyXERHFGk0tWlfW7x2YGjCUV0TTv0N8fGOizc6dPWxNsYnlYZOzR46c2O7cos9KF+TlraW6wpfkZ6+5osT19bZapwbC6Q8h2mvsjL9/Ys5Exa2zutDfj09bR1aPnmK3PCgEq+ZfmZjHumppalNciQ0SzdTO/IdBJd2eHJGIABHFmkYdwb1XwiwlHHgYT7R37oK3Fc32aVDQDBHbR/QD04GcCZzhrOJHY1npGs12sNFjS6Rr5mOB1BnhrIw+qHgZdVWu5tSknb44TR4atu6vJGnN19ub1mNVn0pIK7e5ss1xri+VXV+3m7TvW0bXLUrX1VpPOWiqdtVejo3b73gPlo3v3Ddnho0f0rNnHX33xpYYdnR2t9uvPPpMUiPJuNSvqXJZV4AKTlwhyRQwpmhrq5O2Bh0AyXWv1uUZ1NiWJBLM5lbal5RUNQ2lq7d+7X/uRs4BG4alTpxXXn714Ib8VBnYz89RJrulNnqshNQPMGs4AAEiwglLaQ/KlEgoctm1CPl/EIs70lqZmZ1QhP1rIW1EgEZqVLkMLG8hzT4YNeEIwOHOp3ugdIG82bSNfrxHYxfnKWmaorvwzgI7YH3yPPKZCvRNZoORdyuRrkD6mgbRlXZ3tysfYB62tLouIBBzMHnIY4g4M96aGJp1zMFkqpYKYdh9eOmub6ys29gpvlG07d/a4nb/8gZU3YAGu25dffm2jowt2/OQ+O3HyPWtt79R5fe3ra1IwWJxfsj17huyDDy/YX7742pbXNpWnIu3DQO7Y0SN24vgRu3rlqo2NTlgVv6LtpG3RuU7wXJCtrciImJrx9s1bOrPYH+fPX5C04MvXrwIww/3UVINo8BbqbiexKB4AJDt/7rw9eHBf939pdckOHRpWnsX6ko67BrTOfsUMuKOt1Vpbm9QPYIAyNj6p/I5nxbp16cyi8gSYg/KOwP9GjTvq/LT2vgBOqoXDhCrk+bwOMYhcgudBPcWZw310iUW05Iu2vuaNbiZp0ogPPoasJRDnS0uLWpOSXoRZFAahUQLZZW4BynGd9XovhnBdeFQsL9gH547a6RPDtjAzKcbC+mrBfvjurjTvL/38rK0szavx297cbt98870tLC3bZ7//ja6JQSZxPllN2ItnI7awumqXfv6Jbdc32M0fbtt3mHJnslYkF4kMBMZ41A/4kci8Gy9EZ6xzrfRwCpsl6+nqsPdOvKfz6V//y3/RIOPkyRPKM65cvaa496tf/UoAx0ePH6sm/OhnH9t339+QxNzAQL8NDg7Z3Tt3BJg7OHxQ2+3ttOe8IP/pMXz//Q1Jk0VPvlyDo/jVD/BD1s+wMGhxRm0Af2jo5D4H5KYM5dUXiNI+cMSCygI5M8+Oc52+CrFcZs1B+jaCwjhfIxNW+QRN8yJMr3ofogm8ylr3QSuMuq6ONnvzasSOHdxrq/Nzdua9Q/b6yWPJtz1+9Mguffyhffmnv9ixY4fs3p2ndvr94/Z24q0NHNhrI48eSI53aWHTctm0Nbd32uTbKdt7oN8ePXpiJ44ds2dPntmZDz60K3/+wg4MD9vNW/esd2jQ0g0tduP2Q/kU5do6bXp+yXp6d9vi/JxiPrXh1Nu38pUgz8JEnN4ZATzmL7EW5/ORUzJQPnHypIZPu7p2qQ5iXQMQwXtwcHCvcjQfVDiAwtmTPtin7o8yUNQt1Gacr95fAojl0trsSUkqCZzl4Epng6e8pxKMtonzcT1IGimAReQjQn3S1a18S/VyGZlD5GMdMLeytCLZJ9a5Mz9cEYLamzguUIgk6hwA6/1GZz5wZnOdvB55gxtmO/AYZjM1dWTccL5QY/ElkHI6bbOzs7a6sqaeCIMQMSGCJDZ5guS/BRJ2Y3CXMHfPXbFeuZeSoE8GVrz3obgmelVz83P6zAC3qW8BKO1IxAcmkfqXwTOU50u97z05B+kB+NuZ0QfJbu0DYmRq17l3ETOknD/99tMd+G/5DvQkvekniY6AnKbZgZF2bIDz+QhYu3b1KIigZxylf0iGQO7TMKbYoLHgWoqONhVjIF2jJIxNTkIcD69I2YuN1tjEJhBGCp/08qSH7QdgLNhisFYCSmBbW9PBGGWLIjWO9xJSlMSGxjD0r/p6NRVItiiESeBJ5KVfB7VuG9Rzg4wzfeiCrwOoUJpNbo76Y+NrDgM3wgyYacysJQcE8o3Ds1GfQZqdwaDIP0dVBav0zJuarVxxlG5Mvgn6ap4FA1a+j8JKDI0tzHw2HFWgQArdLqPilftJ05FGnGhomAAyIJHkAfIBbsIk5BzU2YB4VnAUY8U9NYplJu4ub+IoCJrPTI2Df0XQ8IskDDW4g2yUfwYfArxjFPgkWWsimNHxHClESTD4R5I87h0NOSGlm5qULNE8Ioml4QqynmeiAUZo4CKjw3CD585adGOjslCNcwsLav6pI0hBJCSVG70qN/fHtpMQ16SCV8O2o3H02XcSd9AY3ngVaiSYtsnDIeGeDSmQmtIcrNE1uBarSbrIB29Vy5dAfThlNeqa674EE3A1+APDJDKFYiM0DpFYi44kcURhXDdasxxeO7RpZ7bIGyXQML15zDql0CxLD1IJRJDsSoUEU88uXJf+HBBO3ix32q0knUCQhiGi9khANYheHuRvRBMNLBUklWBWYBiH1JIOcgwj11aVHIBMEfIhyGypqbe1ZS3owAcmgpIpEKWbBWtsqPfG4uK8tdTT0Ku1RrTRFZfqVGhgJElBl8rWS/oFE8vVjU0h+tY21rVWhFqo4jdTbylLSkYFBBpYNf69LJkF18EUFRy0Q4hzmXRWqFtnkvgaowirq88oyXMzPAp4EDMu4STWmAZoDUpEWROsIQofmZmLSusGq6wvafonMUV3413JECDpZUk3lStuWnHLKe/o2Se2EpZGQxYvoq2ybZQ2LSnfHafmkpBJOgzhBXkIObuAz8cvzgZYbGiBaj0mHHlCHIpJq9htUGODkZg0rMOwlZgUBxUYhgoFFF6H9UQcIj75eidebmjg4wkwSDfQd2HwSYKpZlRFxt8aVG+5UXVra5viE79gnBFnKLJB4VBcCmlZrcqUmfiiwSlSDqLcJq0+i78QgzO8gEDuMiBZ1r7YyOfFXmvv7lHTLVGTsfGJSZexQtoABBdrWOwoZ7EwtGGA4V44PtAUwi80SSWBo31jVhKTKWGJyrb17+pR0xdU+gr0XlByNIVA87FHRDOnEHRkHY1A9hgxRoNcmEzIX9CQyaRF1QYpxXCH56R4IeO7IHtX3RJFevzNGz0b7uMf/vB7y2ST0uynYcUZybX2D+6V5APnjaQ1KErUNHKUlYrM4Ffz4O4d+/67byVvRjOYe8FnRwbk3OUPJU8y83ZKHgkULDU1GXs28tyGDx+xly9HVUhpUCOaArquAAAgAElEQVR6OE2GnBpy6xuwMiiYaGZVrG9Xt1U5F2oSVptO2YsXj+1v//73NjM9aZn6lHTraUVvFiuWyNTZ7PyqmieVIIPCemJtSPINje6ky/BIIghWBUUtw1Wa35Kt27YH9x9arr5RRX0+jzwBjQNnKnBmM6jIZWF47fcBHNI9NE+RxqTZtbKmWOetdEf3eeyGUs9wFy8Ps6PHjtjx48ctX3AmEo0F9hUNfu0hocaa7YMPP7SRp0/tm+vfuBTHNhJI265Z3Nsnhsfy8qozGhmISmqD4r/eTp0+YYP791mmvk7XtonGrmDHpnu/vLgkbX1iNYPblaVlG943ZK2tSGEUbGjvkNY8jTBkrpC32Ltvn9YSUl7ETrH9DClKzyvVFDZvErtcka9NzDvn5+eEZOYz7NnTb2Nvxj3nQisYKQxYWTQ4oedLvtJzFeUtknF0pmFE5Oq1kwxmXEfYm1kuAYEUBFpNrKPTJ09YfmPNRl+9srNnztjk1Fsx8Do6uxT70IinKYfUAHG6G3N3FflI03muTAMlyjASl/kcAUQc7rsDPCIjklglk9goBSW2r0vK0STgfBUDAhmCIFHJ+qKJR5OZc0ON6hC3HTDhjAqukT0jUE/InzmbmhsbLYkUDg2bSll7H3NphmmrS2uhYEeWlXsOsm/bdvf1Wmdbmwy1UwyZ0xm7efOOvXw1qr0LCvTcmdN284frksC5dPakjb8escPHj6o5kc012tjYW3sy8tqamrtsfRN2bkY+BaAsiSCSUWpulpwNDSQYWjQEGKpyJjF8YHDHOiGWCYyyuuL7FVnJkjMr3fPNwU9IihDnOPdd7tL3DTGNgSwxeU6D15TOoaZm/NwYWJeUa3J/keBggLG5viHgycz8ghUKzoqhydBYVyuGwEcfnreu9gatoebGnE2Nj0uOaXj4oGJfqj5nV7/82gaG9tvL12+kQU+sa23vsGfPn9mL168kB3Xhg/NWl82pyb2yjEb8qrW1NtjPfn7ZFmZmbH11TbGAoRSfmUDB8JFcCBYpsREvkX37hmx5acWqybStrHljhXMFVDXxXOzyDAjkjGoHcjRyLHIOBtMaqFe2bBVZinJVWu/USTS0hXCWprnLkNA8FUOadcvZSu0jzzD3ctvd22sT45N6pl0dHVYslAT4KG1v2SaxSFJNSeVHykMSrE8YjrXae6oFMRsNYCKxt4PWuORsQwFO2GLtKw/hmgKK2+tMb5pSkzpK2xUCHPAGuwSkfkbNfZ1VynuRm4Xh6g1wgADEcAFN8nn3BmS9AVSQmXnKzpw6aVuVoj15/CCYnJftf/yf/gcbez2qhuEXf/6zjTyftQsXDnlNVk3Y57/9zCqlLZuenbdH9x9aIpGyU6dO2Hff37Sp2WXbyCOxumXZ+owdOrTXDg3vtStfX7eJiXmrWtq2QRSH89DZtNvW19snn4pr33wjxQPqkEuXPpCs5ouXLwUSigNSaro4BIqNYnINH1aYnTt7zp6PjGgPlqtleY6Qd4+/mXDEsZg1nlMw1GfwD6NGGu54B25tiR2pHJizN6Ce3RfCz1/itc6b5eUdz0HVrmjYF93jL36xf8V61+fy4Vv0bxDgLDzfoAHoctBJbxT6sMple9WcVKPTgT863wPv2fsGCZ1tSHFRFEzPwn7JWBb/yrWC/eLSYTs0PGjjk6+td3DQ8isFu/KnH2z/vkE7/eGwLS3M2VZx2zradtmf/+0LW1pZs7/53adW19Joa8vINzZaYWXdnj0asZXCpl36xS8sVddgN364Zd98d1d7THlK8OHUMDAoLnD2ScY1FSRlAfUFYB45N+h5JHzu3bunM29wcECDpLE3Y4qF+II6k8xzYAbqrP/opUTPAfk5QARItnEvhvbuFYAMFiUN2sdPn8pniBpIK2g7YesbBeVLYqiLocTQ1Y2PBWYD6EOsDj515DzsRfIFzjrVXyHXCrMOvYbUHVRHbwU/1IyApvjwaFjGsC14g/G7vOKIBZL2cwQ690+AnaBUgc9Ua3Ojzc9M2P49u211YdbOnTpsIw8e2JlTRyUv+957J+3KlWt25PCwXb/6yC5/dMxePn9lBw4ftLFXr5TLbKwC2mqSjOjS6qo1NGdtZGTCzpw5Yq+evdCg4vb17+3A8CH74qvrNnBgyMrJlN24+9SS2XrLtXRYsWyWqs3aPMojDTyLtE3PTNvg4B4NEKIsteqakMfrvBcoMaHYjYfI4cNHnIUqOaeaHWAreRjST+Sj5Hkuee2ND3ov+H3uDJYCMt+lzb1mjYoV8swMXrGSLEXGPUgRy9sVyUDlPimvEYkLAo+4xDm9QM4EYg/PW16n4fyJTEg+L2crtXOsDfmdPpAUURhShBggVlRg5TgixYdknG2AJll7fA8/B+gINr36VJJUJz/zgRjXxpqGcf/s2ci/yyP5dvp7XA97S9LGeMNi4N7SrN4mw554vnDf2Iu8j1h8EchYV6deH/Uoe5qBPtfnTHOvE6WmIUatDzzYj/wd57HWQOirkaP4IC949YZBjf7up0HFf8st+Z+u/f/vDvTWgEpYUxOEUQWJA2ZeaPEydICORpBfWFyUGSMHxcTERKDQbktjmEQIZBxIBlDGEfmtwygY8TDJZZOT4KkRoGa+S0hpQ4ZmexwsSAue5ksRGpkPC9RAU1N2awedxs9KEqfqJqsgpoT4Rh4q0OrV/Feh68FEzIVyScUZxlEqhDFNDqhWDrZkTUINB4IJd0aUdJDPyIpAqVv3CT1FE8GBojD6DZBUc/0ghNVMl5wOTT5H/Ci0BkkPrikmYgTc2GSODeJYzHJASA8aA7hgZqe0PuiOO7La75MKVZprFMBBgkM6niC7QZWgoVyX9YMqmFXpyArUs6hBny/mlbSrIKL5FWQFAoHC9ZBT3mSOuolcQ2xSy2xOCYnfI02AQ74pNADIrICK4plg2oW3ACZeBGIOOoZgHFDcfxJwrt+RX+sqxvmMTMlpgrC2KNrwEZEOLcOEdMqWVle0nt2Y2qW15FXxo+R3R9xQi+VdIaRxUkBhxc/Cc5Z+JswGEm0o8qHZAING6EQSK+mVQ8vE8CmhAowCmZ9BQogDj2vhuXLYuwGcG4CqeSVzcZgWzljhsPJrd/1CEkQ39KUAi1qS4RYzZMGIKvxb3FdqjNSkXCu85EarOkjD7YhJvqSFwrDCPVS8KI3NABV50h/1BlAceEQkjTe5o4GaN2RINrgvNAAa6ur1i4FIR1uHo+CD7jbNsjXRLqGgltSQ8HvjA0DJ58jYyht83HvFCdAeoMTTGOhVrKWpwWpTUFD9OmjAZXM5m5lftNaOLnuD9BNoHgyLgz6kPBlI+Kl+gvnc1NS0kNkJnidNX90/bzxTbFH00Qzk80GFdn1J1gbfQ5MbZkHaSmJegcytsVxtnZLIKKm3axda2+sut1epaD3LUDnvBmCRFePxoKymjn9mUIxl6YUKeZ/Eh8YjHrpWqe2UBi9cJ4PKak3V0rlaKxeKLt0geYOKBh/5TUfY8PqsdUeg+fAUrXWS4XeapD404Iu1yHUIyU8yFxhBPJvoZ+R0XZ5FLE59XWvft3eowYb8Fah74iVFq5hpKTfh9oTUtWWRyaHIIPGUFF7QZKXRTAzX9/P4wrnCGouUYK557/69aniT+NG8olmAlExdFrQ6JqklyxdWtWa3tst26PBBa+vstPbuXnv9ZsJKW9tqwnLv8usbNvnmjS3PL8iMk3vJdcSviDaSXjPeEMF7I8ZbnQWJqq+5ypa1N7VKSkweIvivZFKSKAKhSvzIqEPvni0J9kKYsnL9jB6q5bISaBUzDErMLNeYU2OS9aRzIjR3d/f12crSku3p321Pnz2V8AMeSJ//zefGo+U85eeJqexvCgk+Gwi9WHzwOWmisN5c7qcqObZ7d27bo0ePpDFPHsF1E68pFM6fR6eZAUbVZqamtX+Wl1ZFjwdVjckodGmGaCBZ3Yy9VutMg+A0XilJ6+nukF53TaVszx4/lMTG7dt37G9+95ltVgpYShqdVdlLpmptdbNohYpZGdakNomf67w25wyDNAZSyjO4RzrIgkFlMKxlbc7NztvSwpL2G+bOrGGeI2AD1mQuWy/5ly7Mgd++FV0+iVxFMAQln1phQChddC82iGkwkLa2SvJeyNTW2IED++zt5KzyHVBU7v2CLxWFng9+aNgjWcP1v3z1akeahPyEPU2TkXNTTXMVtEjmMDRosr7dvfbrz39tS2vLkmIhD6Qx6IAOl3IkV/jz//snDV5WFlesvaXNNtaX7fixQ/bi+Yj0qpF3wluA4Z0boNMgD/JEtbVqMEv6rVIWWh2jciQZkK+iWXfo8FGdoTTMYXr6syY/YC8hU4MZZ1k5lyPu8BOrt42NdW9ABtN45VjhS4jvcI5GCj73mNei+YVMBk3/yhYm6UW7eO6crS4v2vTUWxsc2KP1PTY2Ye1dnVrfnOF8gc7n/tO8ouikeU1zTUyngCbkfaM3jArO0JijoS6EonItv1aGccTImBi5xJqzrTSICGtfqNmQR0jvOJz97tnlUpTyFfLkyweVQQta52JornIvkHwhnmNEzhnLdQtQXXFpSBnByzuMP5uGFDRhjxw6ZHsH8aoo2OomppEObpqDtdWUs+XFOdtYXbK25jrr6+kUAKWxpVmx8unIa3vy9I01trTZ9MyCdXb3iFUKMMJlpmqsra1dTRRMLefmFnS+yuOkUNBAA6aL2DdiB2K43qL7R+6Nh4hQtNmskNLcQwYUe/b0Kp9k7S8urbzrZSDD2eDm9aw11gV7gvWL7Cf7i58hltF4ZjAOoy5dW2fzizCn3OsnV5e20uamnX7vmPV2tdnK8rxlUgy+aw2+bkNDvUBSDCqufHXV9gzutdGJSemc1+UahbIlPi+vLtvNOw+ss7PdDh06omb+yLNnVt0q2dEjB214eK/8H5DumZiYVP6aqkHisGD1dTA4ixqscs+zmM2KCZ2xZLrORp6/ssYm0JsFa++AIbAggBRNeAFngr8SZ3BTQ6NYVqwH1tX45KS1d3SJ+UEcInaS17oPDXGYteOyo5ynGfIeuWhX1cTnAOnq6FSDbGN9U+c2MSvPc7eqLW9sWjYHeAffIs8ptlW+wXPaVs7mUk3sL8/3BC4IUk8aSkLNCw2qmEMLbBVyGZdPg7XsYJ4ff/E9NBtzDe4rRj3KsAoPAjH9a2t1j0DZEsP6du9Ws5qzgli8uryiAXmCYXylJFmmtbUle/XiucAy6UyN/fEPv7f/8q//l507e8bu3r5tr0cX7fLlY4oFd++8tn/8j7Blxu3w8RMya1+anhUg7PqNG7a+geRrUgOiUiVvp947YkN7++3K19/Y5MSibdfU2jb7N0HD16XeqJc4E5A5uXP7tga1PNv3T78vs3rkviITmHxFzXk1lGHzewNTuQQ1dW3Wjh05onONerZYLgj0Qz4QGZVIgrKx2JPEMvmDBf87mn+s2bm5ecU4oY7F3PL4F0E9GuyqlsJnwxHUUbZSSg80KoOvIrGV1+A9yPfiCMMR92mPjTDQidsYKCeS+nmxydgXKQA5ZQfBBJSdct4ouxLAYqr9tqvW0twk5gd1ZCZT4x54NUnb3dlgh4YH7P6jJ1axsg3077crf/rOzp89bUfODCoeFtfL1tHWbbdu3JZ/wce//LnVNyFLhC9Tq5VW8/bk/mNLN9TbiQ8u2frymo28GLXJ6TlLpXNiDuKD5Z5uAN1qfThmVflXSQpQrASXfeH/qI15XnweZH1Yr7CCGhtz1tu3W8+JGAAYhv7N1Ntpe/z0sVg47e3twfi33sEEQVKa+8xZzX3CnJn5CfXK7PycckSeVx3gjbUNm52Zd3agpFlhDPqZpia2GFc+QJfErICRTuHxAQVnjgMRPceJe94HH5JqC41gH6Y6C1oMdWor5XXOvueZe9M6JcAFsYFYr75SqaRcFz8aGDEHB/ttZW5ag4qb12/bBxeP2ssXL+3ChXN248YtO7B/n92/88jOnXtPklD7D+yzRw8fW09Pt62v5iVTWU0mbD2/afUNWXv29LUNHxywVy9G5bd287sbduToMbv27fe2Z99eWy6U7MnzN5bfSlpTe5etrBclu4nUYD0ynjUmRjdMXWoh1e3hXgB45HxXvSxli23VnYvLizZ8+LC8NWBJwybgHuGj9erlS8lCIevHfmTPSgGi6lLEDib60dBXgDKPtS6nGSTzAktGYTSaOAdgGgAz9rD3ZdyH1pVNAjhVNYDLwUYALusrMgactQHIZkt9RAblnPWcO5zxxDWUDIhTkSEHiMCBPl4hcgZFdmUEd6g2CuwEWL6KO4EFEuOPy2QmVYu495rXwuwBPgd5QRyQwurk/RUz5JOD4gpeXTCnUUrI7tQVOs8E7iSfK+rcBeDGPuYz8XmjjwavGUG6LgXvQAsfWriklcevVBjwuGLFTi0Zn81Pg4p/d8b/9B9/BXdgVzIVGj7eRCKw7Nm9W4mZ3OnDgQFqFfozicbU9JQj7kslJXlsTJpCNNNAQQlBK+10n5yrWYzUUNCtk1lPaCS3Nrc4+iWgvUkKed0dI2zJMrkunGRSgnyG9K8DIoiGTB6KH6+r6a9TIdn4Ec2rAlqofbNK0ColkUcrmaSfuTSJO4EbIzQ1ATZpwrqsDyg2pC04LBWIa5zqBroPVBJBS4k6SGmCnIx3OZhJfrNq4FDo0LDjwBQtFopy8H1QokbD40cBUJIZmP+EpJuzgcDumnWgN10HT83bYPzF/Za2I81jmlUyuyU59En4rp4uoSLV7AZdnvLJN9evQQ5+HGLFuC4+MhSSiUiDAAfB6JRooUhDhhgnvfG5x4m1muPRKDxMtoWOEILynW8FE2aQfdLn39yQWacakrVZW1xY0jXSmEBOg0NDlNdgys2QApmr8fE3erbcDzF71HTyqfbE1JR0CIV0NkeNg1iTb0P4ciSNfyAM82jm8dz4FibcNLVAiKlBTqNQE30vhmhq8WfeU+bt1W012mn00uDgWnU4WsKampq1R8paZ42eyPH6DKKCZBnr2t/H35uGmFtd+6EsBDvrGCSDtPSDRmL4LNwvN2Jy6TRvfjMIcbk1MQICskWH3498RiJlXmgn3ktGdUGJTb+7sT37xCVSXEua9YQmJAmzZCjqskLGs1fUiAsoOB26klXIWltLq22peZvWfWEISpxh/zNsUuN/fV2SC+xrGrDcX94Lmm9EhdEIgMJJArdVLloamTpklTbWbXurLANlNW+2t6yjq8u2EzWWL1VoY6oAoLgH6Vtb569dy1qnSZ5IKeHj3i2urGg90Vjh3vIcoP1iBgwqkn2uBBC6NrqTm+5JoaEpetJ1WZkOSiu5WFSs0rArmfLESvqXaTVaXDseDxySevfV0WcOgwmxD4LpOw1KDWdLW7adqKroL9PsRF4klTErJyy57TJrFavY4vqq5RqzXtiLOYbR+raVi2XJYGVSGcX9OBBjsCKfGwo/NcjDIC0yjYJ/DH9PgwPEZmx8cF0gYol9SELJJ0HoqBolZ2JbEGfC50M+gPdpaGhSjCHJdr8Jlxvhh7kW9ga6ussrSy6BIwk7BrUuZcA5EWXwHDXte51YAOuE5B//i86uDiHAWcc1CTe9pYG5srRgtdkaq69P2/mLZy2TzYh5g6nlZqkiuYbpmTkNpzBd72pvF6Id/wJpCqN5vYVngRsW+0DI5aAickYNQyXuBRX/kifYNmttxGvDdK4sE4cxmKyU3AOpUpH8kHvyJK0WA1gN/J0dJ1o4awN0nRrbtUzrd5CErCViI6wLb9yUpWdMYfTtt9cFOKCw/7vf/50kligKOadAlvEcc41NksgiGSeksWZh7rkhsKPeNXg2s4cP7tutmzeE4mMdNDfBKtxWrnHy5Enbd+Sgm8aBRsXwfmrOrl//VuwkhgG8FjIRLlHnRsNvJ99qmE18RIpo71C/vX/yhJXW12xtedEqpbx99dVVu3T5jIr4F69GbPjwsKXwjElnbXZhxRLIO6UyknBB+7tb0jKbkjwBVYgEC4xSarMy1HlQ8jUJ/Xsxj/EmBtEtygcYWDx7/lL3yNH97vHBXmzONVgjw4/1dbEUqjA+1BR0ZP78HCj8lFCLQvuBTGMghYOOdHm37dTpk/bwwSOdgf7abpzsw22X9OFrfbMo83O+B08E4gNxeTPvxW1dPWwt3xPIgLEWBwZ2S8+cnKi7Z5eYJxx2sIdAO8N04PPNz8w7khHWxGbB6muztrayZBfOnxHCGKkcQCivR0d1XSBslb+VnbnK18zcgorq+nrkdmqsHvkPGadWtD6If+x1l9KrD0Ppsg0M7pHUmHy0atIu76ZhVUF5iudcfkZFpFk8z388qCCPIHZyX5xR4oNY6fpnaOpu228//7XdvnXDJsfH7eLFC3bt2jVraGi2hqZG2yzicUZTfF15LOsZ9gf3EkNoN2D2poCMnhke4LMgtgZyCg7Q4bNyTtCA0BBVKEFM3BnMOGuM2OgAAzhy3jwUEjXILcgrSHIk/vk5J7hn8pgKHjkuw+Dm4t678vxDLJ4khbXnbzS72EvEP54XrCYYjpzZ6RTNe2S51uyDC+eso7XVJsfHrAtmxfETaiAXN4pWk0lLgnNhbtp27erUHpyfGrOpt29saGhQN7m5td0mp2bt3sMRa2vr0T5saesQa6W8VZbkiwadNSmBoHp6+uzli9eKl+5VtKzYj+QpQ2qXcdjUYE5SV0srYsO5tKtLjJF7gYKkYUYTaWBw0Lo6u+1f/uX/0GfnHOYZqelMk4vhRAX/HoYdtXoProfhwPzsrHWSnzY2Wq6xWaayNN+UX7FXqxU7Orzf2loarLWlwSbejNmzR8/tv/9Pf7RKsaBcHVDUlavfWteuXhufnLKl1XXLIAGVSmtguP/Afhsbf2MvXr2ynl2Aw/L25NEjDT0uXkDvfl0Amt0DAzY5MRU0tEH6e20kfyv5BOStUi7q85PTNDa3WX1Dk02+nVRzNMrXUp8AEHAmEEP7pAHIYADc17dbchT8G7lz/55BG8WElzNDRF/P3QF3KfcLwzUpzoOkTiZVE0YBtuaGJlteWpaMJMNc7Vfyrq2yTc/NWRJppjD2ohklLzM15WqUc6TTSGb62SJ5jyCrEcEzvJ6kU8NwLrJZOTuIe6yjWFcJ5MI+CAApSdnAEMi49NPE+LhQtb0wG6dnFOM4I8hp2Z/EKvIz1uXg3r02+WbM5mZmrZU4sbZq586+bwvzszb+5rXyG4BX//if/sH+8z//swYVyMlMTy/Y+fMn5Tfx4OED6+7aZf/1v1611tZau3Dxgu3Zf9BePhuRAe62Ab4w2xRgpGT9A91Wl8Wn6J7Nz2/aViIN7dtStY7E5QvvHdQP8NRjDbD9OSuok8bevLHZuXnlUS4p6+bwbpjrTfyYX/ODDNzPnjmreMm+glFBXcu9Zfig2hE4eBhU8Jn52t3fp/OGuosBtNeOAS0vKaBKyBO9RmeP6BkSOzOw5l06U3VTYM07rs73nUBoQd7ZJWuQ0fS8QYRAnaUe82AYMawRCln3wpka5I4uY4MsF3KC3hCUTA2vH0yEyQmbGnO2XoTtm7WPL52zE/v22OwYElqb9mjkpeXLGzY0NGw/XLltXR0t9rv/7lMNvgvrRWtuaLVbN+/YRiFvFz+6ZKnalAbyLY3Ntjgzbze+u2MdPV32wWe/lPfO8uqmVbbJP1sYR8hHj3PCWUWet/OsiZ1iQXEvy8404M8AopCVkWKCvCLZo9u2CXtNEoxl6+/fo5iA/x73mmcA4w7w1KHDhzWY/erraxqY/v0ff6dG9517D21wz247OHxA+cHe/fvs2++/U95EXAFIQPpJLGI/I+PKgNLl6WoUWx2I5yBCScTCfqhxVohqb2R0dHa53n/Mcfg38iZel2skvkVFDj4PMZCaSuA7vjfH8N+Uz7ikl7NdqTGILbx+W0eb9u389IQdGNht60sLdv7UEbt5/YZdunDUnjx6Ypc+uGg3b9yygwf326P7jzS4AICzf/8+u3v3nnpl01Ortru/S6zLrYRZfWPG3oy+sf7+3Tb6YtQunD9v1679YCffO2nf37xjQ4eGbW513Z6+GLNqOmvZhjabnV+2/cOHbPTVS9UglUrRNvIbGh5xFiGNRtyS5FI6reECw0y+yCmQvub5HT1+zB4/fizJypXlZWexdXdI4nf/vgM2OjqmmBbzIPaO3yuJ7zn7MgAS1ZPDb5BYrnjJ/vM8Q+DiOgaCDlLi2iIjJ0oDqk4NoAn1+xh0S262Tv0/vp/PI/nJMBTWAIZeX94BkDxvGFkaZhSdkcqXAzNdlk2MHeBIgV0e2SScoT78rCg/Q52DepchCvGe+8DnFiNHvoruLQnwhhyN3tW7s8J9Hol9AnN3dyt3RqpUazSwOdWjDL1R6gjWapSSYzAhdk9+01leAWADoyKyypQ/43kahrjxnPLBrKsC8CDI+3YU1gLIOAJzfmJUxCrgp9//au7AQDanQkDmzAFB3dzYJI1dDhwSMzYkTVQ2EVN5EBlKIra3hdCB5umU2rSSXgIMG4xmCIGGJh30KBIgoTY03fRDSLrcHR16H+n403RBT1eTVy+21HAJXxGUz/tL+1gSFy7DogQm6ErGIYX+cttUJHJgMnGHEs71EdCQjGKCT0MZNBtfUARddsaDN1+OOmPimdKwgOYbzQI/BEkiKiq41DTj0Mz50IQDnSLK/SCcbuwUO0eYEnBonklyJdD0/f18mg1KQBT+kITzPpH5wHXT9Iz3OQZxITyRehFiHrSm0/8pwCj0ZHYaUYjBZ0LDnaDDJ9SRgi0GTo5qIEguLYF2JiiHhDPC8MMkm2RDqNpgDBvRS7yfX1swzY7NdhIYM+vv71NTA/TN5sbajoagaOkyT3PjYp69kBJZqHeenAo1g1ExU2tJXzl6nm8WYjtTa8vra9KR5jUc7YwkjE+i/cuHFJFerP9KuIeFJGx4XkEaTBpLWdUAACAASURBVBR7TJTDmvQDxtkoSFLRyFayLKNcGgnetODaWRfIUznix1ODePjIHClMxyXlBFMI3XKhQvywBj3NoRwTfj+sWJPeyBbbKJhLq3EZjJbiYRsb3D6tdwTBO91fl5Phf24+54wX7kEcZLCeuVXOoHF8u6QsgnaiD3W2JIvBoFNIEO5BBbNhkg5Hw1AtyPQ5kRRSl31EsgSaGsQqRSyNLJpSIIG4NyRmNIhAQPP+YmIFo+YYaygitHcYPFZKkn7iE66vLrtkTTB8zdbnrL6x0RYxyWaoQjM7sS3vBjUEadhu5qUvu29oSLJhNDBBZ/OeHe3tbjwa1j+SHwxTMAXGFBa0tMt6+ffTVENmiAYxz4VYy4BDVPTQXKKZxl5TIU3BFZpLbnLuBtlCb6jg82f7TsoECTKStoQl0gkrlPKSe2IIkrK0/o0kS6+f3LLGFtcfB8XP33tzh6Zlg54ZhQtDBxIqqK18aX2G1RKbgNH/xosNZ7r4INfZLdIYls76O8SeaL4h4WLQRMHF/nAarqmAQ36I63JZANeW1r0s05z1ASqFlGQ9VpY1WAV5LxPk6rYQK6xFDXnxMAoSKvxOAdeKN0GQW5qbX1ATlOEUg0kZgDLoSZSts6vVzp47ZbNzM1bX0CTZj3WS3zS68zDy3KuDwnBlEYPnoi3MLQrpCiOAhJXPqIQ7DDdp8vOclIiC4KEIQN6La0TiSB5N3kUtQFtnGAF1GYoD549QYTRwqpZGg7dUdAbZFoNnl/nKI2eGv1HW4xExUXR8/CKQPkD+KZWS2SDDV54xDRqhslMpoeybm2miYRbXYF99+ZUNHxq2fYcO2XYZKUdn6ikxpulXKCnOUqXqbEEWYnTUvv7yS0dqVYmXGe2b5aVF27dvnx05esQSqWDMV6kKQX3//kPpyGNczL0BRcq6o2ElVPVm3upydVonmE7bVtmSW2UrbWxYX0+X9XS127/92zd25NhuO3bqhK0gA9faLMkF1NIXV9ZtuyZjG0hFZXNCbBGTaNaura67sa6GarAdktqvjRh90iBQk8TjFmc6xQzrBt8bNOuJkUIaV3xgiklmQ9Z9q2C+1LAvyshLpSQZpXmSBtgea8lFxEqsejNiYxM6+JZQsdwDmj6sG3IwoVXlN+R5Fu/hyDpM/wrW3AqK0odiAAzUnEnC5nNd7levXwsZyqAOfwEGcRouahAIkSxKIzozrMCAOA2Lcc0R/pm0Bqholb9+9UqDAxo/3vD02KR9y/oglmsgCcjC/clciiMp9K2kyWA5SOqoJFQ9jSMQ/2gNLy4t67olxUNDXabJpmYWDXc/p9zQPp6Dzt50pBvvQ2whP5RUIw1SUPnptOVgwhVo7Jbs/VMnbWlxXs9m3/4hSZXMzS1aR2en7gfPjz2MdAq/08wk96WhKxNsnWOwQvJqMnMWRZkddrubRhIfGWqs7Jhl05RhQMM1CulZLklaQ4OVrapYMbxePA/IxXSuasDvyFOXvIGt6xrg7wbZIccOzDfJFeTz2j/kKjSuGGy5tEGzFfIlNQO4HwwcGpvqLbFdtQ8vnrPDhw7Ydrkk35lcU6O1tnVaKunMA8AlVq1Yc3POihurVthcsc2NFSGwO7o6hcJ/+eqNjY5NW219s43jV9fTp+EejQnFEfSbOaORcSqSNznTSKxMScFimu5DOjWm1OhE1s8ljfh7DOu5NyB/iXncl5WVVevZ1aXzmGfA0I+1IUYpDVQGaHV4UXjeTh5AI8Ub4khwpayzvU0a5+ShDDfpD0kulvoAmbZqxY4fHbbdPZ0a4rW1NEv2ZX1lzU6fOq6clRrgux9uWc/uPTby4pWtrIFQp7m3oYFKb3+PhsGcRwug+Ytl5V4ocJ06edSWl+dsZWPNho8csdevRgUuYCDO6+KV095KTkI8YMAKo47c0uSJ8WZ8Ug1oNYVqa+X5xPdSr0S2LOvv/v1Hit8XLpzVvmNPzy8uWqYuZy9evJSHGHuBPes5rg8IOM44izmbQEhL9o2mrzzzYK7gXbCmpidyLYVi3og2yOFVJDGLxGWNA6sTSWtrblOMJTr781floPsdm2jOPHcAjEBP1GAhBjgohtzDpStjQzMCi5TxB880nrUPPDyvRuKLdYE0jvLMWgezydi9WhWAgMYWe4jhY1/PLkl/ETcYav/88kUbfzNmbyfGfXiUq7d/+Mf/YP/8T/9sP//ZZQ3wp6bm7czZ43bk2BF5Mq0uLdm317+316+nxWS6/PElgZgePX5ia+tlw86hWEEKb5edu/ievXrxzF6/mrBUqkGMGVryqSw1KzJUrjMvcAb1i+QzfYAHO+nx0yfyreKzyOtAsnBe3yijV9x0uS3YhPgoHD+GsfAjsX4Ylu3dt1f36PXouNdilS2tCfYKEmCspT0D/S5PVyprkK34FxD/nJG+Px3dzvklz0v87vDzA5gVBkqRVaF8W0bSHtPE5g8GueTXcTjv8ZG80c3Xea6Sw1LM9iYlZySNT84BhmduCO9el1wi55uY6pLRcv+V5uYGW1nzvPIXl8/buWOHbGtz1UqFNbv76IFt4v/Y3mP3bz62bCplf/uHXxiKBOTf7XuG7Kt//b9tvbBpv/zslwYOgwYmA7zZtzP23Te3LV1Xa3/z+88VK5+/HLOxN9NmNTT2MTn2oQ5xz89+71MgKRl9Bsj98CYi1uzq7pLHBOfNg/sPlPfjXUAN+f0Pt8Ty+Y//8I/2/Y0b9vTZiO4L/lQg8cmJPrh0XgPFq9euSHbyj7//rY2MPLdHDx/Zvr17JUf5w40f7LPPPrN7Dx8Exlte8ZuBrPdhPDbzLJGsnJdkHp4F3gzXmczwzcn8DuxkuC8pVkfwi9kTwB+xsc66IY9lUMi54zWGr32tnwL1uQM8I7tbcjr0BSRHHmV1KpKBbW6ot5WFWRvo7ZaP0HtHBmz0+VN77/RJe/30qZ05d9a++vKaGG03vn1qn3xyWvfiwOFD9vj+A0kDj72esb3799j03IJyvVS6qn4Xg/rZyWk7euKkXb/yrR06etS+vvqDDR8/ZJvVhH1367GlkSVuarexyWkb2rvPJifGxU7kFgCmQloTIIEM5AMzk/xSkkIJB2iQvxKvARAP7dtn01NTVt/gtSw9FfInBhUDewZUnwo0rD6YKyTAumHPKz8JIEjd+/AcXE7SQaeq/YPELU17SVwL5e+Sb5I8kjm2e6v4kCqAbArE4gikCf2XYGbPM/NBI+Txqs5tqaogzQcIEZm3AuCOrNc/ofexg5ZFNiAyVcMQmp8Rw4M+IbFDbB0HsvIarviQsLa2th0PCPJomMXksvocAvp6/cbPyt8C+SqYXzu9OAd/skYZFrGe+VlUERiG7Dwn+R4BYiYndqNtSRWG3l/0+4hga332sNfjoMKHRT70if2dyKiI3ayfBhU7jb2f/vDXcgf6UhRObCZ1dtUwBqVOsGMjkZRx2Ei/raVVJqNMEQlEbGCaSiQqfKGrLoqdJIegRpP4J9RYgiIYkyHpmYaJIUEXGirJJNPGiKgmgJCcsOGjeVocPrDROXQYHCiwBY1RisNY9AhNpoLbPQkIgqAbncLlE1sQcUg/uR2Ao4SE3q9zrcSSpqOmBiroEYIKyDruF4UkwZn34frf6Wyi+U+B7BQtmmgEMVAr0JmVhAnF4ok9QUnyT/IJcbNdki0ZT5F01maECOOGMXllaOEDH17HTXBJuNysE510b9DzWrHxzjNw2rNTNHt7enTdNA5chiA0zkBgQNcLyDsCtpK1gNaj+UCyCaqTP0dtdGkEqokdofe+OyJlUL4h0fguPLPoBQJre2iwX8W4JEmStoP+5zV5Nhwe0qzlgAZFWHUkJX8vZBwIrdBYd7NBR7JzGNHoG598K4NQvwHuQUKTKQ4Gfjyo0LrkfgXEueh/NIOgtIf7GKnIrFclzaJL+0GpxmUwEI/yABqCyEMk7RriNAwKIIlpVGLQnlQi5zqvrufI98Mw0HtSzCMLBrsnrB2u6cesDhICMY+C7q4St+AFwvvR+BWDJ9CruV4a8lHKRz/HwwiDitjo2VkbWim+VlgToChFS9aQxJksJCEgF3r7emX86IMrR3rxGSIaQIwqrb9NyT/JxArt12zWB5YMN1RguKQKBTXsDPavEK1lb1JEz3k38k7pujypq9XwFBRKLksD1bXmKZrq6qFRJ629E0mPsq0uLwv1BjKctU9cELqZJKYKMienZLGvv99+uHXD3kxMSLf60KFDMgGlQGbISXN/77799s2339rM7Lw+Cw08AiFFCMUGg5mIJFlZWNIANkqfOe3eB2x6/1CsaZ1DH6VUD8mWr19YWXXa+8QPYrASSPZGTUJ7hdq+ZpsBhkvQYb6ZyqYsmULqCKNwL1RpdmAS69fiKEl+Ra1Mf+ZOqY3NvtgEjPtaNG50QOP1BHk6JbjSVHWUtSPfQLQ6EozhaXt7h/6bvS1ZmKYmL1q2ttVU4Ys9QpwX8jHlEmpIK6DjLd8f5ACUfBMnN7THhO6rQv8v+nqA9dfYKNkWN2hd0frdquCZw3DIrDaF3OCGNTZmraExa7W1NWrkMtyi4V2EucJ4VfTxitawnut2VecFzT4a7awLvvBUkTxBGEBRNHCvImpGqEYGBCSvqbRYV9xDDVqRewM1Jy8TN0rzsg6N7KKlMjVCv7OOaArRMU/CWAnNB+05tJxDM4GGrmIpa1tDlFoNRijEASasr67rfEfPWHOjZEIFPXTxn/3i55INkNxL0Mhln2mIBIOEs3Mnsd5Wc+Lh/ftax/KtCD4dAAaQBmrrbLOO7s7AGKvY5OSUPX3yTEWXMxC3NSSBxTE19VbrF4R/165doTlSEso4m0xYcX1dBpJHDu23L7/42uob0vbBR5fC0Kki41Ykn9AAT2bqbGUdtlNCBoSYgrNohMxeXrE0Df4tmE+wntxA0E09GamHxkVojtK42yxUxESiCdAIo4yhbLpW9wLJHEzAacLRaV3bWJNRfBk2KLIsSHJsOasJ5gCNRGcybUmugAUJKgskGAjCyAilsc0+Jeag0RzjA/kVwIZMrQ+PhdJXTkPDA+16Z6GOjr32JisoZYZgMFTYJzAUiLk6cxy5BQsUNg/njkxwAyOS9QtSkAKY4izKq8AWjF/cN2KucggYtgGIwr9HFp7kXQQA4WysF8KTmFsTUNQ0wKI/VU0aBJ4z1QC/wM4hLnmjyY0GHXDggxnFydDAiLmQF3nenEZPH/Nfzq2B/j7Jy8zNTAsJiZQV7IXGxmarra+zuflF7eW3kxOKw3hpUaR3d+9yKdSgf68hSWAo8lz4/LHhqTM2gIGcIcGgIKu1FzImaThLijVIOrhEqKNNeQbucZZ1dnHQ6Scu0+zmuiQtF/JbzzHJnf49C85zFfe2YL8LKYiP0bb7PRBhioV1yRYxvPmHv/+97erqsLWlRcvVZfXMUykYW3ViPTGoAQVaLm5Ifq1S2rT19RWrz2Wtua3Vmlra7PGT53b/wTNraGq37URaTW9Y0JKn01DA2Tgyd5dUQ1oAKoAdNFZ5NvsPHJCHCXuCQXA8Gxg+aNDHAEtyV+79BEOCPcJa5V4weIetRxOEOocmJXuKJiqSVv17dtv9+/fUXCYWwKAuCZGbstamJjccTtbY8sqaUOIMMxlSYKZ99v2T1tkGO7GsJnVXe5s15JBB80F1Ipm2K9eu2+C+Azby4rWGpdzD6N9C06dvd5+zGN5MCGxBHE8nq3bm7Hu2ubZkC0vzdvDIMTFJ+FlJ1+UBS7nWtTeouZfkI2FNJVJidyJtxN7k/kRGEay72BBkfzx/8Vx78YR8cYgVtfJ3y9Zhuj0qthsSTcQHl5xxMI5kLgM5GRkkVmupVLC6TFbXg4E2A3zOvXa8pFIJW9lYF4AoXVcvU23lkEhlForW1NCsJiYNaHI04iF6UAJKqNFJaPLGpBrXQWLGpSS9UUZc9bLG608N8UJ80B6UGXtFzChiCDGHuOqMlLLt6t4VgFAuValGcaUiaTKGCDThuR4GvawNZEYX5+bs/Lmz9vzZU60B4ju55R//+Hf2T//zP9unv/6Z3b97x96MLdjZ84c1fO7q7rRjx08IMDf64pU9fDAittvQvgG7euWaLS1TTyQ0jOBM/tVnlwWkePnyjW1Xa62ayMhrrbQN4MQZu3xQhqQgzF+/HlWcYT8cPnxY5ukY1XMPJKPCQFkx3UEDUSJFty5IgR0/eszu3rvrSOqtkh04uE+D/dnZ+R2vKx6K4hjndkO94hHvyRoCOMJ9IxZxL8UyD81H3oZzz+sa9/+LgEAf3Dtzgv5DBOKRU+48d/LqdDBOFwveZWjJ/Xn2nGvUQsRMP19JB1y5wGtE8mMfiPpQxM8mKRakGARmrb2tWfKAcwztapP2q4/PW29Lo+VqayydgD2/akmMdfMVu/blDdsq5u13f/ilclOYoqfOXLA//z//ZtuYWH/+S0smaGQvWFtLuy0vLNutm7e1zn/9m8+tYjXyJrl157nhlVgBdKWj2GszzjqGgWIih/4IdRx7H/YMawoZWUAEfAbYAMSGs+fPWL5Utpu3b2uP/PY3v7W79+7Z2Ni41nPf7n57/nxE9+HAgQOqLaamJ5UD9fb2CeCwubah2NHe1hYQ4c565QyjsUsu5bLR5NO+PzVE2kIGclPxnD4KcVvyWwF0RQ7A0El7NwwyfNjuPpesLcl64T0Cwr5cEvvdvZv8SzlaaKRHnQRqUZfyy4jRzXqODXd8EPFwAfBSzq9Zd1urVfIbtn9Pu02+fi2JNdiVp8+fs6tfXLHhg3vt22sP7eOP37OnT59pyHj/7gMbPrjPxsen7ejRY/ZydFQ1ej6/pjp4aE+/zc/O2/H3Tkv66+Dhw/aXL76x4ZNHba1YsdsPRyyVzVlNttHmFpdlUj4z/VaDI2TcVlaW5Svh57qztDlzeMYuNf3Os2B5dVW9poGhQdXeza2tOu8YPCHnRZ5IrHszPh48R6hZfF3Jj1UARx8CqvcQWOiuOu19tIjsFNBKNQ8yTS7pTT4rI+4AvuPvIzMp9mJ4zZgnRp+uWMvy/ZEhxTVQW/NvLo8dz/Wq5HldAi74jZDHCEzpZ4Ny6jDQJJ+gx6Uhj3qAyPW6nLZiOoMCmdI74521wvr2/NHzBb6ktBKMxunv8Hljrh6BedSW5CWsba45SkmJIVIqCyjJn7mJYhvncjvnisc/P9+87nW2hAP1HGzjPUFXbfkxs8zbVG4mHgd7Pw0qdsLCT3/4a7kDfelaN13mIFDhkhM1n4agF3pOmSRpZ+PQ3OCQ9Q3tci8yEg4sAdBMTNLZkBS7PimvsbfTU0pEhcYN3gRePCZUiNOc4pBkMELTnuRKzS816fxLU80wdeVHPQD51DYi6UkoaSALucf3x2a2pG5AwSJP5drGkpSgUJIJt9NJCdyuW+mHA/8QkzoKOg69KEkSJ7IEJ+4H947gDMqXYEWDlSQNtDKo1WTCp7XRSJriRE00kMWSevGmI8E86ozLvCtbpwSMgEkhp8kwqMbarA4nPg/JglCX4cBG05cmEzI0QjeHAo7nSqIBSrK3t0fPhPeNSANQoaD61LAEoROMiJTEWY0Q7SSpGhCkg+QISPyAAJfEUKBWq2gPBnhiugQU1DtkE88nYa3NTQFlTNKM14hr44thE7rRoOy4DwxFeN6u94zslq8ByVjBKJCPiQ80JGtQ2bK1jQ1bWF7aMS+VfA3Jn+qYOGR49xkkoxUGaW6c7Z/DDzAv0jhYhAISSgNkJ3sFND4sJP9vH6R4k5LDsTGHP4GzLTaLDAGbtU5JJF1TGjkG1/ZWY4+GdWAg8T41aU+oPXfYVnLBWtHnlbG0m1MpcQtoBOm4Blqz2D56PphG+9SfJiKDNh2CkjRyEyd+SVYsPDOtw0ARdlYQ/UnXeZe/jKRuanWAQzHH04bXQOLE9dVrtS9ZP86woUlUFoouNuspJmhcI5XCNbm8wDuqNp+XphAxSRIraEMKjYveNo0b0CxudAVSnHuNFw2Nro7WJr0PZs28B81Y0PU8w+mpaSuUCioW3GgyI0Qs0EkKZzQ+aaBB3Y6oEdY4aOeW1jYxNWiucl1Xrl5TY4XYIlbU1ra0uGtFXaUhlLSchjMMGh1RIUkXpKbEEqHQdNaBD99ApIShI7mimCzQUNHXdekKR2QwrPG4Jbm64BuQrkGyjQQ37QbS5YLlGuqss7NNxRvxgT2DrMrGZkHMkOh7o2YozYyAbPThkRcg7KE4KPH15nIKfEnqBNRyaMCxphQzhRpGioZ7UXTJq4By9gGbNx0jel3yY8Ro6Qc73dWZJR77+bzsL31pwJKyfMEZVWpIan9kxCCIxm0gjfBNoIlFIUAjEZYVmq0M0ElcM2mQ646iw7ibvcZgABDrlsxMaIKh3eo+LBFNw+CHZLhYKIvxgXEhCarQiwzC0RDf3NiRglMsV7UA5R2db2QbaGBHg7SElbZcO1nIszD0r6GJB5W5pUWDCOLh5vqm1bKvmReL5ZUUoyJSqYUyDMwAzvfNjXVrbmmydCgoabiwF2hyURxNTIxKApHLowi9/NFHdvDQsOSKBCAIBofPR56r6Y85PDJANRigbmxIfnBlZUnrcHJiwuUhKxWhlxYXF2xgcMA6e7pdF7emxsbHxm3k+XPJKkkeMZ1x6T8hezPytsBo1zVeF21xflamtduYsa5v2NnTJ62vt8uufv2Vrayv2q8//9SK+Q01ULeqCVtc3bDJmTkrMVdJpeUtceDgARlTS2ZraUnGyYtLaN/nhMomnuzu7dSgqam5Uec4yHoeBs2eYrFiHd19du/hE8vm0NB2c3f5EYW4Ri4kfyVM6BtylstmbP/+vfYi3Deo+Xv6B4QKh5nFWgco4Q31snT5abZwfQAWGPT4IDEhlDIMHR6SzoFUSo3nxibYIs6E1P5BJkKynil5wMzMTLuZKPq+IJolo1erc50CnnMfuSwGUeRh6PpyrtDglbcNrJzqljzJhg8elGE2awdTaX6GuMC+ZrCMpJ/7InkOQr4DWhPPKK6ZnIniE++KaIapBn+laH39vfbixavAIjHdR9ZFRNkrDoVriYwEziGtqeCpFM2VNdjX37uvF/KR7JdSgWK0akePHrbF+XnbWF+zEyeOCUHO+zQ2tVilXJWUGmAQgXqSCTUCJenIWc6exrNA8kne5Iqxj/ckFxFoIOgr+9ALD5g6W11bFZI+Ns7k24A0oHyPiiFndn8wPmNsNrMmaYKTW9BoRzqTZxU1jD13ChI3oACDaa3nDTCgXO6FvDn6lyQw5q1iZLlpnR1ttrq6aLWZpP3i4w+tu6NNQx20+Fmr2bqcvAuIg5JsXFm29tZGSyW3bWEW9mpJ0hAdnR1Wk8rYk5FXkrwpSHkjrfXFecpzICcH/NLU3KrzHc+qpaVVPS/Wh4YyyYR8FiJjem3VPawYmrDmALqoEZFEypE82pmaMRci3ruOOgMdznXitg+Y+WLttbe16oz59NNf2jfXr9vE+Fs1oMklOG/QdMfcVpI3wViTI7ec37CL505bbRqE65Y1NbiZNvXG8PB+Pff6XKP96YuvbfeeIQ0qCpWKZbL1un8MkAFQEKPZo/JeSiRtaX7BcnUZ+/nHF21lcc4WV5ds3/Cwzc7MKa8w4/l6wyWHXGKpoGEiMYBnzOCUPJfBcBz6wA6IjBuGeOQ3rFn2IlrsnJnImzDcoAk5i1dhvqj8B2mTAkAQyW9qBrHjI+A5TN5S+GnV14lRIUDa1raAbzNvp7U/uMfLy4tWYt/SdINlTv1FrGLgXa1aQz01YElsQW90MuD7ccXtQJ5YczC0iGA2b3b6M42sTA32QNXusFS9fmAtaR8jhyM50oxyE+47a4f8jlxNLMhUUqxfBjfyh0okrKev18bHRl0SNmlWX1trJ48ftZGnz2x9bWUHSPbbv/2N/dM//Wf7/POP7N7duzY1tWAXL5226akZW1yct199+ply+PZd3bY4Ny/TdNY9Uojr62VbXS/r+c4tztpHP79gXe2Ndv36DXs7tSr/JQbxAJnI9WGhFQsVGz64X2zAO3fuixlI1nji5HsCGWLSi+SYN/ScPS9mmoY+zrAgTyWOktOcOvmeTOfJOdO1NTorAC2yhyTBG1jnMlVWbUWemNB5sVEo6LkTN+OQbHPDJVm8qem1LD0EcnjilpiOAYzDGRjPNv5OnnBBykuyuKWy4o/YJPQciNUZN53eQR0HkE/0qAwYfh9KIa0XpFSjX0X8b9YSsbuztUXScKsby2ogf/bJRdteX7Xa7Yq1t7ZYMpu2rv5+oGS2ML1ok6Nj1tkBaKGi+//h5Y/tq6+/0Zn0mz/8WsPN2Zlpa21pt7WVdXt4/5EY/L/87FdWSabs+tXv7ObtZ8rf8EeK9hO6r8FjU2A8gJgM7WsB1DAsQPEgKUN4cjGGujAeyan79+yxQrliM/Oc0Rn5TMxMz2rg5g1U6lz3ByFnEcJ+GwBZSpKg8rKBJYpHZkCT83ewzSUZubGh9xG7NzRs2Mvkv/IaDOxGfnZ1ZdVej405kCuCAgNAUA3yIAMlT4DolSCvpozV5eoFuPIhlue5MA3Y695wd2YVa4Y1EEFM68rngp8edUKe/kevYraV8tbW1GA1WxUb6Gu2iRfP7ejhAwLonD13xn747qYdOLjXnjx6Zu+/f9Lu3r4r2bbvv79rJ04ctKm383by1EnJX9Y21tvy0oIY8709fYp7Z06flmzWwcNH7Otr39jxM2dtZnndvr/12LKocGTqbRX/no5OMfFamhu11xi2tXd0Khcg2K6vrlprW6sGDfJfhakQWDULS+6ZRu2NfCCsp9fEprQDXVGUgFGB9Bv5vOQ8A7iD++a+P66YEIcPqj+DaTV7QbJQIbZ67uVgLIGRYeLjdxWmRC6T5PKU7FvWKD9Lrqm9HwB41ED0qVw23etgvlZW1xVD5L+lGtiZx5zx9Ly4fs543o9zR+AEMcAbNYClJ9bYluNrSwAAIABJREFU1OznWwDLiRmcxf/D39/rVfezlQqJhgMA9DyPc3lNr6354vOR95MzqUeACgiG4UHCl+fE5+XsAgihmi+oiTjjy71FY/8QUBHxTIOKoHryTobb1Vu85nX2ILHR2STOUo8SwHEwo74HoIifPCp+nCz89Oe/hjvQn8kqiSWog+gkqGBSR2IRUbJC+UkjMCeZosnJiZ3mGI0HGuguJZMQSolgoCkqQwkCGzTZzU3XqJOubmh4BQ8JXoMmpqR7ArKhvaNdenqSBwiJIfc7In150WicRnChGI9FTEycVJDKvBXZpmqggEFRTYuiD7qKotsTbh92eCFHQ6VFKGwKFIIVTTwCIcUlgWhxEbkslzaRZ0ShIM16rkGyKrUZNa6FIk57Yk9S5VNcZ4twWPKLIpOilIOGQ4NrIIFzCliQT9mqKqmmgcKhQWJCM4ihkZucuqGi2BRBC1QNzmAG7b4RjjxX8C1v7fiLeJ/Pm2MksGiiRyQkf8916fqLJIaYXCMp5UwH14d11CBTbXk/UIhz4CkBcjRE1PWPSEdHfCatLoMEQ22QBvLiQ8FdCB+3a/Tn7rIa0kgNwy9PXMvS1ZdmYY0XKTrcQrOOPHyzVJSJnOTG8Njge0FQB+aCK/j4kIRrFelD+rsucaTEnSZqkLfxyfU72Z54rfHQjpRJkMw0UtM0Nij0A2Jchwy66TUZvRfNUyRlOIRJPRkkcEj7wM+NZEkakangebBf+bw0e4Va4udgSNSCtPSD05XiXdM1Jo7sR8ls6PX8IBTSVYhtUPO8FpI9KddtDMat8kbcpoFBA9ERlxpkgZCS74ffv0hPxDARJBfP3w9qNNEH9LnQ+QaFLmNwScL4NbNeGO5pkLnN0MOHVcgYiXEhWS9/9sQLPh8HPI2eGBfiYEf01EBjJTkF6Q6ynoKysQGJsbydPHnc9g4Nqvk49mbc3oxPCDnL4JLkCX1fKgQQRULscr+C5Bga0JIlq1alL9zQ1KR10tbWYV9fvWJT0zNBigWjYRDdKdG02a8UvlwbwyPQh86kAqHvLrGgwyLLib0if5gMaBUvAll3FHb8am5sVpyOHj+slVx9VsMZniEm0TSFFhaWraOr29E4FRD4xDQSOKdo0wQ7cuSYPXj4SDrVHgtddozBDMke1xebAS5dBsrRfVVYC5LSYFiEXIXk8DwmeFxypDYxkljJOowao4ofgWmh80Z+RAwHfCAYi1OPH26g6FIOVaEVSeZJXEFeEyNkAhx8WOIgmaRRZu7pjF4fJh0NsrXVZRVmSeR3qiZPARpsdbU0VNHTBiFm1tzSakuLy5YvMtTIGPLkPHsKan5xj2guga4mseTZQiu/ffuezNM5mzwWRxkvzhH015vdXBct7SBrIlRsMJNkHfCsxGzDABe/Dnki1VlDrslWN9aFMJOMH8hIhouJGiHghXKGaSEUt+t7c89lSom8jBqhBevu7BBqmeeJ7AVnSE9vt01PTzgQABRUlkK1zg4OD0s/ntcE3U6DFi1/jGyRjQSxGan3rEueu87zSsUbPuzX1VXt3wuXLlpDa7PYHaC8GBgw3AT9hTY3bAr2HEUVjW3en7OFe7C2viLj2JpE1Zrqsnbs4AF78QSjw/ft8eMHdvv2M/v1bz7Q/aBhtmVJW9ss2NzCiq0XSpatb7CRF2PW1dlucwvoHddL1537JZnLyDjJZpQXrawua1BCEbWRL0hD/uXrV5J4G9h70J6OPNc+T4Ls1JTb/Z8Y3kiakOvAKFsBuWxnTp+ym7du6QxiX/Ts6tU57khDp78TN1lraGNL9iaY9cn4EEkgyWpwTheDaajHCRVfSAVW3FSeuMRZzq+oE068BXXJ2tIl0TSF5aSms7NLkqm0N+honIpl5nrCSCLp3PiRbxH3jyIN3V7lF8jM0QDidYlVNMWQ4AvyHy5D4zq9/I+fh1HDvSdGcD7h04F3i3TqJZkJ4ixhJQwVQ06yUzQHQ3k2a0Q/O8jGz8HIcgBcobMcTzTuoeICLJGqXbp4webnZ6Uv39yMFEJVqMiOji6bmZnTZ1tZWwkG3qZr7exisLWsuEwuAShF8a7qKDrOSvYD1wJKn+a2wDphUBH3pEwYNzbdByhI+ikfqXJv6tRQd2NRNzcVYGV11Trb2wPABfmgBvflCmc68Z+zg79nb0e0nc4aDRm5LxVJ4G1zTpBpwapAkkwNSqRVtm1zc9XOv39KQ0EkhQAz4RVDA6W2vkGDffLShhznTtGsWrL52Wl5SFArNDY3WNeuHvvzX76yxaUNq29okV/F4NA+m52fFSCB4Rifra2t01nP2ZzueRzYIJPC/WvvaBOAivifTjEsrdrbyamALA3GskFLnzVFUHc5Soa9zsJhMOgsAs9nydN13zRgcp36c+fOyST96ZOnGuq1NjUodsK6ZF/ArhGbgDy6VLBMTcJOnThq9VmkL1L2+uULO3v6lNCx7IuGXKPVZDL25dfX7MCho/bg8RM1NckByU25TtgnnBU+gMpZJlFjz588s57uVnlUTE2M6hzBfHt+fklDcmc0UCsgmePAEj4Y+WFdlvpiQw1l1pHOA5o86+vO6CsVrbenN8iQeqxBc50z5+jRIwIvAE67c/eenh+SIbwfZyBgJv7ddeVd9kIeezB4kKdjWE2uiBxeMmW7urpscnxSZ2xDY87RqMmE5alXkO8puDE7z4AcHkYa0m/IgJK/85k0rBAYwdev11xueOoo1NC8CYhenbXKiR1EJ5E9Mbu8vvBY6br3ah7luQaXKcE7jXvIXlOTts4bwcQwXo8zG78OYlthc0PyaLTJW5sb7fjRI3b3zj1JgAGAoJb+9Fe/sP/1f/nf7NPPLsvcenxi2T755Ly9efNGa+7UqVN29eo1O3jwgJ0+e1Zx48XTJ5KYSSTrbGMTQE7F1vPLdumD962hoc6ufP2tTU2tigFoxNxqUVKpQj9bjQ0N7tF9Gh97o1jF+j167Li9ePlKA2XuzfY2OTxx3+vG2HyMkssuPdhmp0+d2mEnkB+98xf0ut6fP01L91HTeZ9DHpOaOa0mqcsGIx/DPW8MYEU3r2UI5vWiSwTLPy/4U5Dzczaxznhf9gf3nTqcvaq9m3ZfMsCAPBt6BmIAlhwIw+BVOU7V/fNYY7xPjKmsA4a9nPWxNxHPSs6elsYGxb9CGe+4vH3y0XlLbm5YFf+bjjYbnZiwE+fOWLax2dJVZ7KvLMzIu+Tho6d26fJH9pcvvhII5KOPLtmuvh7tj4bWThsdeWEP7j+SPN3Zyx9YYT1vt+88sHuPXkpiDpYCwAoB12ozuheSphaDnWaoy8hIniaw+ThDuS/d3Z2638hUChAnJmJEjbtEKmc+uRZroATIR9I/znKsbiN7435HAjagpgALPtfgUuEyTi6ohxGNzqmf3KfJJR75ntgcjpJ93Hv2Eaj5sYlJ9VZUg/9oSBHrSWdapbw5DJCNeF3M61krJ9CBta114cMJABI+xKZepTbjHiEpTa1J7stKJx+CNZVGibi0ad2tjVZTLdpAX6ctTk1Y365uqYqcOv2e3fj+rg3t3W0jT57Zpcsf2MuRZwLzXPnqhp0+fcgeP5m04cODtrS8aHUNNKuL6h3V1dbZyuKyDQ3tsxu3ntmJ04fsm29v2JHTp+3tworde/zcci1tVk3WygMPKcmlhXmdA5ub69pHu3p63KNQAAxXxdAgST5bDCrwlSvZzJyflweGD9q9+/dtaGjIpudmd2p5JCvdo2JUeU0ElXGfGfRrbzoeakfRI4IbAHrFvFg5Vtif7D/J7LE3UzXeB0TdRLWjy8bzFZkSPKsoz+dAl0Yxiel5sYZQC6HG49mQ9/M+rMcokUQRSkyl5o/sYWICZxvvq+efrg2ShN7gj70QPi/7Ql4pwXNDfcKES7izZumniDkS8m9+57qoPcghGPgAjGDAILCmvHBcnpYBEvcmAvTisIOf5/46e8WH58RVaj+GIwzSeG48B4FHA/A69mxcsSD2V9Sp25Epj98T+1fqnQDG+WlQ8dfQmv/pM/z4DuxOOwpajZTQ3O1s75CZDH/f1tqmJgobCjNtNheonFj8wBogmaMII5iBktZGD/QlSXDU1drEJAZwbgIaaVFhB0o7k8k7wYvEkUNm8u3bnUlmbBirCA6TeS/kvNkd9S5JXjSUCDIzJLZ8BppCKvIogtGoDMaKoKtI3DFFJcmLpje8n5gcXE8OSvm2ra5tBJNZp6jyc0LNqVnnnxn0cWy0q5GfdvMjknXpsZc9qPE9Mu6hWNyqqgjj+6J+u4YhFE2JhFCLIC3F8EhzwLtUAAhLb965PmNEwLuHRHQe8CftB4QPPiKzgaBKA5fGxztDS9CSzliITXc+m2R2RLXzZrhTZB29zWeQVp8oaRQv4f6HIRSHmAdhD7gRfaxmCI3MVMLqsxh5eqJMoSc6/I+M8eL7a6KOth9NexkRe+GiyxW40QdWMjcNJpQJDM23XCaAAz+fd9YOmugxGdZg4UeNWMepBLrtjoGUy1d5seMDlYhY1IBI8lcBTatBAVqnGZk5ozu7f++g5eprbfLNGzXr0SLFlDdRk5ZO7SZ0zto6NYiVOEoyZUuyLQxJ8FwoFfM6bEnshYYs4tkARZkCMejWMzjA2JtikESRJEfoXBCZ7mPAfQIV5Q3mtPaeDNfFjKmqMU/jkEJNfhYBKeoDNrTP0ZWOhaozpCIaSfqL6bQaCpKMy6MH62tG5lbBf4F7xftynzRsCs3v2OTWMI7mfmFjZ5/xnjRupFdZKkomDkovcUdsEWRaSAaQeKqlsV9VI9s9dEqaBWBOCVHqxPFjashixPnq9YRVQKUz+AFhY3hBuEY0P6N1glaq5INAYvp6RhYEOi1FM9fU2tJm17/7TqbajgAxScKg4y+3GwnTO4qZRjGNXGIRTVzeyJEbNIazkocRiom1Fc2zkf5gINrSbD19fVoLIFBVYFLk0RhImLW3uFQdQ4qaVK3tGdovBJMPdGlsgggh+aeR1Sj2x4WLl+xf/vf/U2uL4jLqvTuS3/e6ZHCCdATv6TILAdUUJFXiXlfT5EdfcYgsHfBgchglWGgA8ffsafTpuY9i1hVd31hUfsnGcE/9/diyrCvyStY6z6fMkEJr2tHPQsTJY8kH6YqnTU2652grs7ZcFhDjz6Q8iRg+tzbnJLOwse7PsbmlTY0zGjU0dGjS8l7sk2TKG128f19vn70afeUDts28TAaFUtOAyeOGZGBgDW0g75TQHgCOyfXR9ONWg2Ik/vFpWb80lAE8pbNJa2lrs/7+QavN5KQxv7qxYTPT02oO43OBgTr65ho80wwKmtpRoot9CjLLkdc1iqG7+/pU1DUpLs7Z6fdP2fLSnIaEAwODYkXRqDp+8oTt2TPo+tCKpQV79PCBNNDRrmcvx8ScZyxN3UTi/2PvvbrjvM49z6cKoQqFnDNAAMw5UxItKln2sX3CnDkzfdvTN/OxZvVl30zP9Bmf9nGSlSmSIsUkZhA550Khcpj1+z/7peRZ/QXGS/DSIk2Char97v3sJ/yDnTt/Xs3nns4O29nalknpXmbfki0prYOQ9A0NQrhRRFGQc3YxYIX15IUnBu+OWkdjuaO1VegzKPsXTp2wb29+be///H3b2Viz3/33T+zKW6esGfNyzF0TTbaTPrBcqSoEL/Jdre0duquefP9E+0jSk01NMtmGer+1gccOz77dVpaWxaoifqXRMM+VLNWK7E3KmlLt9v3TZzI0JU9iTwhlqqqDeIN2L4anPvCHQVgq5hVHfUjoTBp5/QR9bwEWWlqlUaw7Pxi9Rs0TaYJLkoqf5XGYQgrPAr5ghsGqihoYkVwgd6To7fj3oI2eBs3WFPIyGtc+lBc7FIR2qSSDTGIXxTG6yzSCItRj1NQh3vO6/H8aF+wpsQHCUJs/B4UdNRVpetAYch1wz10ocslzNITVYAOUOQU7hZyj3ymJaUiIAStwhRdtym1+ZARJjJIhp2SjaOC6dItiVfDOkVRJLC4fLlg3U5MTGoAxSLtyiUHSPauUKgKfJJPNiosUo4tLC8o1Iq8pGtqYzXuu58adOv/cOxqAsV994MU+d0ShDyuiAb83zZzRqMG2Jx9vzBx57rx3Gi0aIhe9mc3Z5j6PWG5R1scZ9MLbmZ1uXMr9jq2Lx0H+HOkvDVkCUrFQcKCGon2N4Sqs4pidPnncOlqahRoH8Y03D03OlfUNsUd5DtwntUrRWpoT1tPVYdmDtBr7PX3d8h159uq1zcwsWXtHr5rrIOrFrqyV9d44i5wD7vK9XZc203MPjFbyIJ4h+Tifh0EFUiewO1hnwDPkqA4mcSNcMe503/jQirubZgh7wtnGLvfCPiWPiLSh8c9BipNn/OrVSzFJujoxocdvptH29tNqrCu3SNSblQt26fxZDXIACpDDSv6pt0+DRskPNaXsiy+/saMnTtv3z15YCc8g5HLb2u3gIK3BHAAP4jMSbbB9Xr94aQN9HfbW1QvWWIf/jDdzVlc3JKmTTh/Yq9cLwSOvZqPj45ISIhYjTcaQBWT1zvaO9gP1yebmtmIHMhUutUnzxtnI069ea0+Oj4/p87FvYcI3pVplpg3TGnANsl2Oos46sAC2tAYGMd2heHSwNuwkGoODfQNCJ/NMAQNkDvbFMDsA9MR+BCDHgB32GYOvnl4N4hgcUBMptxGAyEFYkVeQ2LMBvOGALDedj9gFkWwGg4YfwF9er7lMjKn2lOZ4qaR4qGaXmKrIusLYLKkxNjw0ov1Dvcv5ZojLfcFwgpyrmDvQ+Th14pjd/faurS6uWiLRIITzjRvv2v/1X/+rffDRu3b3229teTltH3x4VV4j/Nxr16/b7377bzpvXT39du3aRcVRmor0+vIFGJ1F6x/qtvPnj9nc3Gubfb1opTKNvKTVwTCoqwrMQBwFkBMBqSSLCntZ8qoJNTFV88IyZZAeeSUJaOasCmcjOJMUBszkxIQGHpIjrpUl7XqQyUpGitdwuSkffpLA8MuRo4c1KCC3XFtfV1McoCOxB3CQN98iFhqx0CVuHTDm0tACHsnjzwEryuFCU1T5TGAcc59xt3DfyR9I9Qb3aiRl401Aobhh9YpZ7rm255Y0CmleuyRm9BVJUbGn8bvLFjOqHX7z8VtW3N22ZLUqNYAXswvW0ddljU1NdmTqsNWKMC/jtrqwaHv7B9bV2ydj6oODot24cdnzi60t6x8dt931bbtz5zs7ND5il9++Zns7e7a1s28Vq7davFHngv94NtxjrjDgQ2xp2Os+wH/Oay16FgCxOAuwMTWwrdVkao7fDM9enjmNCQOFr2dQLIvVxj3jyhIMG5LyEBN4UabCdZbQeasG705HwBOvo+dFHUjuFuX65CPOYnSZSgFmlAe77BbnFznOL7/+WufeoW7OIudLoMGAQhcQFjZ2c0prS46PEgjnlMEo74vXJO9Qsz0wMXhNvDO2Njc1xJBqEcCgfF7guThg0ErBWhMN1lRnNjbUadsrS3bk8CHbXN+Qz8T9+09sfGzAHt5/bu99cE2MqRMnT9rtm7ftzNlT9uTJrF24dFaeMgxGisV9eWD29fbIHH1s9JDd/vaxTR47ZJ98dtfOv3XeNvZy9t3j59YE6r8aU96JtOGrl881/DrYT2uPkndqQKs8x0GuDjbys+DAizrb2t5R/sn340E2jMn32ppiPKwZ6nFy+ZcvXjijIsifvelFcSZgSARJaJdWDhJ5KKAEmamoFhQQUsDUSMEB1qDvNeKrZxgek5VrSC7Q+zXkyCiGRDURe4jnT10klYRC0SXTg/8G9ZbyJ7GlPL8SUBkgipr/eJ8AZiTHrFecYx+QY8OsIJ9kn3P/0YsTSE5qEd4zgInobAhnT0RsCz6rZHkVh5ALdYl2Ygtf/BvOMbmFFCUS5DEuEy7wJ9Lv+/sC3YkVE4CjnLNIOYXa0Rm5zrj98bAiJIJ/NagQCFNANnX23gxAHFv706Dir5oOP/2fv50VgFHB5cUBgHpLkdfe2qpmG0mzLghQCYWCKOoUDAR9EjWhoDo7ldDTaOdAy5wqNP1JIgugjxsTQhlDN9ekXrqRriVHMsKf0TDvH+hXEGXSzmsRWChmOcwkm1HDKjKeFGURrUlYEZrsevNMwTSMG3mPboDszXVHqSZUMEqCRAmZMyq8ue1NVy5q0ViDLjpISYInnzVCEUToRwKXm9C65BRNHya1eFuwtiQCNJ/dyKvgWnQB3U6Dgc9OYP2BEobub871gmNIHviE3o2V3ZSZ15MpOAE7NAXVQA8IeX7/YySdLgqmz6CXqjWnAwP+DHp/ukS4mDz8hWTCkTYEdz4fewB2SISG5jm6Zh4FRBhOBftx6ScHvcMoySBwk/T4s6V5XLK4Vay91c3poomDaMcyxHNGgzMy/HIDieUS8e5/wBMlUWaPSfZBiU297ab3NJmnQSJ/BzE/3Jg71dQsto5CfZhke/LnwwYNP/R2vPSPpIkcleUMF12Wb4ysXasxajb5n/s5qhTzljtI29Ejk3bqxFHb3FiThuT2XtpqMaiyrdba2S30TAHGSIXhAsZxnqyzLKDQCgf7atWwNlvbWy7nFPNEhfMRGZeyb0Gaae34DEIhN6ghjUybhi1B35TXiIZ8kaSULnhpKjv6qayiwpETNG4ixIE0SNlTouZ7IzZCwTAs4v3zvmR+LRq+oxcj9g1rL8ZIzNSop0nN9yFnI/o3VHwNBrzhxbPBowVpGH4OKArpGCtxc7QbSUFjQ6CsSyLEWV4qdKBWoovbgPF0zU6eOGpj4yOW2c/ai5dzVmW9aCJKh9cRIWUavlG8osAJ+t/4AFA0YOBMw4O1Jabw6ze377g8m9C9DW6eTeGEaWy+KBYAzJis0MUMa5wqDQJViZrOuRfgNGiJNzwP7U1RlzEedOqyxzoa9WiE11khl7XDkxM2OjSkQcVKkLrZ3s9IWsHRiPh1gCz2YoQY1dvTLzmj3/3+T4ph6pYHTxnvmXkjNKrh/Dn7YIWBgobA0u50iRGhqdVMck1ivmjCR41L/r20PSVt4kbaMm4XC8SLVTktgIIBCS7/C/RFHbkp9obQcrQvebt1zh4AbQ2SuODNTA1JKfmCRBZavBRnvDd0lCPmW6WEiVyDmkMUoh0dLTY40G3F/IHWJZPOiXlBc5eY0tqCQTPGhUVplkPPp/FO8be2sebow9BM5Z5hX0h6RMw99yKJ9HRllhaPW1dPt/6OIaZQYiTGDMI1HIpbb1+/HT4+ZU2SRgQNt681g2pPcV4GcbmXttXFJd3jOiPFwht2I2vm5pOZYHbq+uJxhuaNjbpfKzLoi9k719+2agWj2aJNTE7a7MysGstHjh4VwlzNbM68EHUFu/nll/oemmCtzSmXwwoeU7ls3i5euqh4UiBO1Wq2s70tSRHkX3ifnHnuzLHxccUMGDBu5g6aicGoo7bYgLxeItlgy8tr1tfZbL0dbfbO5cv2xSd/thvvXRe6+eubX6lw4YzSKAI1WtfYZDPzS5bVEIdGOB4dyCVkXBIOqTKa6bpzfZjAetFUYM1AEfLed3fTNjw8ImlA8gWLNdqDR4/VpCjVXOaHshImFuwDecWo2nevGWn5a1DBfsW8nCEmngBFFTNuHO0+BJwjBspQPinKuD8BF/B9kfQdz1USCaFwkrRfQ72Q6vhvdbZ3BBN1Z6lR1Ln+dr1kG4jBsP7YA+6R4xJl7HOaF/v7B2INYILLPkM6BIAHX5xBFXj8mmyywcFBxTb2PyhWGhvcL8RmZ8q5vKJkG4ImucyTGVIipZMAiVnWMJeDjYTMzi7G0zSfPSaQi8qzSVR6vyPdI8sbGxqCqgB19i77hrWiIet7yOMWz7a1iRgA7d6lUvIFvBX2JZ3BHuX+YBjN99M0gBUDapJYNzY66oyLvj4Vq5xZ1op1lYRBaAATt/jiuXgbxqXxuGOi/IEimC8hGJElCu9bEgnyxfKBO8+PWP/XaEjkS918VnIgobAWoCfEY9d/9rVx2UVi8g9rRxSVGWade8IxZIOHVC4XzGplO3PypKWSCWtBXjRIiXZ2ddv61o5tEk/VRKpZNrNnvV0d1tneYnlk1yjwq2XJUCB9sZ+BsUCM3LLB4RH54rS0IzvB54/L744hJvESuSHqDO1ZfE5irru/n0krByPfIzdhUMEdrJgTdJx5/tyhESiKLA4pow8+uGHPnj1TDOHs8e/Ij9h/MBBgK3sDrd72kTzr6FTDSAzF+jrdlTDJVBuJnbBv7c1Ji1fLdvXyBQ1OGfYCKKHZhM8FA1VYMvg8fH3zth0+ccqev3wtVh4yeQd5EOHUXTExRhhwI83HGVicm7Gezla7fOG0HTt6yIr5nGQq5+YWFdO4A168XLJUMwzGqh07fkK5HjJ+SJPMzLzWM0BqJWoUMdxS3hyPa2gPMpk8Q5Kj2ZxiD+yhdDqjs6a4XarKqBVJzvrGpNgEDgZyRDN7mmYv9VoKqcVyydrxYoLJilE7gLB0RjGe2M6wkzw+T5ypmobH5LyA3PiZU4cmnbUPOEdyhfj+OGtdCFuxZT1O47HAPo8Y1DRH8VGgae7SPwxnQfe7PEhkME1Tm1jEsIEaqA5D2q0t7RsG/eTuxA1JgMZMgyt+BfUcNVtdLgp0f4O1NCUsu5+2a1cv2fbGur18OS1wAyCADz+4Yf/lv/yf9uFH1+32rW9tczNj771/zV6+eC3pkctXr9pnf/lEOQ6SZ1evXbCOzna7c+tbq9WQeYTRytA8ZX/3mw9saWHONjd2LZnssEqtwcpx1pCcpyrQBmcBJgfxL72bVg3KfQI6G3lF7ljVcngPUeOIBOg69OQEzpTxeowzx6Di/r3vgn9F0Q5PHVY+gL+BUNSA2RhGAy4KzNrjx4+qnqU+4BwwrJC2vWKhD0+c2e0/6gewkksx8Ty5vyM5vYjNK9lfmLENLmunwbjyYG+NEtu8Bsq7HKoMvh0ASW5VDN4rb8A9X70JAAAgAElEQVRz9DhKLrsc+SZGw0t+NsMVGD7UDunsrurXf/77tyy/sWZdsGWLJVvf3rbBiXHVnGPDI5be2hZbm9yipbdPzVr2z/37j2xkqM9Gh4fFoujtHxDr+auvv9Wg4qOff6D8Ynlty8q1uGWLDHNLkpvjXvQ7j8Zqwb2PaFTTH0H6BrlexUCz4eEhrQ9eSxHLkXoCydeNzS0NZRkEsqHp45RLznakHyKvqFSzD4/rQcq7dDfMGuo0VtlZeT5QYt/wXpQ/4pESTH4dGODKENRp7D96Oc6adqYh3iqJZLN9/uWXQqpzrgBpUZdGPQNnVvu+UW2OCkMq+UYSkNrPUenuLcg9x71Jg5rzi69OAomeYLytfgcD1ErZRkdHlV838TmRIGyos972BttdX7GTx46ouU8cffDgoQ0M9NmDu0/tZ+9etgcPHtj58+fs9q17dvHiGZudW7ILly/Z7Vt3rLuvx1aXF1U7D/QMKRYyEHnw6KmNH5myP31y085cOW9Lm3v24OmMdfX1mtU32tZu2oaGB21xYd76e7ttb3dXd9Pg0FCQZgvgl+DRwx6ljyEQWzym58qfDY0M2/Pnz21kbEy5GsMDB7buyjD91atXjvpHEUAsNGSZvMHuBtg+0OTXqEcVMSsYRvv59eGhwJ3q0zjbXc+YXCMYYMsfK8QT7nhirYADoceiGpL+XQBnqN6Xogq9A7zOQn9B3hbOhozAxP5zHRzrvT9AKJF8kw84YS2Q1wvwSQ4YZKB4DWpt38MAyZz5q7oUScBg1O35g/8c9iPvDdAbP5OYBojKGWWe0/H9nCc+jwZoSZdm5yyRx9DbjL7oYbKu5JLEsEg9xb1JPavl68e5nvLHMOD1GjkEz7CO0RDjJ0bFm2X+6Td/Kysw0dyqoKiiSeh8GqxtnozLDNFNUilKe3p6dMlsbLieMn9Okx2qpSjpzc22vbWtQys0K9rpNAcTCYO+HR14TQ0jI2wZG6aUEEFJ5ZKiYUAgpMkJ3YoGpAJyoE5J6gI6fSql4h19XL64LKPCP7qwkJkg6QcRRyFCMo4nxs4eCI82XfJCEhAUGWRICx06ZJOBiyeAEOyReiIID/T3SV+ZxgJDGwILE+GoqSxZISb3QapE2vMkVvXuXeCFpu8emRIrMWhSsOKSjwzBCWAYvEUGRARKkpFI+5h/D4I6QqFwURCIGcpQdFDIsQYKaGEKqyaK6NneyEIHV8OJwHgg0GpYE5qiQq+E73XJLZ5Vs15Pz1YNFDf3icVqQlxpgg6aN4TRKMFkbSmMaEzSKNHnF0K/Xsk+F5q8OsrhNcKEGHq+I5H90gA1hGEVDRLWg6SDNdLAhkZysWzZfMHlUoI0Va6QU6KHNMvo6LhtbmxJmojP6wmVI3wcue5JIZ/bkX4uHSHEBk1FmBJJvCZclsdRON7Y9Sl/gyNK8zkhikHQokna19NpVy+fE6uC/TwzO2+vp5esuT1lyZY2a2rtMDDUhVLFEiQg4TJXkkYzEb3GOpPnCn9HkxXEJEUfZ0vPvujSSKzz6Nio1qWjvV3FGagwzhZrrwZlQJzwvrnI1VyWga1LVOgsvBnkuAm0Gt1hkBXJVgj9Lz1TR0BRGGiIE4u59024vDW844zF40r+ZURPUlNf54NIsSQ8oRXVl/0V9BlpuhF32LegRDgDLudWsxPHjinhTDQ12YP739ni/KzQnRjldnf1hL3pDSKkPkC9oV0/2N9jg4O9tr2dttm5Zen8HhTzSvqEtkDTv+ADF/kosLcio3nR5k3FIE0VybCQECebhPKkuUbBAaKUJJpmHfrH7GE+017wiYHyyp9Ln1OyUr7GQgoJqVZUk3d1dU1yG960rCnxZ6iLbjAJEZr9MDBAkF++cM5yoEgaEpZqa7cHT57ZLjEHDfnNTQ27ZCDb1KjGCH4KGMHdvXvftrZ3fTBAQRGGoZFHhht8OeOG2K5YIak6NPPRac8K8RlJ1am5J58Yb9TRxKBBpGS46ugTR5E4CpbXJ56ia0zMJl6yXvJriddpv/Mail94JSUbg2knXhN7ev7odbPH0hmG5f66NB5oOsIaUwMx6F7TqOMcshcpCJBLADnX1pyy8bFBK5UONPRKNBKbSxrAR2a/kvIDAVgzNRUx2YaNE52hehXr3twSUymSYAtmctw5FJjs/cj/pgwiqKlRhr0M1Q52dy2pZmqTHRobsytvX7G1zXVLY0qYRm+7Tt4nPCdQoYP9g7a6uGw7m5u2sris+4TCk8KlvrHB5mZm/R5naE9jGCYPOu5BYxUk3IVz58KQqCJNXs5RS3ePVfI5a5D0UsWeP3mhBjcNo7GxcYEXbt+5Y/Nz814YyVSSRiDSIS4bAEK4q7tLMdPPeML20alupNl3EJr2eBABRnBfBeIQuQMFNGdhbn7Jm/wUPEhRJRqshWKjVLCP37th3379lb119ZK8V2L1dZbLZnS3Yyap5iLIxr4BS6ZaLZPNi4nCs4kGszCc+DP2B/ukp7tTOsOwl4iPFG4pzL1bkIYq6XxLHiXZYs9evLL9bMaSLc0uJRbDh6ZJzfsIwY5xMDIOsJkwcWQNkbTii9hGk5acKmJGAPygmJGsmUyBobU32Mb6utYSlguoepoyAioEZKWYeBqjeJygcSR0WvCVEXItQVN2X/sVqS0+k0wO8Y2RBIo35o4ePSaJGYovDIsZfPDvKNCIaZGUCvlTb3eXnTp1yra3NiXnNTM7Y10dHW6qSZ4SkHY8OzwpuDvFEq1PKDdjIMtekMm8UJ5FxaetLdDgbgQMqljG30xsZbrqCMPIrJv7Tii7N0AC1xVmaCADRekQB+kXADKSnCP2lOzkqRMybSeOXbp43h49eqRCtz6OjGTFGuoabXNn08glKMBpvvOMWFtem/cF+4PX532JkScdfAdzeP4SFcyYG3uD3ocaoEA97yTDEEM1VKTEB/ZZb0+P7vP1jXXr6ep2nWpyqVLBmgEyFPLab/x8DWiCdKVkWUIjQCxhNQbclJOfJlCR5Pncc0AWzmL8MlRjgJa1q5euCiUfU8PYPc1A+Xb29Nji8oo3yUp5MQoaGfS2pmxjfVUeaPsM+dpabG1ty/azSILJYVUsi530nm1urysHlpRVT5/Nzc3r74ifXZ0Mbx2otLW9aUeOHNZQqKe7WwwKYglIbRprSPWwh4mFsMIEyKjDRBdJWc5Xu+oDZOVAeXNv7e/u28TEpJDh5N1oukfAFTEFkBTJHmgfM3zgLmS4yhkn7jI8Gh7oE2NhuL/bRof6rSnZaMtLyBxVbWpyXDka556c7uY339r44aP25Dm+PpwL6gRyvpzqjYHBAXs9PS3poVI+b5n0jnW0NtnF8yfs9KmjykWmnz23hcVleV7wGi9ezmC6o4a9/J2sZqOjY2pUslY0m9X0xegUgIokKyu+Z8M9LpAKg3gAajucxXYNoYlxsALzxYrNzMwor6/WGFywv7zRLA88kNc6y26qzR2QzexbW0ur6sLWljZbX13Xvzl86JBt7WxZoVyyjZ1dizfCmoXJDRuU+zYp1gzxgf+qjHmqRXlfkAcA0CJPYbAk6R41bxzIFMlqsPeRp4oazu5hcqBchKGz1x6eR8CYYqjBOca/R5kig5B6mF0MCuO6kyODZfLoIbFZi2q2JhMw4ci9Gm19dcN+80+/sImRYSscZOzrr2+p3nzv3Xftv/3r/2PvvveO3fzqW9vfz9qNG2/Z06cvxXw7dfKk/fGPf7SOzja9t+Mnjiouf/7Zl5YrVC2TxRC31za3V+3Dn1+X5OHXX9223d2iaoYaQMIya+X+ZNR9Z06fUV0/83rG2b8tbXbx4kV7/OR7DZ6joabyHmqcAMKCre4gp5rqF4bPRw4ftlvf3BIYhiH76dOnZaTNAEyAHOSaAJJJxpKmXtFOnz4lUMl+9kB3BrGSLyHwybcCwI3hrvsheKxW408sMR84ED/JF2nORyxfZ3s4W4Ln4pKwrizA65A/sZ8j8CJ9AsmXSgGAHKT0ht3hMqP+fsjVvTb3WlLStKkma25qERAvk93W+/mXf7xuBytLNtDWZoVs3mYWF+3Y2dO2m9nVkHt9bt6GkIpkYNTfb8lUs9U3tyjv3lxeVn/lL3/+xoZHhiXd9ZfPvrbB/i771d/9UjKtX9+6a0vrW5KHy5cYyjM29qak+9A5il3gCVjWsBGCrABrcHhyUmu+urZiH//85zYyMiJ/n2xm13r6+1QXb61tCADZ3tYR5NBoUONzCbuCvCOjMwqDaG9n14dCeFnCUJQRMc1YH07gMaZ7p1xyT4ggl8u9J7nf/Yz3SOR/4MMK6nQBXUoVu/Ptt7a4tCSWF2eVHlKk6sCd9KaJG5rSqsHDIJreEzkc+a5yT3nu4LfqPgRVehyNDZaGKU6dhQ9QXb3u3EGkWgt562xNWX21aO1NjdaaNCse7NnQ0JitLi3YubMn7f79Z3bkyIi9fjltZy9dsIff3rPTZ07ZJ3+6Y1evnbDZ2SW7fO2KPX78yPoH+sRo6GhrtXiVPoGJuf/02YwdPnlEHhWnLl61xY09u/voubUSfxoTtp/NqW7H3wKWDl5Z7OkeVBficQ3+hfRXJgeA0L1aJNVVq9na+obq06nDhzVIQfppbm7OkFAnlnE/cte9mp52NRD5kPgwSQBY9leQGIpyDx/4wGbG/8yVGSIwp/YiUqfysPBhEveBK2gEkKUAPyWXdwxqCh53HeRITyDKwTl3DDLIQTlj+xlAYg4IlDwZTEiZr3sOE93T0b4XXEV9LGcCCqgFq51ejRhlGHEjGVyTF5tAB/G47aV3tDf5Ps5MJLP0Y+Al3xfJzHH/AJhDzYG9R7xyhoep/+mAPu+XKAbpVzcsZ59G/jqREgr7lv/UwwIQqjWO5LqDEklgzigyhWekOPdG+8nBxfx7/feT9JOex09ff0MrMIDBYmBPqNkbr5MEA4aXJBc0IjSxLhblpcBBo2igOUSwo+DigkEqhksNRIea28HwlSKIwIEJTWRwGBnKRAhbRwV6wkBA9CLWpXP4IgGlSUeCETXVOdCRJrOa4UHKwiWFXGYjCqpcYE4pdOQhlzuIUAI0+ojegAZF78mAUNqBhqaCTsyB6DKGqu7JPgVhFDR5/9FlLCPOeExIeFCIvD0a65hpk1REHgvSbIwYG0Ib+CBCaONgOqRmR0CreMP+B3SB0JM0WCmWg1SSLufIDE2BMiCVCeLINIl14Aa9QsJTmsqsxwt+Na5/JKXgKMAfKJvR0EAU68Co8AY/KNuSNyZCwBVKWhqabhQYNfy5ANWcFJW3Kj8Qf948+7xr+oWGZnQxgZ7Tn8eqVqg4eo5LDWSVhgZ5vBcoRHJqGkdmryDIUOGBCo9e7862My0wDY4GZz6oCHIIgaLoqDOnmUfan0LaBu1tSRip+ePPBFM6lxxzSSi0nFPs2dyBQUbnv/HRQevr7bKJ8VHbWNuwFy+nhfDdTmct1dZpXf1D8jMAbafiSw37vLOOygXLZtKeyIdBUdQo4nPTRGXgxVBM0/+AchKKpeSa4W/Oi1AwbswUXY6iRAZ6o5t5+xArMt0SnTcg3p3m7Y0XhopOmXR6NckGDWBJ5AQZMRIS9xVwvUoSGgoP98RocOkMSXL4vojMo0kseA3OE5+N9zAyOqJ4IIMskOhdXXreDZKAK1m5BIIdKbWsra1veSKUozGflLQdOtqJ+pgN9vfaQH+PULFLKxtK/XNQyJEWg5WEyb3kWdijJjYDCZPo12EAqDMdr1cMxMcAtsfw6JhQj7dv31HB40wCb7Rz1mh88PkG+vuV1FBw0wxlqEFhQbIqRoZovi5PwICTYos3wmAOg1IQIQvzC3oGVABzs7N25cJ5G+ztEZ2ZImJ9J22ff3PLGltapU9LTKGRYJh3Jhutp69XTUPe950796yuIWFra5tB4gqUlLMO1Agl+QyU7CgG8zyj30eD6R/HIdYnYniRxImiG3nHBMYBe7unt9eRL9WSNEtBK7vET6OGNDSfvNhJqUBBOoJmSiSlRWJLMwizT4pghhYej9kHGb0Ga8yfIeEHSszjkSOZlYhWHT3f3JS05ibkDZett6dDA5P1tU29B8zoaDzNzM7Z6tq6GlkHebwJGiyZSmrIQ2MXVD4xRsNUUZndS8bl6Zyt5awsp6kzMCY2u3F2Tcg1vBeK+xkbHxqSnMjg8KDFE3XSo97YRTqOgS2G7XENKvGXyGey1pZqseXFJQ3jD5DRGOjXz3r58uWbgQDSEJxZDZKEQPO7Dao6DdDxQ6PSp08kGYpSUOR1lw2PjArVtLm1pdcmTkTSXOxpkn/JEbD2IBgDgohGM1/OAnJ93fnFJUnAsKl5Dmq65mE++nCQIaRk6mJxS2EQDcr6IKeih+fP/q1jaGY1e+vCOVt4PW1Hpg5JKx8ZPowok2qU5WxtfRO8la2sb1kbd8BexrZ2dnWGuF8jls5B7kDDCOn7B/kEMpm+vl5Ja3H6JO8kRLoJvNDd3W/bu2nb2NmSlJW8o3I5safwEJB8FU1pmJaS7ElpqO+tPfdL8OIa1ldNcj4MMGjAMkCgwcbAgmGkPAuaHEEYSTpwHzDI4Q4TCIOmWl3c1tfWBCwRipSmb3eXUIbUNngHMBTR0BHWF8yTwQENB0Cos9cP9g/E4mHgCzMENDV3CQwD1glZE0fkYZjZrM/53ns31KRliDjQh8/JijMTymXrHejXAJG9MX7okE2/mn4jh5TJZMX2w6eCe5p14NwMDQzYwuKSGJ3S2K64BxZB0RuRfn7VVHsjAfMDyiwq3DhwynmCbKPQgjTo3RhIr8PgtlUN/5zkHjC6ZY3wAeKOl09SstEWFucVD4nTrBN5BmeA98tzYX+y3kLncW+HtxMZS9LE8RzQC+7o7JETuTGss4KdLeeFJ8MuB4O4fKAzB1yGL94QlwRcBNxw1KkPfn0w6cMqvY6kVfwyg4WCvFZU8CLlRKxjrR18gReQr1CykYFbUYMKzNS9sRmTX0EM/yX0qHN4SzTIdPbY5ISVC97ATrWkJCezskIjBYRuUmj9FE3x9K4aaN5UhNnlYAWuGZiO/J6cxXNOU33BWVWDPci6ksfV875DLkM8uXTpgp4PJu98TrH8KiUNIoaHRzUwJy/f3U7bkSNH9HNev54OxqswNZyJ29oK0+tAEkptLSn9TJrCxHntwTia7QeSfTp1fMpmpjF+b5Af1vbmhu75/tAYZKhw5+4Dmzp2wp48f6U7oq7OG+cYaYOsZ++Q8yA/VibelAvW1pK0a1fPWU9Xq9hqM69e2ezsgo2NT1j/4LDNzC2pucmxIAdubW/X/orkNlRrADICSSxmpMtOKBcI0rHUeKurq9oj3BvkH7BF2fcMJbL5or189coaGYTFYC/CVmUNiFnIvtYkNyQJDHlBYcDbKNYo931/b5/NvkYmCDZzQvko0lc5Bly1mFVl7Mo+d988GuTsse098jdkEEt2/MiEzszrmTk1is6dOWszc/O2u5NWAxLGjPTH8XFirwpY5dLAAiShGa9BniNWHcUbk7QfawWzBYaMpJIYdHAvIiPC/gtySDD/iKfyEqprEJOXoYHVStbanLT0zo69+7MrYrYiJccdSG1N/vm7339mH3103b747LZizLvvvmPff/9cDfOpyUn75JM/S3qVJvDZc2est6/Hbn5z29LpgmULADtSVqxk7cOPfkab0r747KZlD6pWqtUpt4s1mNhLPD8abqdPntJzXJxfVD7HffPO9Z/ZrTu3nD0QzMQjD0DWR6jq0ORXniJwV78YFLdv3QqAsJpdvnTJ5mbnJJ8rH0EKLF3lNZenq1bs6NEpNUQBlTFUpzHMHcV6ZmCeSQWA+jQML6o03GGGO0Jc8jEBYKe6RZHemapiJsKosJgGoao1AkNPIEGQ0MGfCUatcizJmbocK/cLMYv4zvnEl43+RuRxx2uzv4kz1OgMUOl17O6vWX191f7572/YzuyMDXe2W61cs4XVVRuZHNcge2RwwHY3NqytGUBEznKVqvUMDlpnd7cz6XJ5y2Wy9uzJC+vs7rfdTNbu3//eRocH7Je/+ND20gf2p0+/trnFVavTEI8Y6x5PnF15CQaGAbkEsZGz7OUrl0TVxkZGNdCgYX79+tu2tLhsU1OH7PDEqO4J1dH19ba5sup3AWdQ9St3CoyxtMv7kRszgD/IBt8ZQAQw/l3aRixxhjFdnWJwy19AspUtku6mIcz6giYn/+TtnTxJY3/eFhbmLdGUsmtvXxejYn1tXT0eyRxKptplhdT01R5z1H4gRerz+h3ovqHUBZxHYif/ls/J/mOwzMQddpfMtIPYBjnt5KFJy+7vWVtzwhoqJetsTllLsmJ1laL19/Xb3s62jYwM2nf3XtmRo/028/K1Xb6CD9pTO33qhP35z7fsyuWT9vDhrF2/cUlDwKHBflteXraxkWHb284o32tqbrKnzxZs4uiofXnznl14+y17tbRmT1/OWUdPn2XlDcb91mLrq6vW09UpTw3uYwyhBegSINT96LgjJFuoJrgDgZdXVhXXyOMAYTKcmn49LXAm54ge0cjwiL148UJAxEjK202s3e9J51GMQmcX8LPosag3w7kOPboIAItMslQxlKfgN5P0nIO1DmwEAdASrp6hxrqGD+6lJLkkmDgCSgJUQg7ZexfEMAEjec6SR2fA6YoW7ofjTfsIZMo9Ly9b2KENSDEj++tDEvKx0CLU3Uc9JoZ5XZ16C01N9KdgJbq3I6/j4Dnv++nzBVklgWs07PKaidyP9Sd3FrAbecQfDUtcdtt9FaXWIuk2H4Q6owLpJwaNrrIS9SCjvDGSoos8hKKa24cUUa7r54IvXvOnQYWvxU9ff0MrMJZISUqGBA+ZApL0nuBRwd7X9Bkvg7bWNzptHG6SIA4FgYCiFFScTAH3M7o8ZXYWJDhIChhUREHCL9ofTGIkPxACmXTaSJhkqIxunqPmZDIT6ceFi1qazo2NjioU6jloWUYoiWC+rQazUENQ6Bl6+OSdxgpBAjM/op6a70FTvKuzQ40TmVc1uJQQFzSBhn8rXc4gNUVixmUZmTETbAjQyItwIZIEEBiJLTRb3uis0iCXfqNfFHyeN4k10+4KF67T4URTC3qAauYKTeJryBeXl0xOFUBBuTiyMLpUYMiABvQ/839LwsY3KxkIU2qQVwRFmX7H45bCNwEERJCp4GdEDTiX0wpeIfUeZLlMaLrxFb1fNbjD54vkCFSchn8/Mjyo5+2ae/6ZeV5qpmvQkXyjNwpCJ4ZGZTBxRvLkjWRCDs8GijQvTPh4XIAd3cjb9Gg/gtDk+dEI4+eLTSMaoTddnSVCEhyknwIjRc3zQC1W00G6oNGAA21X1jI0bl25QnIJoHsqxZwN9HTa8EC37e2ACGy3qfFxPS+aZzPza7a1d6CGcmOyxRKgB4LkGUUFSKa6OBrVQUoINDpeBsEbhmYTl6zWPDSfpP8cmhoRUoIL1LUT3cfE9dRdsitCmNH0j0zqo2GAN46Cpq1MTYPMFesWKPYkjIoTkm1wg2AoxjJGJU5QLImR4ftNnhE/Om9CZwX2AnGCBIkhIUUoDV3MBI8eOaLnNDu/IHmKyJxY7KxaVYjAnp5OOzRxSNrzIIcYXDU3t+rcI51AAt/T2W6JBjRXYXPkbTedkUdNHpmBUMzIdyMMbpWw0OSKKOpCwqMbTGHlnhJCVyearLu3W0hEUGuwLXjvfAYYNhHKAv+MocFB10tFFoJ9Yj48wluB/w/qyimwLoXD2lIo05R2ppsnW0KfQOMuV+zqxQvWgOmepE9qNreyYtMLSxZLJG03g+andgiHQjRwUJxjYxOS2ltYXA2MBxpdDW7ajBYqNNako62j989dEcWaSMc0QlQJyUpShzcRLJhQIIIAomFFPOTzse4MEoibLW2OvKThQdwkbrCWiaaktbd2qPiI9HBBP1KsaaiL54r0tf39iPpLM4Y9TBPfYmpWbWysuTdOI+eEJogbg/OrF8ExSSchmQXtulA4sJnp59bZ2epyfpiqJ5PW0dZhQ0PDuusYqOC7tJ3eExq0oalRzSLl0DHkbCohdjN8ILh4bJDkYYgbaoghaybplJhVYh6HJPFWqVpbMmljg4PW29Vp+VLeUm3Ntp/Pa1BheEsxhNXQzC1+auWKHaQz8qmQzm8spqYrcerh48e6x3w4LIqHD8yRzVI8K6jAjBpYNEMUE6Vx74ju9z/4wBaXljXck/FyFSP6ef38VAq/ELRYU2qYR8UAP5uiiiEQ/441YM3xPijSeFY8cVcgzpk3Ir2hwD6TP049A80gcRS8jmgq10p5a25ssEOgFzNp6+vusMHBPtva2bQaw4C6OjXzbt66bc1tnVYo16ypuc32MgcyHwQ92NfXI1aT0FTxOp1fhhIqgriPQVricxXADgJIJJIqUFiDkcExW1hesd1M2vIVGETOFKI5xWASVqTMgFtadJ4YOMAe5XNSpMgcW0VbxZsBMHFkzs6z9YKGPU++wR7X2eMuVrPW10xNWos5qj5Qyh1h3ug+P1n3+ZH0idh/7BlvMvC8dT+AzOWOlk6x330MBUCfkw9wTinCvOnLM/E7XrGo4A3lqakJ3Yt4nGEWSuxYWV4W+qw+0SiEpqOcKdAKOo+KFUG+RXI+0iSvV3OeITRNJIZHurMxjA8STz+WKVGeCOMr0ukN5rARA1CNypATeqHnnhZJ7k0xhuMaxHGIkGqYnJyQAanYrk3NGjrJZDzRaIvLC9oLNFT5uSBiGQrpvoAlCAgmMM2cDeYsxOhXH5g4SINfxagiZlNYK6cMDJGQvwgBH2Kb6y27t5cM2sUeMdve21FDkQaBo6FdHpTYACISphosCvJTH2qZJBVpDLnfVE1yXsX8D/JUSDnhT0FsqJHTkS/EavIckCRpHbJONcU8DfNjyPGYcpSTh6dsf2fbOrs7LFfMW1d3j0uOZGDr1Gu4ocGT9NRdX5qYyJrigwKKdMG2+9gAACAASURBVGVlTXElMvFk34wfGtP56e7ukX8LLB9v1LmRKrXD1NRhDb1gDzIwYw8BrGKf0mQmjqytrrukTLzeJg5NSM+bffD48WPb29tVrHv+6qW99dbbltlPy4dHz5omOJ5gAXiDXGOdVe3Q2KidP3tC9dPW1oatr2AMn7SmRrzx+AwtAqTc/e6RHT991r5/9lyD08Z6zjuSZ41W30gDCoPZNfeswu+FgWxj3D784B2rlLI2NNBvSwsLYoUcPXbC+gdHbGl5TQwDmA7sRcUC3b8OfILVQCxQ0xiGXxieqUarrxc7SmAHmhx19WrCM8hkTSU5GzMN94n7+BIxYAEQEOm8E5uQ5SIaOOs1Lt+GQvbAZcLizi7b2twRivrdGzf06+dffyVQTp74D0hG8nUxrWHEmtzbd48e6D4///Btm5yYsm+++UbsB86B2MGgeuT/ZdLgl9wnn58MXEAPzxP5EoI4kh0JdzFMLr5gg2PerQY9dWXQHY8AcZIqkrF2QvnG1sa28o9qpWSJhpjAL0hGffj+NXtw/7EVi1W7eO6wHT9xXDkaPgTDI4P2l798a5VS3q5fv2aPH7+UzCTDsj/98Q+h2VSzS5cvWG9fr335xdeWK5iYSAwq8oV9++jjdyVf+umnX9rBfkWDihh5fL036nxoWLArl6/Y7s62TU9P+wAnkbBf/OIX9qdPPpHJNfmjJFXx9ZKKADJJDjCMGmDkYpwFjIMfPnzojPNqzY4dO6bhNQAQ7oWI9SBZoOCZgyH7xua63g/Ibmd4uYyQS/U2vonX9BLcEN1jeGSOLgnUN4NZ95oRCDE06XgN1esi8XuzlO+RhAwstTCY0x2KPBbgKLGK6GkUbXLykNiC+D26Hw4DDr+fxE4PfYZ3f/auLS4u2dzia2tpjts///pd23j9yiYHBiQlhfTTyNQh29rdtjbABbs71tzUbJt4w7R12O5BxiYmp3QeBoaHLL22pRw72dIuMNU3t76z1paUffT+e5bJFuzPn35pi8vr1phqlcky5zpiAyKfHeWsklZtCH6IsI0FEAR9jsxMWiyof/j739jNm3dsZKTfjk6NKdc/f/68ckVACXxOvDPJlRjAcu4zB1kbGx232YV5S2cABcGMjNvz56+stblJaH1ympfTs9bW1mJnz5+1L7/Eg6Ngk1MTMgb/9NMvFPuuXLmsvfftt3d1Fn/1q1/b40ePNEQhzvzmH/7J/u9//VcBXdVz0GfwPfgmF1DfA7Y5ShrB8yDMZWAQ8Rk4n6DuBSJVHwXJsR1rxUQ9FlMc53GKyV2tSabx2JHDloP5xaAC366mhDU3Vqy5IWbtMK3NpXlfPl+w/sF2e/Xitb3z9lU1+0+eOG43b35rFy6esUePnts719+S1wZ7anZm3ibGh6yQZWjTplrk9cyS9Q332mdfPbJ3f37DHr2Yte+n57UfYLxTuwBWW1qct8GBftvbRpkkYT29fYqtyLB6vh7OECCj0DejwY+HED069jBsXVQGGCbCGCNOsu8HB4fs0aOH7m8R/D8iGW7Onvs14DPV7L6rIUY6OMKBDhFo1YuO0G8IwAGZX/N9kpp0sARfHlsAPbgCiPeoAMv+AKrl50niuFZ1jwqGwdTZQYbcpVB9cMDfC7QXALEec9xfh0GFmIViSQF+dDAmMYWBGzHF65XUG2AQ9Ya8XYOccTQ0ITeOgBKsgefSgEKcpRsNM1gzGPuRzwr/n7PJs9AgxZztFfmLqa+Wwq8H8CB3mHtueF8wAlh7X0+DiiBxFTEoXI3mB5+KKOfj+wVw+YlR4Yv309ffzgqMJpIKbPIMKPh0FAQhep1vKJCgcXM5XVgU1qsry7aXzlhTU6PQfxpQoMWWwCQUyQySEBrBNTUMKN6hY0cTVZIBJqlRIzsKEF7Q+VQ+orSpGJa2eoScc9ojzS5+nprygaYp3edK2eWjAhuDhhuar0pc0CuWGQ/GrQU1DwgqkXEPCRDsC4IFjSkSW0eIQEB2mpx3bzzwRYmPDJygLSfcQDYb9Hl13dK0oFHT0aEgDWKVQOXaxd6Yj9Bz6CVTBLIGBGMu1Pb2VmlkUhy7Z0bV0FrnUgEl5sajzggh4FGAOXUu4xp9BzkVEBo+ICkiRD7vzNciatQLbSf6GoZIbiwWeY1QAEvaJ1DqlGiGJFIJLxdMMAJ1OQYvztV0leGtU+FEQefyQb5Gfheg02M2MNgnqqa0mmuuMS0dWhoJ0nYmwUjqEhNaTGbnjnx36l9MVMFCzvVKRVnEID6g3Un6ee2V5RWXGwpoRlD3Qlcp2XVkuoqcN7JLXrQINR6aDawBa0NyT4NGzc9A7yOZ8nl5MJgCecvrF8vW0tRgJ49MWL1VbGV+wfq6m+zc+TOWATFT32T3Hj2z5fVtK1fjNjQy6okyBmbSMCdJ86aUsyMcaUKhHbFXWCeZ3Ql54zIq5HdCB0fIRBqBSGDwuqAXkS9AHkTJm683BRt6wKCCaSRLRkLNLX8tLm8xnUKTLPKJkRRHkC7jdX2I5bqXNC4HBwa092jIgIbljNLEZo90dXZJVoRi2hMMf77sj4Z4TcgI0Kv9AwO2vLKspI49RcMYzwcN8eQ/gfakI1H5exqCPHOhk9GjrlZ0Dv2c1etnsm5IwJXCQBQ5Gpc14WdAPogKQJcBc41vzBdB0GIA5gkUn4XYJ4kPpI0kY+N6zbw3DXJb8XMwGxzsd9RgrSaKMJJNsJEwimttR0rKNWLRdl5ZXbXHjx4rFp05c9aePH0ihApSMSCWWaeF2Xk7f+y4jQ8PiQmi4UFd3L66dcfqU612UCjJBJimQ0KGfDRPElaNVe3K5bfsk08/1yCoUmYdY2JwIIfEWsqAmxgJOimgSBjy9fS4pB6IUBJk5BpcZswl2vDPgWVAwaQGZLms9abJRDxvaW3zprWaXnF7Pf1aDVkKL9hI7HFQeNDbWWdktvzZOcIHeRlilQbGkoHhjNSLTcHwmfhEDEVKBFSjjPwwNKZYjcWVjHd1d1smva9zTJMIbe+Tx49qULAwP2OTk2NufgtyqFi01lSL7gUYLVwFNGCX19Zsdn7RCjABKIZLNJeb5DkjGbRSWXJuULAxSmTAJsSmBqEh5ogNVFSCzdkF9QWGbhQ0WkOdawPX11lXT4/NLS5bHahEGswEhXhMAwDOEfGAO4OBSjGbt0OHxoUGRALpwZNHrjcuL4CEGphDgwMaECG7poZmI2fOpchqVvah5hvvGZfAwIdCNGhiZ0DwSLot0WClQl6yLULBBl1/muvsG56j5LOam3WGVjc2WKA3VGf2McGfZwGyjDMmvVwNKzwGxc1je7aQU2O5lMtaQ6xmI329YlbEq0V5Ae2lt20vvWuxhgYbHsPI8J61dXbbQb5oL6bn7fTZc/b85SsVkT4chVrvpt4Mx2TCSePDYD71yRyVtaThd+bsOTE6QFk3NTVbqqlVjI39fFb3BkNP9ik+IendPUlAbGxuyEsEvW7k0Rjmcp46kfni3+ztihmouy4MtASIyHkxFPk1EceJu/19fUIwiu2ah43QrrjsQwtnC2kgqMYlvi6eT7kZqg/L+JVzJbnEKnKJeUnj+fAPFBmD5qximMAJ5AVxmC4Y5wLq8NdN72fs+MnjMnNkiNcoD50GNXAye/u2urLiPiANDdbd2xPeA2h+b5BF0i1Cx+5nbX/PvV7Yi+jBL62uqKFJM51mO/uDHE1otGxWa8qaRLrJKh4DKlhsQU/CHHEbmvjKJ0HVNjpTjHWZPDyh58swYGLCzz33Bp8FJDjnk5gyPz8roAsNcIpMGgJIngFqIfdQEyAMJ5xZjASX+7TxXFxKwXNKYgo5mvKQoE3MWpNrKQdtAmEYmgN1cTXp21rag9+GtxNpYES6yXyvBsQ/8uTgDJGj8GfeqAWI4RrOagLDhNVQFeYuZ8Elc5xtxoAqaQUQf2LmxjT0ak7BgoBVydCExoEPGzo7WuU5Njrcb11trba9u6uinuwJeTy8RpAxAURBSwEUPGbklSrgIW88d3X1CHFd4t4ln0iA0oRFx5DBQStiosVi7g1SrekskIOSl/T29ltPd5e+V2Ch5mbdp0jaiIEr1kbJ0nv7kjeDPR7ldJzN5eUlSbLMzc2KYcEzlrm7wBAxeRGx//jMSRmIl8QmOHZsynZ29pQz0JjP7afVcILVxFpv7+7ZvQePbXh83NbwrhFb0xs6Yo7Vx6y3p9ul7vCDo4G6tWHdHc329rULNnV4VDIlr54/Vwwm3z9/4aItLa9apcaNRd4RU8ORRjSyKvzanGxy6Y89NM+rtrq2qnua9WK/Y5ZMk+bp06fW29Orv588fFiNFCSxkAvBX4BBE/uEnJLnSayTb10+K8YysUYswkSDtaYSVm8la0k1Wktzk60ur1hnZ588NU6cPGO7exmbnacJmhEzL05OEtDrkhKV7GRzYK0XrSVRZ2dOHLWjRw7b4ydPJA8JEIS146yxZjBl8LMA1LC0suN5CHkY+5ocXHJd3hCK2NwM5jkDLm1ccgNvycc5+1vgLQBNyDI2NLqnYbGgfJE9gIQiIAj2PIMKGLj//E+/lPzoNzfvW6wWs4uXjqq5Sc5LrvD1l9/Y0uKevffeZXv+fNZ6ejvtyNHj9off/U6Dtc2NjL19/YIajJ99edMq1Xrb38tZa1ubZQ527Ve/+kAD1c8++8Y2t3PiC4hREC8rv2tINFjuIG8XLl6QDN/S4pIQ8zCSP/74Y/v3f/+9N3YD8yCSz9IQO9wRUTOUJhveBIcPH5Y8D7kruR+DCvbO/PyCYrU3I92TjHXntWGfCqHcUGdzC/NaPw3Fa7DSGY66PBP/IxfzM4hPY0HAiEgqj3PufhbILHvzWj4i3GlxR3QLca+hgtfaLmlGLgVYxmM37FCG60gVk6ecPHFMTWAM5F9OzwmswGDOPTaK8k1kKHvt2iXl4Qzen09/b7u7efvf/+Mv7emdWzYxMCCfnOWNDRs6NC6gExIvO8vLOnfzC8vW0z9gmVxWOceTRw9sdGRY9VDvADKULRZrarb0bsZevZi2VKLZEk0ttrK2JaZuqrXdpS6RoVaj0z+7GG7UcoERHAEOifUCE1Ud+MLQFA/R+/cf2/GTUzY8MmC//90n9r/8r/9o9TWzb2/fte+fPLdaLGaXrly1F69mAoO5w967ccP+9OlnqpV43jB1vrt/X3vnww/et7X1NXv+7Lk1Jprs4198ZH/8wx9UZyI7d/ToEftv//pvqjEuX7qsfXXn9m3dV//pf/tP9uUXX9qDh49sZGTIPv7lL+23//bfNfjiXMqrkIAiuRtvkEfIefUg3sjNOSiVc0pt6cMHPIZgMBM/mvTZ8Y+TBxagWUOFw8F+MECPHTlqB7s71t/dbtmdLRvq7bK6WlZDi97ufsn0AlYCLAG7lVoSE+2nT17ZyZMTdvOrB3bl2mmbnZuxK1cv2+ef37IjR4/Yw/tPbXS0yzCPaW5qVSybnp23gdF+u3f/hZ27+o49evHaphcWrA0ApWJTWUC09bVVeZiQN7GjYUZwHhgGa7CIxBag26r7KRCT8NKgtqapD/gWxjO1L3fYQP+A9hB328jIqPwr2N9C+QtE6OxNQDPeS+FedxaBVBRCrui1vPtWsO5iGQgc42Beahcxh4N0uA8EyWn52e6rRjyRpCnG0qqtHQwbsQyi/iDfI9YH8Yi+BDlpqCt5HXlyBna/d2J/YNES57irubcZRsjHpeLgokilhNjA95EvIfdH/qS9V0CylgGQ52rERs4Zf896eR7tfl7EFCQo99J7GrIJbBBYEg6s4z3XhZ5ATM9JYgZBPpmhGp+Bu0vvntYiAG3JWwH6dQbNG6pE8FDVcCaAiqWeEtRMoiGHBrY/DSr+dhr0P30SX4HxppSMjCIjKYqoocEhW1tdVbNSPgkBeU5hzICAIYZMmaVr2qImEoMMjCBp1kXmgPI1CCgJzGdUJEk+xiesBAo/owGN7vxRD5gB8S/uRZAj0u+lM0hw9YaKBhlBkibSpvNizxHKfBEQ+U7QRWqEtDpCj8YVTS1p6JEwBxkGijompBSt8mnAL6OAQTZDERIuBgKuQewTUEHOdAFqClwjoDuzQQE5TPhdQ9bRivwFAVlNWQpcGs2SePGkBISslwQxBXZ+pdAS2hwzu+YmoelAxtG4dP171tWLKrQnQZVRXAiBAboul5V3gzdcA0o8NOKFRgxSA5EMlwInFFjYNiok3HRI6LSgXRjJCQh5LR1+R7Y4qyQ0msQO8eSUgoY9xf6Rx0SsasODA0Fv2pGRbAP2BwkdF5OvO9rIThmOnq2jidHGLGstVWTrAnd9Ud4HlzPfR4ObdWOAg/4raHeMpSIEzw+MipqM/jSzlomrSTtXTY7IV6Xqxb+aCGj1k0hwmYLUrIBQoZkdD/JhJI4V66MgLJesqzVlHS2NVm8560d6h8ZD2awSb7TFlQ2rxRqk386+KjPcEbPINbmZ4pPoS86oWBYyjS9Hk3PhgybwZqzTOR1hI9+WsE4UDNFwJioy9LMCoyV6ZpFheoRS5ax5UeMoCqHQNThzqqia90E/nsXj35M8sW78HWueL/jQzJNRhlc+/IhkqpCbk5FsE/4qddaSarLGeM3yuaKdOHFMqD4athRevDYDVRJcnhYNEffXQL+f5+AGovxK04kzBvqLptHY2JhiG0kb7x29Z99jnF/O4g+sEiVlJAQkaZidVoKfR6WixsThw5P6rBRINItlVB9Mw/i38q8owAgpaohKMknx1t7SYrVy2c6dPm3NIFvRkq5W7OH3j6RBTaOOAQ7NYai819++roYW+1iNm/1MQHjkrJzP2wdvvWMNSv5KSqoXV1fs0bMXVmSt8iVLgpJBVqNMU77RWlqTas7V1yfs0aOnMrWDbeTaoD7E5Fmznq0tTTY4MOgm7PIHYWCVk+SfDNeCXr0QvYHFxdCBtSJucuZ4LZA/rIf7v5FweWwnfj188MCOHjsis1S+N4ppPlBF+9Sp3q5D77FBqBrph7rOOvtcBuTdXSogaVR8/+SJfs/3kpwWiiTksMEb7drVa3bv3j1HLMuPBx8T5BwonqEkF6VtvrXjVH7Rzw3WQFJrz4CG5sDKxrpNzy7Y+uaeWR0DWZqnoIGgDNOsJEZUFEeEtKH5QVMaeSOfe6uRocSUYqw+ZsVszs6cmLKD9K5ir+TeGN6UKra9tyuJH4zBaWCAJCKeIssjiZoG5M7ytrWxZVcvX7F8MW+La0gvOrNQ0kVK5t3cFPYO3i80JSXBFpgXnEMKERqTxFeQtewh5D982B4X8h3ENlS6Y0fdgFBst3CXyLdGsk4UjzClipKVTKLZHOTIukKzjJyjB0ZD0T1BADkhscHQiyFapRITk7O5rUX7hHODFvhAR4edPXnMFmen7dLFszY/99rSmbTYNafPX7BH3z+113OL1tXXb/NLazZ5+Ji9fDWtu5zNIM+GvR2Xh5P8RoOGiMR/Cr7nT5/KkwCwxekzpxWHOSd8lqGhUXv89JnQxisbeMZ4AcTQCKwjzXSKFJ4BZ4K4LEAB/kXBTE/7O6DD+LOIWSajQ7G1XMrQUcuOOuM/fwagoH04wsCKpqxQzOi8c8dyBnMHOnfsLdizNNnlVxM36+zstrYOtNFpCPnARiy+Opr4NA4o1gCcVK0xiScCeRJi0xXr6++zM+fOqQlIow80PJJJbaAIY3WWBYk9N69mNmeS+JlqTmrvinKfAnzAYL1i2UxOB6FaJt6DMsMInjsRCQwMcitWKlY1COEMuhQXqAbXDxZTAMCGBuiukawcMgBBJL1HjkTOyYBUd1Y8SH74EGdsfEyfPwLjEK/IP9wY2+9fYiTGmjQfiPu8V2csej7N3o2kFnjuxE+dqfp6AWKEQKb4lQSBfwZQ4GoIcB7UTHfJUxWs8mLDvJxBzr5724C+bEGmiu9Fpoyhv0uHkTtyf7GmahzCBAxM3GjPEN8l9xl+hqMc3etLyMpSWfvJBxYVNGWsVvP8jgEgMpOVEnkvuTisDMAf5CGwsppscnzI0rvb1t83oKE3TBNpaKsxUW+7+xmdK5C73OWxOryxktof/BngAPYTSF/eJwM/YhwSOQyFeG88c2I9d6v2Z8j3h4eGjHiiodABUmPkrw36Pfcnd6d0rJFy2d3Vr3x2nhlnBv89sY1gfKqJQlxGsqpBeYiaD1n8ihJqVKdSCffOKeINF1O+0dnebhCO+vt69Ay4M5dWV21je9cOCgVr6+yULExne5ct0qzqaFeTWob2NN8xkK1VbXtz1TrbUvbBe+9YW2uDBvgvnj4RG5FnfPXqO/LD+u7BIzvIFWzyyFH75tZda+/stJNnzij+i6XQgCyKszbv3Lljw4NDursiSU7yxZcvX9vo6LCtrm/Z0WOHQ6zYVg6ysbWls00sYB0AimSyWTXsqzXyUJfxZLAD6CKVqLN4NW+nT0zZmVNH7cWzF/bs2bQ1t3ZaocjaumErQ0bAG4AxCEbITe3suTQrAyX5INbXCeFczGXsl7/42La2t4XGZlDDHqK5x59pr4b7s1KL2bPn07ovYXFJhjDE4WgYTD7GejKoUWMLMEfwQlQ9GV4vqosjDXHyYFiDAPS4LzOZPauW8mL3kR38z//yG+vqaLHNtRU1gjvaW+3w4XFb39y2i1cuSuLm7rf3BCB49mzeBge7bHJyym5+fVMyVPz9tbeu6u764uYdi8XwtMurUZzL7tnHv3zfMtmM3bp13w4OQMInrC5Rbwf5vTeDGe5o/ChghS0uLOosEK+uv/Mz+/yzz5RHqTYOgDWhfYMJsn8+15RnE+C5QL5Mk5q/Q60RhgVnB7P7aADqgAKPEcTnY8ePq4dAnfrs2YvgbYbcCfeKI6nJyYnDAPvYz96gg3ENmM2RxVFdoTikWtzPruqiICEMYE+yUgkHWggAlUFm1HNG4nA8zlrhd5OxoYEeu3jutBULFeXapUrNpqdnFJvEyEg0WmdHmwaeSPlU1EeoWvpg23a2l+0ffvmBvXzwwCYHBmVWvr63YxPHjln6ICPgTekgaym8apZXLdXSqjvj3PlztjA3Z12d7Rr2b+/t2fChCUu0tFmtPmlzL2ctn0Wqps3K1TrJsGIyT+u4whlTjQc220FSAMoYrBCveZbke/zKc+zr6RLAsbu70148e6Y+QXdPhyWbU3b3zl37x9/8SrH5T7//xO7cfWRtHc3263/8R/vjJ5/a3u6+fEFh5Pz5k0/EqEDqi3jxpz9/oiHsjfdu2KuXr2TMDmji/Q/et9/+9reWyxdtbHRE/iS//8MfdaedOnVC8frhw0d6vvixLC37YJ89wCD32fPnQdKYz1YR4041qRD5rr0fNaN1p+by3kcJqH5qJaHtYw6mVL8mh1RlWT5X7BuaxzH8LemtIIW0f2BHDk1YmTqmpcnK2bSNDfVYKZe2toZ6a02hqJHVgIvnhzw1g/ETJ0/ZsyfPbfzQsH315UN5VLycfmU33n/bPvvLbTt67Ji9ePFMjIq9raKlkviI1dvM/KqNTQ3Ydw9e2akLb9mz13P2enHRUl3tlqWuFrut1dZX16yvxxmDxGx6bpLZkpSjN+xroKA0wGMY5ybVeHwAAqIOWttYt+HhYZt+9UpSycqnDzLqhcAwjxgVkUy3G03D4PWQwD0dsSioBYh9kQpIxCLg+5D1dk9UR/LT13H0P7WF50zUYJJjlx+oAyMliVmtBo8V8lOkMN0rh2cDaMYBqS4/zX/eL2BQ56yGyMPk/9vHhf1Jj5Iv9cIEmPRenACMYbgp9k3SPzd7y/sYPrSmZ6bPF5hXUuwIMqf8BbWaFAWCjxjPQKDZasiXqFlhtoW+QySxKuZpkKXjWbGmAJc9B/Yc0N+o52JRThl+zBtfHgFOgrqMM87cZF5Saez2nwYVP7X3/9ZWYCzZJBofDWi/EExmbhS/UQDh8qPQ5TAQPGkW0DTmIBFIO9s71AAnINHcF5tBiKs6Ff8khSS6EYLOqeLRxNBXNEJXOJosWEeFKaNkIcL01YtzLzIdHcj79n8v2ajwGWhIEigIogRUUEoUDSDaGFSo6Z5EimHHte1CUCTRYS24BCiGoyCLWSbB1Ol2oE3LKgzVxJRkggc6mcYifcOAIdWsNSSA8Jpcpq4niQeGN035Ofq7EshrUGveBMpnoU1jwtPqCJGw8XS5yI+QwFSW2R2JJQ0dNWj1npwOyWeLUHZcQdlCVgmOPhvUvvAlWYKgfxw1ZqP/T3HP56Zhgoar63N7Yei+HV5MRvr1NGNF0QxDCl6by0nsFBq4RTdyjsyZaQqOj48KAeoNz6B7+EZXNjI58mJSF2nF0TSSnQhapv7cfU9FKE0aqUKO7e1p8i2D7GRCEgOLi8vB+AhqnVP0CPqSSwo68nTS5RMgQqF/RZ9V0gXhcqkGpKZQh7rsAwOD/dKYsPzBgUx6J4YHrVrIWWE/Y5NjnY4gb0xarlix9a1d6c4XyzUhbfJCgbgWsgYLIDADdR05Dv5TMy3QFdV0CPqlaN27VrwnNOxJ9t6bjopruugruvC4iDVkC9JX/DzWJJJ+88aXF6Ts0chAW8V8QEXQ8IhMkiMkTMQwIIkUoo1EhCIXqmQ2L3RchCIA9ejGaZ7USPKqanbkyLgKUxpxQ6Ojet80dED80fCRkTSIX55Tvcus0SCkUUfhICmhZDI0p+qEpL979zsVH6xtS1v7X/ndREVU1OAh7kVDTz6Xn2mPiZJtCwwhPr9komRUjvGj0zvX19eD8WnJmtudAYL8ExJMoCg3aMbVx61QLor1JOpyvE7yR0jq0Ihh0AOKcHV51RvzdW52SYO0OZGwK2fPiHJdLual6X/n7j3bh1Zai1m26LqfYjYU89Lbbu9otatXLtvde9/JqLi+AXQNUjH4nBD/6uQxACaZoofPEqE2JMkDUkaDM5dKk070gdNihaaH/UOTgEH3G2+LKFl0CTKQKzRLQA+yD5CjIobRdIwYXDQw1eSTJl+FJgAAIABJREFUdBVSJkgLugm3zkSJgTO6qAV50NC4IMHl70F7UyC5Pwpnrd6KhYNQ6LpkCEyQuhhNu5p8TkCEtrWmbHiw39LpXatUira5vWktyZSG1zIdhg2EQV9mX+yKZvZyqSCE6KvpeUuns9IWlkktvdQGl7RRvCQBhVnGOYrRKMVI1OW1dPeBEpOPStyGejrt6NQhNVEPMlmZMm5u71kl9sMwlT1IEULzis/IwEz3HmskL5RBlzUrFjRIkycB8VzIYsxAk2p0MrjlTkXmhgEFTWIG2zRlKNAkLSMklsdxp+V5vEV6DPTe5MSETAs5X5LMgJmFiSaFoZ4fKC1HaeaQHdIwMyfjQBn8NrikGQ0fYhGsie7OLp0p0O1zC8tC5RPL6xvjaubhU9Hf3m6/+Oh9++aLT+3K5fO2tDTniNgY7LQxe/zkmS0sr9mhycP29MVrO3HqjD159lzsD/k5xWKW3tsN0o6grVw6olSs2NEjE2JUTE1NSu7r0qWLGhaqSSDkfr01NqW0R+YWl1wTGdRxpeb+TDRmYiYJHDwOuI8pYhRvg96uqOvSaXfghucLzpSkoRflQ2qWS0rOG9DEGeQTNtY33IhQOtvIZZS1xgwDOEvKM8LwHtSwTNSLLjHFWeLcuNSVe0YxzKqvI19qtGy2YA1C6MMYQS+7Zr39PTZ1ZEr/jjO4tbMtORRAH7y3ZGPSdja3bW15zbY3N9U0GBoZUa4IW0YSREkGLi5PQ+7C/t7c2Lbd7b0gheWgiK3dXWtMpuRzgVQXjS2mNgz7GAKytuQ0ovcHcIvLhcZBGOjzUeDr7gr3nrxZxL5jbZE9dMQx+59nj3QQMVveLMhOFXzQzffBakBWj++B2cobYF9IzqDqA3r2LutL7iakYwDmkPtE6MHIND26a6K7GARo1EwRm0bDTM9PNOT6kf+Fe7cxtCZ2+uBEuZx3IN98uY6z51wa3oQBhbMlPaeKUJR+Rh2coqEnZt8ynndPH+UEyvsYDjVJWlHa7hWYmej219n4yKB7c5HbSpuZRjDyWc58YW6CpxDMAA2COBsJvy/xfSEWcd7xdOM1WDdydJixxBpp/x/s673QzOYDcWaEAi3BJmV4QDOBxh3PwyUp2GvOAAHc48xpvoRUDcwTXoyhRqKpUbGe+oIBbVtbhxr1kY8Wa5FJ76m5j3zc61cvPX8kh+V81sp2eGpSuRFAIwZu61vblkS/XXrsKY9zcZe6JXdDzo4BEOw+GJfLC3PW0ZK0j3/+rhUL+zY8NGDPH39vC/OLdv7iRWvt7LHM7p7Nzi/Zzl7aunv77fXsomTWevv7fYjG2pQr2t9+P7jUlBi0SNruYkbu4CchlEOjxGsCmI+tYp4gfUNWK6xOvE7NX9iN+IERGyJptmRDoyXqzVKNMWtN1tnZMyek1w66nNy2u6tHvmuA48jLz5w7a/vZghDW8XpQ9WXb2U1bd0+vjY4eslevXtiJqXErFbIaELpkCXmt5+W8HfJJ5UfbO7awuGCjY8jwpCX5p2cuOQy8gEpCVUcyp9xloK75rHgVMnyOGGdRLP5hQOGebOwrgiXnpKOtXUMq+VRUi2IeffDeWwJfjY6OaLiCCfvmxobdufvS/u7X7yin8wF1wb74/KaYliPDw/I04yysr+/Ye++/I0bMnz//yuLxpGX2yVM43wf2wc/flQLC/QfPLJ0uW6FSE4uiWgv1o6QlaxpU4AOAXxo1K8/4rWvX7IsvvnSJucCsQ0KOeOMSfF4D+Rl3Mf/h4SEx2wCS6Kuuzo4dPSqWDWbdquODESxr14SqQalkJ0+fto31NYEAQXbzyKIhA+eafEiAuBAbCc2cXf6tOPJv2G80lqlTqDkdfBaxNniv7NvIk8eNph3UVirwrJzpr+ZiPQCiBiHtj02OWUreN2aLS6s2MjYuWSNAbvq3Jc9rASHhU8BnaqBWS5itbyzY+z+7auuvX9sg6PWNbVvd2rRj585YDvkoYkDOzxgyS82AN7N5O3IcIMWM55t1MYEaWju6LVsu26Ejx23mxayVSzVLpdrtKb+v1CyTy1mJO7LkMsi8P0n2svcByImt7YBApJyIgXydOn7MP0OQLmKo2tLWbAfZfd2D1y5fsY6uHvvz7/5o9+4/to6eTvvFr39tf/rL57azvaPhwckTp+zBg/vyq0Byjz+DQcE909nRKaAXfQ6eIaw02AbkE1F+GDWSyXnZu44c5950vzkBNQSqrMrPglzdcyAXApXEZGAA8pn82f/gFRDJfEWMNL438hThfDFEVHOf/lBYK84JuTaxA4DN4fFDtrW2bv2dLVbY37OJsUEr59PW3dxkTQ0w3hiA4We5b+3tzdrvJ0+dkqTW0NCg3fz6oV26fMwePX5hf/frG/bHP3xtx04cs+npF/LU2d7Yt/ZWpJeytr65a92DHXbv3iu79M4Ne/Dslc2vrlpHf4+knwBjSBp0a9v6kF7f3REYiprD2TTeMxNi3reBD7VDv4s17BSTsMGWVlbFeMfDcHx8XPUAdx6M15nZWQ1wGAiphxM8L7jzyCl5D2JFBEUEZ+kiNe7N80geXT+Xcw+7Pfi9ChAb3o8AUYH1yr1OvQ4rijVVvhD6Z/IHZOhCXBUYEvmxvPJcdXIiadswVHXZUPfA8K+/Zh3wOsQ7saIBT6p57x6rWi8Av8Wicgj6NeTG0WCD9+Z9RAd2ek8oyAMHhol6HKE+iHIHyRaHlMsBnSXd+YDHFM8qVQ2hI39RcghyCw3M1Ed1CVzvv/j+V3vGrzn/lGIyuqedZJTlD+vPxAcVLhslsPFPg4q/yn9/+j9/AyuA9JP7TTjqiwCILiUmiBRZBHwlcgcH1tPVrck6xmsUwVzqBFKhyzj8zc266CTJEZIOGkego6BUo9VKwJOGOLIYoeiKllHDCtF0g9yOJFwCuv1HJqxq5suUxhxtqsZd0JgLzVsmpZKgAYkQEPFcsFKxrKENB5MCOQNQjzklsGQ0EZpampDl0KgWot0sB3KtDlqp683xOiRXFMYU+Sp+E42ik/FaIBOgsdN8oShG71joyPBZuOzVuJC+pKkIA/0FWi6fzSmoUijI1yEEWgoYL7BBiMStf6Bfl4rT69zMM58taHIODZBiNkpAaTwVy0FnOhjWOb2Md+uBjuDJhSJaHxT70NBm6CIpkGBIqcZAkGtSwSvPEUf+s1+iolyyWWEwxYUgc0fQVAEhDXIFbXqkIoj2oukGqRj2pDRz29rUbKSoior4KEFW8iaj1qyejWtxl62vv9/RYBsbMuimEQqSlEk2kjm8d6EudBk5hZQvlz3xhqGXQmEIRuM46Kqy1uwt9gjvQ6qZaoKQ4PugIjIE49Kjedjb2Waphjrr7Wi1xljNCpltyZRkdOnW2/rWllE/5KSvn7RMriAdaNBhFBOgTCQXJsSoo8olK6W95A1D7a1gcK5CIzQ4eI+Rzj6fTTrosE9IWEKSoXsRVL8aqk6X5HmQ9NG0kCRBMHrnebPOamgruXSGFK/r7Cs3WuNMqFmhpkdZ0jh4WnCBcxb4fphW0UUtg0+QkQWSB4adVWtvTtrEBLIre9LIp2nFa9PM+Pd//3c1UTva2mTa9uLFc5nWkUhsrK0LfQq9n/ONzAoDhslDE7awuGiLy0u2u5e1ttakNaVa/NkHA3F+73vdE0F+ryFb+NxiCmSzNjA4qJ+vRCzIRDCYdVmuOjVU+exiAiCxQQMo2SjDWIZMGOuVSZRAnNSZZZBKS6U8oTH3DqDBQzOZmIPUjCjSNJtFbS8LgQoKuKUpae9cu6RmxubWhn1z+7bFGRzDpmhpFQsMWRcGFQN9vXaI4qOr2z755C9qPICG6mjv0hnhfbOHQVhjNAYFHkQf54jPh+wP251hNU1pzrKQvIFxw5miMAZ5SYLM8yJxcy1jGtv7kpKhWd7U3CwUIebYUfIpWbUiaNWUmg+8LuhAoTazuTdsNpmq13mMBA0JwwjddDTmta/Qps1ktHbEReIaZ5TzGw2aud+i/zBax0S6WipK/qW9tVnx8tX0S1tbWhcaenio3wb6+iQTwXNC0gcKfktbm2IO72NhfsVeTs8IJZXFfBZ0Oh4AoFs1LKIgdw8mYntjU6OGK+jmCn1Nj6Cct+62FpscH/YhCmyRbN7yhbKVYe81IrFDse3N7b3dtP4/DwYJD+4WkGzIf1DkOGWbJpjL5vD++dwMEhgwMfAg7nL/OGMg7ayycDkz3Mc3QWcbH5ygj0ujkLNxkM1IMivJ+SyXNSTH68qH3JiqI/eX13M5feqUVWNx202nbXNjSwMKjBelDV0qWLXEnZi0gYFeNXYolPv6Buz/+M//Wc1nfj5o/GIuZ9VCwUb6uuw//Mv/ZJ//4ffW19slyQHu5f2DAzt24rQ9fPzEllc3rKdvwGbml+zkmXN2794j6+/vFXoM+bhcVDDU+P+t+gy5g6wNDg7Y0++fCJnGa1JwcA8xkGfvNzamNIj67tED207vOyOrWHapwpIzzth3oIfZJy7NwCDCDfg0kGlpFVo+8pVyjxZHqBIvoyJIQ2fOXzYvpD7PkvwKNB2sF/kISeKnpEKc4oWYx/eB4qRJ0YZ+vLTdaWrH9LO7Orr0oIsFl/ASIr8E5b3NdrYxPG7VM9rYWrPTZ0/YyPiI5QMrBKDEPjEITyH2BPKhtZiNjYzZ559+LomF/b20zi65SmdXhyN821JvJCMlcRWvt+WlVf3HcAfJH+6U5bV1NccYyB5kcr6eGtIHZp+kGj1vIV5Fd7nyhCD/ouEA92PwX2JQyJry3oulfBiqeTzt7e3yBlqtquFab2+fcjQh/GruS8R9RY5MXKP4f/H8uV7D41G98jPuAHyJIpq+ZBzFcnRwC+vN73km5DYCrxAjYQAyvAwSg2Iu6vfesFfDXZJsEUiEWOmyX/5F0e/NeB90qMJ949+mOw15oCz5EsPA1jeD5R8beEcY1kRDg+2n91TME2sjUJDIKzXyPNf9VxYUr1p7W8rGBgeg9rl0E1rQBpNnV3eQWMVIe3CvljHJbLFc/sDq8AlpbhEYobEhaRubm4pn5CnkbjwPkN3UIZh4xhN1trW1qe8XAxfmg2Tc3F+MIZiqe4p4mDo0Rktla8Gvquj5SdTolmRDHc3qrCIej4caJhog81mTyWY16fUcGIbQaIh7zv7O29fkU7KzvWndnTBRShqkjQ4P6c59+uyptXd22cvp19Y3OGxLa2uqiRrrk9rHui+Rd6FpA2MPDydYiNWyNSfr7O1r520/vWWjQ/326P5Dy2aydvjIUevtH9Sa3r//UHd8qrlNzdIDQD/BoJXHwsDPmZAB1BVytAj5yhCD+E8M4vPRjGQv644TgKgs+bpIFhJTbZo9ff0DtrOzpWY9z1RGpvxaLUkKqb5SsIa6mp08cVTMK84Q5ye3v6u9BDNPPidWZ3fvPbBYfcI2N/e0LxoanXnEfrt+9bKdPnVEqGie1cLCos28ntG+YO1gBILgJ3/jvc8tLCjWE/8fPH5s65tbavLm5bOH76HfauRX7ZFpeNEZwHxFnnoCvlDLBHaNI/wd1czexoOOPBX0PNKu2Uzarl46b3fvPrKO5ri987O3rHewX6bF3969ayMjA/b0yayNjvbapctXdedxtgFNPXr4UE1c9vP1n70tBtlXd+5x81smTb6M3E9eg4rNrU17/P0rO8gxpK1ZgzzOXD1A3kLlil24cEGylxvr68p/YIC8de0t++STT9zHT3sZfwuvZQHKiD0eDGzFps3lNKAHuPjg4UPVfvli0c6eOWPzCwu6B4lHArOFxqHYsMmkWBfUWQDqaLqyhxigiAGLs0sYPBA7GB740AEt/YB+DnrtksANcSxC0BMrudP4lToeWRfyILGSErD/ASrlrVaJkM05a2lJ2pGjE9banLBaIafcu7u7V9JH9eSGDS7HR/4NeIaeCEN1wHkYZCfr49aYqrOVlRm7fvWCLT57bgOc9VLFphfmbWjikORWGdLHqa8a62xhYUneP5RSE0embHFmxpqRQ83sW/oA5m+vZctVO3r2vC28nLX9fUA7ffaXz25aHBBPqSS2UH2yweWbgwygK0h4PSFpMnJA1jPUsBfOn7P07o5Nz8zbqRNTyuHJdZDYI/fv7+m3uZl57Y+tnT2rxOuss6dXLA/qjY72Tp1lBr3yEyPGAjRDySGZ1DlxZnQ1DIZ9yM/eVd/ETMMJYjW1I8+JoT2A2IiZLqkx9VEqGlR4vg+AFC8ubzJrABNklAXWCGBUZwbW6TPLLysoa4glKcAprMKS7kvyIzEt8c2MsWYuLUV/5djhI7a3uWHHJsZt7tULmzo0auXctg10OCM0hT9oqaDcmnVAvndqaspWlldtaHjA7t17bJcvn7ZHjx/bh7/40H7/20/txOkT9ujRMzt/bsJ2t/ZtoG9Y90Imn7WGVMLuP5ixt977yL599Mzmlpdt6NCYbe7B9vD6fmdzS1JWMPu4B3j/AJ64X6P+jAOrYPn5OeK5kEtzR5Pz7O3vS94PsAXMCs4pcRO5YPpCUT+AeMFeIv67nJLnELwe3yNQVgA/RFJQAmRowBFXfhv5WXIfRj055bhi0Dv7QWAqZJ1DM999QoK0dwEAVdaBhAlkl0uSqpXCg7r0EfPe36uk4YNSyv+o/epAWh9sysMrBqD1B9Cm/1lc9SwAL/J+wCnO8nBAaATWJa6J4SpWeMMbNQUAR8QIcnjWAYWZCOjtP4v+Jn0fgDtR3Yd85YHqgmjYzVpyRqK+p+qfgg9qI6q948G8vyMQMvUPdQXgE5pNalu6NJjnlj8NKv5H++KnP/v/+QqMJhK6YDgQaoTWaqLz0WgQtVzo2noliWiyUSj/v+y9d5Oc15XmeTLLZZb33qEMCq5AGJIARRKU1FJLVHdPzEzsH/sh18S2Zlrd6qZGjgZ0MIQv771JV2krc+P3nPsWubP7BVbBYiBAAFWZb77vvece8xhkA4TIC8UXhxAbl4CEXpsoVGFjUwxy+K2vb2kqHfkDuCYc1EUou94k9uLNg5xQGkEWKpoUcjgRGGQiRdCCVSF0rRuqqvFadaQGASZqwjeAbJS8EhIDOZuYGFfQQDZjdX3Vg1Qwf44KfQIKKCGaSn19vZbJZYTc6+rs1pSVe0DAc32+oDMrwz03BSNAuY8FzQNv9OrPoCMCU8OTNZAeJEo0jiN0S2j+ytwuI8aKmqf4CYBwAwnc2qqmCQ0QR+r6+BUUdCqV0ftA0QflGNHiQRUVy87ikIEyicIPaGQX2qzBtMylp1xeIjIm47NFwwBHNrl0lWvUlqwSdEfVqP+hjiDPVqbEjuYlWeZQ7evttixNMWlG+8TdqXowNZBqqNro2Iht7+yo7qQAZa0ylJERbAPTadfHlXcCchuFgg0NDUnOhIEbhwivRUN5fW3dk5dqVete8mGhEyQd4iAvFg0aokGNmplJLyZZuxRxQrQIKuTmxZwbkn5SYyFuyQSDMJeLqY/VbHpizPYpojpbbGyoT2grPjfPiv2FBBGkQxgWVt9oR6msxeob9YsClMJNUgkyYQ5yF9LYdvYBz0vJNojdwPjg+uTdoqGds36ipoeMgi9knxzxRCHBMxa6KAwEI6kfBj8XA4lgrMcelRlekKmgEXFh5B4lmxhe0shCLqvmRl6sGdBzxJyNjY0LfXU3nXItbZ737fk5mQK+/c47dv32bdta21Bh0tXdY//x7/9uq6srRjMFRMg777xjs3OXtcYo0J4+eaq4JLRkfb1Qd8jTffHwKyUpFDaFfFkFifvdoNftQxhHK3hcomCDKsrz1v2hodXfrwJNZqDVqpq9xE4GejLADv43NIJpLMLe6uxB8iGrfzs5OrQmhjjy4QhDQrEqHFXGAKguTlziOdTrM2ezDCWK+kVTi8HC5vamki4kggYH+uzeu3dtYeG1HZ+eWANFRaEsnU/iI+utLZm0/t4eGx8bs9XlFclKdXZ1K0YjvSAfmmpVOrMMPdD6XllZFopPNSzDWTVfXduU+Cj0UxjciYEk7Xn5NVstsKc8efRmXmQGGMUUXo81FGmTRqbdkSlbb2+fUMvyoGiC1kusSCjBZr3AZBDr7px1VrLB4SHb2NzS8EhDsHNYM21eJIkiSwxzNgcxgTOBOF44y8hMu6+n2zraYBIciHnC6x3tH4jyfXSYssmJYQ1WOPe4btA/anqWijY2PqG1srWzY3t7R7a6sWlsZ+IiQ4Zo0C0ZA84LEPf1ZmcycPZ9USnmLVY9t+HeThsfG9L/u+/QmTUlm+WnclZyjxdiiwbtGH43Ja2tg9jmXjQksgxKGIQx6Oa+MejiPTh3aSJK3jAet8MDhkVdFwb1NOoyuazuH4Pi9fV1GxgYUmOIgo0hiBDmqZT1dPcEg+SzIJdS52zCM2/qwtSh8eaFZ836evpVwKbSGenpsi5gRnF+0BTCw8Hl65yR8avffKyh1e/+7V8tnUsLNKCYF49p+NtSX2f/6//yn+1wZ9tymRMxNBiSNiZbrH9g2L579kIyCl29/XZ8krb+gRHb2dvXPmSv0thAjgo2UGTkjfQR0i40nWmE8X28r8v9xTS4YOgSizdY5uzMTjIZO01nZDTbBgo/X5TUJM+HAc3G9mZgmjizTSxMKPaRuThNwjiDwaQaqlwHZ0PEPJAUotazU9qR3CGHofjk2pxRwzAI/eKKGDCsbZ6jhvhhsC30rIwnm5W3aI+cY4LcZPkzkI4lDSCR6qK5RYxmcIkfGajdrp52u/f+fQ0qGJ5zjtOEIpfgdw3uK2Z727u2vramxg3nIZI9E5MT1tnVIZPl45Nj5UreIM1JIgHD3c2NLT2PUr6oayrhg4O2uTxLOF/xgQrGjkE3mZxPGuYyZg8ggyCXKMaMYhBI+ZzOCgdVOIUf2REMQT13PbEKppptrWrO1GpxyX8wcAXFSk5yfHKkPEP+IPmC0KViH8O6gNVK8wSPKEzl82d+r4kxZ6DOCz70Z7jXnHRqf2gY8ho0r2Uc39iowj1iO9Lg44uhBg0gYo5o/sgVNrjMV4TW4+/JN7nn5EXfI/AcbScfDZ3vAX0npoEbyUYoa9fshxngyF18jchDOS/JLTs6WnU2MTgCcEBjEpm8cjmv67k8NWF721s2OXlJ3iU0g51ZouQq8E0BYFTUHKdJz76HWYdBNnGe85T4JtmF4GkXyUZ093TZSfZUZr0MzcVEkzyVDx9iAeiEp4YaKYCBBJYgT3LpQmdae15ITMIjrSnpTAyaAciJZHIpabbDNkwkWy0Wd+kazqO19VXFa1iMEYODfUfjA2ZeazKp+8ZgkDz1zcKSGoHdff22vrWjvZJsahbDI3uWseGhIa0b5HQ4E/DQqKuVrL0laf/pv/7auloaNCx88e1jS5+kJCmDMffe9o4MtYlDSD+9XljSXpGnC9K8rTAiDu346Ngmginy5Pi4YtLW5p5duz6rtcyapLFFnF1b35AJLqj5nr5+DY1glRBvevv6LpCuxAXuKUkB8ej0NKMhIzmGlQuWqItZQ7xqqeMTm7s2Zdfnr4sBWS0wEKjKNwiW3FmhJNnT8ypyiXUWr4cBydChTU2ZmJVtZKTfddsDI5ehn/zHkAU7Zxgyp+fPmidW5mgSNdTb7Tt37L/999/pzDsrFuzw8FRndTRY5bMjRQUgCnRrNJxwRDGpPexhz+cVt4MEUZQn0/+Ehdnb1W6x2rn97KMP7c9/+qulj5GLSdidO7f1uZEWTGdO7ff/9oVlswX7+Dc/sf6+Qevs7ZU83lcPv5TcSyZzbj//xX15bX3y579apcywOfJKLNnPfwmj4tS+/vqZZc9qVo01WEOiwc4KmSBR6zIpGCaTV5MHO2iu327emLfPP/9c+zUyHUayVjK9oIvz+Yuan8BEDAQ5zlmP0TwsUAYbV+bmbG111fLyfXSwHnuQxioADO6pfAPEBK/Y1vZmkAp21nMEqCBnIacuFTnXGJa4N4FiT2DxO0I7ZulMWrGP+MbadXR51JT2hrYDrMj1qWu9fhCQiprRavaP//B31tfbYaf7e9YshYWEbW7v2PbOvu430DQYnuRNUmwg966nIVu2ga4O6+hps0r1zO7Mz9ki0k9Dw3a4f2TbhwfWiz8cTEHyuVCnI1VLTo1H2dT0tO1ub1pXR7tAnmubmzY8MWlwGC/NXrW93QPb2tqznt4h+/zht1YsV+2MBrQkXr35KoaAJBm5R5wVwaCcOjgw3Ylno8PDao7jMZdsbLKlxSWbnp2w7q42sXdGBoftj3/4k5WQ7yNfR3UAKedmhsaw01usWiaXxifAmTaR31LUVKV2FDOH60JJgDgd5GjI2Vij7BU8K5CbPDo8FkALpidxBQADbGTkI1dX1xx5XjV9rmhYpXge5ICiQUXE4vX61w3Z3TfLjdC5BgywJeuI91wAjhWRZyPON+KH0yjJriuzs3a0s22XRodtb2PZbl6/bHub63ZpqN8qxbJkd5EKyxe9hwMbraerR/F2cLDbnj5ZtPvv3bRXr1/Yhz/7yP71v//Z5m9et4cPn9r9+5dtc/XAxkZG7fhk30oMb1sStrC8a3M33rZHLxZsZXPHBsdG7CiTkfKCGFV7ezbYPyA2EvUqPZ7Iz9NZ2XRknB0JYC3qqTDsATjDfTxNpwQ4g7UGmA4mCPkN+e7r12/0zCLZZzeMdtZuQGUGNoGzeuXDKNlA3+ffDyqcES7vUXm64dHqgxKXyXQfKXIY5Vb0CBgSB5amAga5T8jh2MvyjaAvk82qx+X7EHaDA0i9d+gDm++BGf9zAzamnB3gixgR8lYlV/leZp24QO0muTlJPrustedbDAV8oqK+mVirDj4Us7MKoxy2jvcZyacACvK96iNKhSPm8pRmGs6hUuB7xfNW8hjYuHwe6i8Bg849X+Pf6b1EALHI7yzad37unFuN8ykomcCoiMUAhjp77EdGxf/Pm/I/Xv7/+w5MNlP4nGo6LURXuaxEgwIgMspRIKocPqWOAAAgAElEQVQjECWUlPP93gCvqvGHxA6FVjSo0FRbaLZzIbYIAgRN0ecVfL7XfHP9PU8KXfrC5YvUMFagcxQuP6sACzox0H4j5L8fkG7cG/liEGC9EQbVzAcwJO1ujuzBlYSNBEhBQPrP0D6RIqh3jXaKOChroB8xSw0GcqDeCAp6/WDmFZmTQQkHEUcDloYVJnY0Hgj6MBwYAHHoR81+Zya43JGbV3uDgj9joirkfowg3uxT1DCW1lABHI2a5Y5U4T7THPLhiLMX+JI0CygMc6qbJEkiTdDAYolWhhLD0AjXoIcEVEg/UKJNKvZByHJ9kSdFhN4jwQSdEqEBkeSRkXbE2ogGAjTJkkk/AGDFNDVIfiVKmN3ouRTQOqCunIXCcAK9bWl1SvYheAcETT/Rlms1SXpwGKiQCs1JinmGARTGFJp8Tgqz6EBwqp93DtzIjRTSm4kahnEQi0XQqORBMj/VqhpcDEZi+ECApGO6rXrc1zkIY75gjLQn622op8tKuYw1NzZIS5RDslQoqGGigxCEHalIU7OdZguWLVaErkHFSSbSAY2poURYy24K6jqH0SBJBp5B25731/qQjmckC+F0ywg94TqMFfdUuGATOIpBRvRIeAU9yghFAWqQmKA4QSNAjA5nIXF/hAILZk+sTaR3SBjdSJ583qUUHOHu0gM0yZzFULLr1+ZkVAhd+t179xwFD9KFgqVm9t9/+8+2B+K2em53bt+2u2/flb4lTYD+vn77/LNPnZIc6KOYwv3hj2j0lp3FExDPNO0iVCvrxT+L0+AdfeJJibQ8ZdheLxNV+drEMTn1PR0ZBxMvWKv8PUUJt6ACCh3D4XNH+UDxbWtOWlc7vj6hcUX5jmJJYJ15J8vXelOiWY1RpDGk5S6WQqsaQBRhDKeq52Ub7O+xHOsLqS4Sd+6lKOFQcSrS3E02Ntjk+KT99dPPvMBQguPybyS+7777jt2cv2GHhwdqKHD/v/zqS8VLmqs+9HWNYDdE87XE2nJZjSY17hgYOTUb2QUfGrgkU0ZMF9aZy32c2MrqhqMsDXSey3HQCGTYyhnC64JOi2TCIsSVnzMg/Gm+B+3Whkbb3tnV85EefEurEkeQbBS5DDeJJ9rvQRqmXr4c+ArUrKuj1fr7utQ0akwgEYPGd1IDIZg6r5/jb1Czjk7kXzoCMruk2IgkDM2u5lZvbIEI3zs4tL2DEyWgGmjCfGBlB5kwjeb5HCSyaM4iS1DO29hgn/V3d6qBTOwhsiAHl0W+q6tDsg4UNayTQjYvGRQGWpjYssaQK4zXNUjqJ4u0VtDMZ+8xfKDxxBfPkX1HQ1HnEF4k6NGnUmqast+F4G9u0TPk52gi+eCpoPMApKy8YEIsoqHHXtEZjjyFZAGCLFo8Qny7DJU3IH3AyWs6esj1Vnm2165elTzMwvKimk8RLbJWLVsj3iN1cfvVzx5YXQ10LQNs19o/Ps3a/sGJEvqy7r1ZmeFZzc19NWBHVgikYDKh4SV7j2ajhiXFovX39gVwgMu98fk4p+TPU61Z9qxobZ2dtrqxITkrmvdC7sc4D/DWqKjg3d7dEftGpEOdDy6JQJPGBw/EcI+3fA//5tIHbmwsI/RSyZu+kljjDHY5MXKrra0dDZ7ceLwm/XYAJxcFFCyOYPin1wuyY9xjtPeFRNMQGYReUewZH254/EPeZXp6wpaWQaA2WEt7uwpfziSx4NDNllmqM4PKhZKGVZxtPEMaF3wGDD2TLbDYki5vVeNMgi1QsUwqK4PWOiR/FAd8TxwDCpAcHt9XEtrRTW4p1t0MnHWDf0XEopDPmdi4fkYR19xg3BlNNH1hJUn+L+S3HK14JezvH6r5zzkGypM8qiUJa7houZzH867uLjEAQCt6/ur72RmssF4THhPl4UMzzhkOPA+Q0zTSyKHJkVlrnCnyXGAAFxDwOl/0uj4wd2BQQsWtcuggxYTkUnRWyQuMswEmw4WnlhfPLuvjgxxv4Afj7/D3nMWcJ5H/hvtoFL1h5QqZwaQaeTCa/5hKO2uZwRreJYlEgw31dWuNC3FI7JfhJqbsVZ1h9Zyv8shh3yX12ckBuYdIxAIGAi3PZ5XxLnJzkkB07WjtibpzNZaRqkOWBKlUYiSAEgFTAF7Jy4P8izzWhxg0Q9nzDAM0FA4DHQdnuJyrcv3zshWKOcXY7d19SUU1JYl/NGEcpMXzQu6O+Ds6OmIvXr7QsIt9f+utm5ZMNEg2kaVIQ/Tps5c2Oj5uaxubQlnXxzlXHGENqhwmdYQUzmczkjvq7WqRL0H8PC82wPNHTzXMmZmdtcHhUTvYP7KXL9/Iy+Ctu7dteXVN5vM0XNc3Nm18fELnEjHi+vXr9urVSxvo69N5zPUjWzUyPCIZTQZrnBUHRyl7++4t20W6p6XVjk9Seh48H2IYEkmskd3dbV0zLG+kipABYxCvJjDrLJ+3kcEeSx0faA119XTYrbdvWmdzUsMTZPISLR22f3hi69u7li8yPG8TUAcmutDoirOAR0BsIxPqgCTuKZJ33rCtt2RDvYxn1eQkB/+Bd83i8orOwb6+Hts9OLBj5OXYV8jedXUL3AbrGSSv152+l6P6M0LpetPWzyexyRl88T7kqM1NlmxstF8iQfjZp3aWS8lTZ25uxmamJ0L8nJRnxONHz2xoqN92907t3ru3rbO727LpjC0vLdnLV0t27/5tsdg++dNfrVCoWqVU014ols/s5794X3I833z7zM7ysMnqDUOUcyvqnBWrpa7Orl69puGw2EjVqtjlV69ctSdPnrg/iJjgNcmEUUMKWFdfZ6fHx6H+LKneZOBNP+DF8+cBdFCntX64z2AJxqA3k/ldDe7A0Na+BsByzqD7VHHRzdeL8rbx+tnPu4ZGR887GxwWMd/jubeAfIlk0JL3vND7ALAm3ashej7UUi6R1yjpRbxe2IsQflqaG+3de7etXMpZb1s75C+x19jLyytrAtQQ4BgqwAIB/AEIkIDTnkzaYE+XJdtp3J7atctTtr+6ap3UwaWyZJz6x0ZMeHTOcGSVa1X5XwDuQLZwfHJSjAo8S/DUkDzP4LBV4nEbm7liu5u7lkrnLJlstzeLa1bmHmnYzjAGaTh6KigrOLpbQxrV6q46wSBd5vKKe3H1aI6PDzTsZ+/jqZA+ObT2lla7f/++ffvVI+VA2ULJaKE2tbaJ3U/OzT1ua2mzdCqt2hZ5WnIkyTfV8LvoEZMM3yHOGeTBMG3nq6+/V9e3tLSsnG52dlZnJIxohraTE5MaoB2fnBh+QuTQeM6wdskPxSAMflxivQW5o2hQEXmGuh+V1+daN5GPpIbU7i8QsXw4TyU7HEd60OWUOb9uXb9uB1vbNtjXYbmTA5u5NGrZ432bGhm2XDqrvO3wcN/OqzEN0wGVMZjf3dm37p52++brRbt3/4q9fvPaPvrZR/bJf3xu82/N28MvHtvPfvaWvXmxakMDQ7a9s25xzvTWJtvcObWJmRv2fGHNdg6PrKO3R0MiAEjUoEcHB2K6M7BA1pP46v039oL3csTCCyxL1atNTYrfDH2of4mTqHlwn2FU8Nzo7ZGPbayvK49kQO5y5O6NoGa5Gu+A5xouGJnsRQ0gJPEUZL3D/eZ8VbM/sKnY88rbA5gvEmUivwVIQc4noBrAV/OakKGiD0pc8pmfgZ0tJrpkoZwBEYEmlLME0Nv/Vz9XwF1JhHmu5QDeIC1Prae+nqmu1ABaoDrvt0XXwPv5gNR7kup/VZB7d6lM4oP8N3Q//KygXyFGGnLfUqapqsby4YrgE6oVWX/Uv/LyRc60RF8RGWIHsXgPjNzW+5/EVg3nAmjS5aycqc39cQ+OC7Eo99v6Ufrpx1b/39odmAbde3yijyWUc7lsfT29QlDRGGTKyQFCgYFREoOKvf09FX0UijSAoGFysGOMBjo1MsemMHbUYt52dncUECMdO58QOkqA94m+VJwTCEFzh4RRiUkwSYqaXaKtRnqUwbMgomwRUGUmSLMLamiYPIuJEailDE3lJ4EeXigiSVQJDhQxkY4r3haSiioiD+WI6Uw6F8yCXEDOTb0C8yCOtE5BCCMPdM6a4F5xyNHQ4UuIDyVhTplTk+cH5ocRxT5C3WowESRnHKkSdFpDI5Xo6ywx1wFXkAt6ngRYvrgGmv4cRro26Ty7X0FkYi36f5AJUdKuw5FCmPuJjA0yOF40/jCwk7BgnEszzWWokpY6Obmg5EeoOBWGGNFqgOXGSry2G1C7fJcXC/6+HLKRgbckGRi3BJkD0CVK2C4Qlmh2d1h3T7dtb29L/oT7gHzH+tqqGkIkXKCLGFJQhIfcMjwjH1tEmtDcH7EDQFIJqePrAhkKCmLd83hMTVGn55FoURA7DY8Eor29K8iP1YQwK59lbbC3x9qamqytJSEpGiQ3CqFBr0YXKOlyzWKNSds/SVst3mClc14P5GKkLek0Y9alpvgBJRohFjTgC4bmLjXi6BOXjPBhjOQmEk5FZB+Q0KmxgCRZQEkIvRDQl9p7wXhPey0kEFEjRbTDIAH2Q7Mrb9CwzKpWQR5Lg0o/nPm3TjxuMmk3mS3DhPKmwpW5WdtcX7aPf/Oxnhm6vjSAQdH9+c9/VgKu4Uy5bP/lv/xnl0Gr1oTiHBoesT9+8h9CCtIkQg6HZ//Vt4+tvb1ZmsRuNF8nJPqF/4IQ+75vuRckadxzDX6QUsrl7Nq1a7pHkQYla5Tr9cLsXPGQxIzvJRnifYTWTjSJmUUyxcAUn4qRwUGXeUC+rqnB0flJEkOXDxO6leZXxeViKPQw8ZaUUQOsL48bsK7SqRNra0N2z1ke0PSREsODg8JNJtrJhA309SqOoVfcCaIQFFMdwxAkpmL20Ucf6Xv2dnekTY6W5+PHT4Q6Oz05CYakIKe9gcaeYHHRRGQ/MKSh+cJr0WBmmA0NFvSctGXDwELmzpwxSbwpfD1xv6TZTcGaR7u8Kchn+RkUFVIk26CGaKapYAEdLhkVf621tQ2tW3SwYc4RR0GGuul6i2JfJINUODuz8xIeF20a4oBibWx04+kIQcN9HujrV1wr5vIqvhYXlq1SidvluXGnZ0tL2U39aOYMDA1Zc2u7kLTVWtxeLyza7t6RmvzsU5p8MnxjhiTYkCMKJT53XrbJkSHr6Wi1fC4rlLfku5LN9vz1K5uanZJfCY102ANQhiksQYuBVBaNmjgJa4NGfbEY5LecbQhansY89wi5DAa4UYNSTQcVFc5K1PAeajrDb2RTaEZIgsiNh/kMNE8pPimsaARHGvesKZJypImINzIEFiIKmRbkzDDYLkoHm+b89s6WEGNIOnCm0Jhi7zGcVJMVeamkSz20tSStUjizSi5rH713z7qRakhhFt2h9ZDNV+zR0+cyjE6L3eFIxNY2N23lfoJ41JmWSIQzwBujDGy57pGhIVtdWblA5tEcnbw0qb0Nxb6+PmHn8bjtHRxYBmaLmINVa4RFkgEtVRaSmdyIvc1eAenNewtFqrUeGEl1voYl3RMKFxCAmYyb/rKODw4OxaIg9qTTWevu6RXyFcaRYjwSTgXYrS02MzOj/Ip7LH1b9mMBEIXnK+w1H4b6EARWGgNccj9iCsM5/hmWJhIIszOTlsmdBDnAJq0DpCmk9y8JG84hCreagC5dHV2WTqUkY1KLx+RlMTqGkW+rfiFrJRTaOTIsDba3c6B9SxGbrG+09rZ22zk4ND/1KQxrLmkVwBpqJoaGJHGI3I5rkPEoCDyMEWlM6BN6c4yz0FGINF2Tyi96erskL0iBzDpAykkDfK4j0aIYJM+RurgaFwyEaDDTwGOPyPQ3oPai3IvFKhkSWEF4lgW2FOeGSzh6nuaSJS594o0ZHyRETTox+yTv6M08MX2CzKgAIrDwigVdt5gS5y61CZjC5aowx3QUoKQugx+bgxocCaviWw1XH+xwPrP+XL6vTnFQ0jBIziE9UOE9GD7i5YKXVtG6e9BgzshkenZqQihxmpzsLYamvM7JSdqHkpI69MGMQA5NDDE4B1qUl+GrA6qf6yBOATjhHEa+kevCu6Z0XpAk1clJxj768AMbHBrUYELGoeQSgfGNISr5I+himmKABxiG8BnYw9xw1+R23Wfyce7Jgw9/YqdHh3o+i0vL9ur1onXJXwHG47n2IgPDvp4+7W1yzifffac4WMwX7R//4VcCSuCpc3l2xt4sLMpcFx+JxZVV1QfxOKArcoaSGHqO4PcmCNr4zU311twUs1/9/U9tZ3vFpi9N2jeff6lz9ycf/dRSx3z+Uw35YeOOTV6S5CCDCtbB0cmJEM3InyJRyXkJstSR7zB/3auFZmIkOwvClbVMbKHByt5lqILUj2J2fb39/d//0r599EjNUNcbLym3JD/VsCuVsc6WVitlM2rwIluFmTFAKRbk3OUr1tvXb89fvLL27l7bOzqxQpkgQL0Iy33D9xTMqpIbBvNcMlkf1rAPVX/QICqB4O9UrGYIeSFvhfdMYHZ6AEBir1UDz0KpYrvylWnQkJnYxfuRqxDvIiPUqO65QHGH5pWGzUF6E7lDgBV47bF+f/V3H9qnf/3Mqudu5nvt6hVraW225aVl+9WvP5KkHWcQCPM/fPLQLk0NCN3M+pm+MmerCwuKz5wP3z55asVizc4yRTe4Lhbs448faOj98tWqHZ8WrFKrF1O5XGPIQjxF+q9i169d16ACJg17h1g6dWlKBsgMDXl2yG7id0XsJwcTQAhjZtXDPvCgPkBRYHtrW/cFQAxxQQ3SUA+qZqTBmENGBWlWR+BzblCD7B3sBbBCg56Xy7HUBbPbqmWyqeA3WBK4j/tDLONMYP+RlzBw8Yao+0hwfS7DxjkKMIpaErDQuXW0t2qdg2aCQUdu19/fadeuztjp8YHNX79mVckA4llQk5nzaSqrddCEpGTwdEu2Nut8YAjW1dpsA8M9dm4Fu3ltzurwdDkraMD0emXZeoYHdT1kcM2KqWZLCyvW1z8g6d7xmRlbf/1ag0vi0eb2tuTJrLHJuvqHbItBRebM+vtHLF+qSgYNJjQgC/UeJLdZr3OIc1C1cGDDE1PlqRWG5ChftLYkNVje2dpUrdLWmrTToz2L1RrsVx//wp49fmYvXi3acSpnzbCGx8dscXnN86PWFhsbHrXFxQUBFpA7Yh8Sa1hL3d1diqGsIeqI/v4+MbPJuWBJsM/w/EDmKjJedxmoBrFvPfZ4vCXXJ3+JPG7YqgKCXgAo/Sz03Np9SlgXkukJvopi/ktKsKLY5j4FDoJxhDr+HRUBGmCekndwH6/Pzdnx7o5Njg7Z4daqTV8atVI2ZbPjo5ZLZzQogEkMA4hYgccJzWZYyW3tLfb69YpdvTojH533P/zQfve7h3b/J2/Z1199aw8e3LHlhTUbGhi2l69eWLK9VQPFlfV9u/rWPfvu9bJtHxxaH2zt05T851jfsM/I6am96GV0YL4usKX7bQncoWdP073JYyB+Rjs71jfQrzOJ3HBgsF/yeFPTU0L1A4ZgQSBTJBmvYiWAtvw+sZbIlSJwhYP5vFYTSwIgcGDMis0ZjwkYEuUQXIfiq2QzHVgsye+gtBAB/XgG8lgBNEC9px4QwC0AMmXVxuT+yBfy9+xJ+Y1dAJcdWBL9WcOT4NmioZX6Nw62JT5RjyuoBxAe18M9ZJ1IXkrqIQ7848tZEd6X5HfqU2fx09ejX1Rz2fqS944ieSsBRDWA+d7TIqqbmpu93kOOi+8nf5Tk7tmZ+0DGYhcevurtSVrLJSZZE2LB0sML+4B+RMSKlydXksGz9xnpFfw4qLhoI/74P38rd2CmrV0TWBVvwYgP/V0S2zQGxGiWtjQraJAIkjBB22cTcTiSRIAQ82I/qcKU3SpDZZrbJBuGCdWBF+k03AMDQKi3oAfvAwo3KKaQ0cak+AxoQ5ITggTBTclo3JF+bgqHpIwba8lsLbwu70UzhQBL1KGZx6HG94EAEtLv5FjJFAcjU1a+OKgJcjTleB/QdEzjHb3sk21Pon3CqkY7dP9EQkGDICY5opA48D4eXFwCyg9SmgrOyoiYJiD23OinxdKnfniDgKaJS/HjrBZobc7AIO3Xa5EYxUGBOJsiKj6jqTAHkRBA52UhUmm6KXcP02AdfoFOFw0LomEAFYiYE2IUuP61X7Prz/OwfRrtg4syhmrNSQ04mhqa7OT4SPeV+3lw7H4CrBka1mpeB1OgiyJZBbkX3N4Ud3mgyIeBYYD+PqBJ+XkNU+oaVIixXmggUZxRHI9PjAkZzn3lvk1NTdna+pokDDzJdR12H659T7lz1g50R187QnEF4zJng3hij8HjwdGRGnAkhDzTRBNGjsgsYU6MZFSzVYpFJbt2XrJc6tgujYxKAx+djMb6mG1vbkgTkx3RBMvprGTnsXrLl88tk2e9Qqt0BkRk2OS6iTBbvMEMKozn5LJK3jQmORRCP6CZ0Y1nGOmTeDc1Zo/w2WjCUXhyzfyZvehazC53FDFjhMzUoMtNn4VgULPDtcC1doJ2rVM1/RCNPCrYCwz3XK/fkToyQJNWZL1kka5euyIN0OtXJuz9D963zs5u++d//mdb39yWLwNNIj4zcYoE/Te/+ViIQRK17sFBW3z5wr768it9ThhfQ8PD9j/++KlZrWRtoN6R4AiakTCXIoYTSR0SUsTEzc1NFV4gyz968MD+5Xe/E0qZJgWIQD43r8H61r2JxWTOCIrqm2+/cbm3eNz6+wdsbX3dRsbHFDuhpqIrjgcOzW/MSkHQQWAvauiKES+Jd0mIZrwpaMCwpkmUyak0NCxVVBxSlBHyxkdHrTnZaAd7e2q6QetGCgjpFO55S7LJZqYmNRz56utvpGPNM1OT7exMz4BkamZ2RpIFmdNTe/nyuWj+oIxphojdEfYC8UNDCQxOW1rUaHbN8Jq1tLVasUJTznVF+XuSQ34mYtuAcuLMYKjBoBuKrAbjMGdqriFPM4sGPOuFmMDa3tlF6iJuly5duoh9Sp7NtDZ4tgzH0arm/ZA04hmyH4hvxCJiNe/Jnu3r6ZFXSEN9TFrE+BygO51Jn1pjsklN8oP9Q8UqkInEhp4ujITPZTC4vrZtPT1dMgNHCkT+TWJBIUVYtUtTM0ITIwt0eHRqz5+/sBx7WlKBTUJ2M/ORV2JEpy4X7caVWclANQkFnBBKCAmO3cM9m708aytLyzYwMKg1B7NIxrIWU/zDWI9nynCJc4jihudL7KQxIdZLIe/+ETCZ0Ezu6lJMlO9NZNKI9FNbm85vfDjYs9DMKUh5jngcsHf2D/adSYV0WWiAI32nMwE5tYYmIdTYXzSzOKv4Ik6xPzkjeUbNijfOzFEDrBaT/ARrlCalhq+1qtC/SG7AqMgep+y//tMvLc65Ucqracp+GxydsIWVDcViZGUwnF1cXLFbd+7aw4ffWl9/t+XybjI/dWlcr7mzuysUImckOcj89ev27dffaAgKYjhfOLMHH30otJo3hmMWa2iw1c1NDSpgFhDEQf8jpUGMwGySISUSCCCY2axR45B8iUb02PiYHR4c6r5ggLi9taXYg8zN8sqS0FnE7hevXtn16zfkIfHy1Wu7du26ilQMb/kc0umn+VoDResxUigvzoG4azerqcG1C9FVkiyWI+pKMhGGXaOmV12jBrw0vIUMr5Xsn/7x1zJW3dnauZD5Iufo7R9whGsRbeiKs+Ro6pYq1t3bY3tCVRfN4jWbnpnS/QT5rGFkY0IIzlcvXwshXh9zfzCedxwzcPxCgsG3GzqiwVUTEprPydqJUJViYUgjuaYcjyGXml+sp2AiK2akpH3QvI9bd3en3Zi/pryNIpkhxONHj+0sjwxZuxrnSFWQHpdLBfdag+ESDCqXlkGPejEp4ITyKoeFRj5QxEdvuLC2Xf6Oz8KQQcNwPQPABY4sdFah55ewTYl/3A/iPNfJ6zm6mGGsA414DfeS8b3lEk747jDAgQGB1COsIM/nBNSR8WuT9r/+PjLWpkCGrUJTKbB9GRcRH9i//CqV0Kh202nAFvUNDGfqrbujXVrorHEfwPiwRCAGvJZaWmxvd0+5KmwIeRFwliSchegMahjBGNo7MObk9NiGhobVsGFoUjjLqpFD5ra8tCJ0LtJYOTW4XeqV+4SsKGjY9o4We+vWvIBTL168tK3NTQ2i3MwcSUGvTQS2yuVscKDX7szPux52vM4ePX5i3333UrmDfMfyBTs4yNjtW9fEWuDsf/L8mT4z7//u3Tu2f7ivZzZ/Y94WFpfs5YvXNjiCjOmeNTQmrC7OZ3REpbxbBApwRm4mdWrlQtZGBnvt1//wCzveW7POlhZ7/uSZGuLzd+7a7taOLS6tGOkWTL3RiUsaUufyRfkzIT/GYJM1RsOFNcewkmdCHcS1wmwklvuQsybADIyyzu4uW15dly/FyOiovXz9xv34KhUhqAGHsH4AWUiqMQaYywESdbW4FfCWSzRbb2e7jMVjcdiwNIZitr2dso7OLklTnmRyVod0GOsNgEexqOty1GhFz0uAjdAsEjMqeCxILz+XlSF5hO6X/jcSPGENEE/5d6QsiRXNLa0aqBydpG1pZdUSLa1qivF+5CHab5ILCoPDAADyej9iIzvrQohh6hEhWhnut9rf//xD+/Qvn1m16oOKu2/fMcBujx69sLfvztjm+obdvnPXBgeHbHFxMQwTUra1tW/3f3LbfvLgQ93Tz//6qe0dHltjQ7PVKsg7Il1Ttvfef1sI7sWlData0uJ1CcsVz6xSc+Z/LdRPszOzaiy7fnqTJOqIgzs72872jtc7IIbmGkh8eeu5z49YMrAlCz5Yj2SY+P9jgT2Snk+FYSvyX2Kd19cp9rCPGFKura5ZqeIypcQRb0bDJHNJaYYi/M7+ZFACANKZrwwwndHBe9NfIK+P4qEY5CG+afAe6lIYFcQ75IUAKCkfQXI2ZtbT3Wbvvv2W5D0ZdB7u7etzDw4OW49qqbwAACAASURBVCqTFksFKR3AFuSO5G00bsmvECTb29q2kYk+Gxnrt7mpCZNQVM3s+ODEtnZ3rLMfeeisNScSVk5nlB++fr0g9j77/e579+1gw2s8zmR88rr6Bqyrf8DiiRbbXN+2TK5gXd0Dtrt/bKWK2SkAgXNYIy6RTTwTqj5Wp7gd+SWxJwA+MXzlKd66eU1xur+/R/kEw2PIIfsg+y1mDz54YItLq/by9aIdnKSsPtlsl2/M2/NXryVZ2d3ZocHWwsKizvTJyQnFqJ2dHQFTkCQin6d3Ql4imRuYg8TKGP2ChAMCqlVdI0A0+ZcqtuNjBlPOzzbiN2xL1irXz98hSUX8pjaRb2Fg5UcAF7F/AsCSprGj290bsbvLgSecoeRPfFEjwbyBKQeL3t82ZvNX5+wslbKJoX5bX3pll6fH7WRv125emRIDGVbC5uZG8BOjrwEDN2HpNACdhK2urNuV61dsbXXZ7v/kA/u//s8/2p23r9sXXzy2Dx/csI3VLZsYu2TPnn9nXf2dlitWbHPn2Gav3bZHz1/bcTZn49NTtr61rbjENedSabEw8MXjviNZyzkIC5ZzkZjLoNoZJo60Jw4hRS1ABTUQ8buzQ8PFS1NT6n8MDQ5JahVwH3ttampa63x9fU35DM/yB+Htoq9F3cjrklcRIyNWGXEWnw/OTxjg6pth/B18FwR0IOeRJ41/4RkEk9XHFDEHOrW0OnCMQUXId/g+ck735iA2+StInYP8P4A1o6FKNPTymODxinsm39oAutVVBEPsKK5IApK8SGC4hmA67gwtV1Jw5rGrmbiPaSQjHkmi8T3EGvkfhn6n9wL8drKG3ULG+yL0RXk27Bn2xcrqinoCI0OjdnJKvmSq36iN/TrovXiPh5zVhyt+P9hD5LL4c1bKRdvc3HKfkh8ZFWHF/fjb38wdmGgi2cupWxsVUjSrSDopEsQwaHBkOwkDaEYkMSg8OCAJMjLt5EBsbnZUJxR1mTo6khgkNAZgkusJXzKYDNPWaMKuVDBQ1NXEaWi4oFHp+kLxJCPF4I/gSChPKghSEd3U88qYGlGRiSKJGg0bij61WpW0O1VeibHMhB11RzAHoeXT7DrL5jI6sC6MrGQO5j9H0K5UfbBC0SMNdaa5MrQLzVx9HpoArlvM55QHBlNsmUCBnHBZEpp3NBMY8nixWNKzoJPl0jpRFPRk2f1CXL/d5SJAHfhAKGI9UKhAbefwiFCVXAOJhIpmSaGEIjkkAX6LQIq7tADPnuQyej/um4x+MVkT+hkUrw+cOCRoNoCAVPO6UlFhiYkuE38OLLJjmlHcK79WR/i5R4kzTiIZHjEWuEZhK33AA1MGai9/L+R1Q6O8AEh0CfZM+Emeo2umIFtbW9P9b2vvEL3SUYw+secQjJrxzhjwoiUytBQSPOiiahikJmiHklsNf4TCNxmSIgnCcwUpxblFYkXjd2KoTyjgarFks9MTVq2ULJc5FRKPfaNBEcV8W4dlckVJSp2kc1aqMExzZAOPn7UiU/VgrK3PEPNhEqwMN1VyyqSjI3y9yQhZVO3vUZtq3qp54cadzrgIdEPMfikqQhIRUUW9GRPkNcLa8aTE9deFaMD0FK3XYARFY4piUUOQoLcqKmPw2KAAhVExd/myZTIpeVPce/cduzx3xQ6Pj+z/+N/+dzUd+ZwUPzIfOwEt0ipd9uvX59X4AK32+vUrPX+ahsjxsGZp9M/fekuGYqL/ytjeGRCuR5+w27duWd/goP3H73+vYoy1TMLK8+Wzcd+5N9xnBooMCWhEbm/vKJlnbfPxPQ54DKJQBdnfCDVW+volOzw4sK72DslSsfqg3+M9QIHUiD49xX14P5rJxC4Sy2joSLMk0u0kgWuMw3IiRnjDsae3Ww0iqOxQqYkHIMvo8RE1dvf2ZbatzyXZvHN5EEmbF6Zce7saFjR+fHgFQssTJy8UvThA+okzgOQx8njhHFADoclNLSI6sCSKkLoBLUKhgpSIzFV9jSmZVGx3FI/iSGOjBkGUYPgfQdWnyOM+UDBz71hTxFqat+z9d959Ryg5mVMH+TOGcJxZnG38nAaj1aqawitLS5LhQu5jsLdbg8POjlZb31hzY1xR6l0TmXjGc0dyhEYw+x+0JA14GB/DI6PW3pbUoAtJB1h67JPWtnZdC8bteI1g8AkdngIc5oP2rMywidvCj9v81SuWy6QMk28NR3p7rViq2Mrqshq9aP2CJG6UhCHofUZdNAu9gcN6YYBL44EmfGSIR4OQzyCmXTDajQpDzkuebUdrq/StGUTw2VPZjBo80aCD/2cfs8cYKOELsbe3K5NhCk9+DrRhJC/jEmBugMizJe5T5LJZGEYR0yiAaaRQRNIUQXKM4QbgBKSMHj/5Tus0gQwMhRqm0aW81Qpl++gnd8WEaYjTMMHnp2gtXd22f3hqS0srOvdgsoBqnrw0ZSsr6xqmcb8i0AENeu5DZ0e7ngFFPv4UaPNz/rrUUDAojlEA5+U70tzWZlu7e3ZKo4u1UourOca9RPJvfGJcEhuwRfBkIt6htz57+bLlMs6GYDi4t7OrJhyNTyRCQLLy+RlUQOHn+eLpgakwa41mwejYmBDffibjJ8Z5V7RzcrfQ8I48f1z+x8EhynFAdp0VDJ1y+QdJEso9FmBJ8Bz4LDyrmZkpSzTRwHO5kyKxKO7IRaTbonvIuUqzw3MGs8HBQfnbrG1tWV1jnR0eHdj45LgGMMQdeUbIQyxh66sbMu8G4ICReXMiaae5nPs2qXFFM95jjk4amWzXKaay92Py4iHuBmZAYLixtpQ/wSgMAAQhMxuRw6zofLh3/x0Dfc+QEdQng4qjo1MVyi3NDOOIryVLZU5lyMzPcO4Tl2kaRQOIaDAUIfRk/KkBvheWnLuRv0TkraXYErSaacLzLNlbLqfnkp58D89W8ikMwAIL13XKHdnHviY2S7ZEOaYzA2kuRTKgFLsM14llksEKAKVI8k1SgMEkVUw1DLfJGYt5l2W88C9jkIH8isu/cf62tTPwr7Oh/l6d3dQL5D4wKjAgdfkyb2qSBzpTxMEXDJ2kXS/ENNKLVaHBASTwTLhukPNIbfrvB3b71m27c/uOffIfn9ibN4vW092lHIpcygdzwYuknnM7Z/2DPfLNYNj/8uVLrVtvSDhamV9IwdLoLJ7lbHx42FkhADYSSZlhP33yRoNQkPKsy83VDZucGFejaV8NdqQ06jSUR4IRr4vxiQk9w2++eaym6vrGlqRHks0diuecg5FRObmMWGT5rJULZzY61GN//8sHZrWCwAuPvvxW5+HMzKziz+rapq2u7drw6JD1Dw7b8WnKNrd3NVTmOQJyYMiGXwyAD4bkNDdAxsM6ZuhAbCEvPj1N251b85bNnOq8X1nbVm6PXNXzZy/UuGZ9j40Oi7UFGrS5KaH6j7y8udU9UeT3gV9L8dzKZ3nb29m2vr4OOzza89ytpVdSiGelsoa7wJ3qGhutSLNRzG0aghgiI/+E4T1DC5eNJF9z6RLyFM8FiYuAMBz4kFBNoEE7bLaxURsbGZHEiBjsyRYNKA5PTm1kdEJeAchCnaRTloP5pLzG9cL5klTMxdf3gwonQNJ0A13gWuctiWb7u5+9bw8//0KxgvP3zu1bqpGWl1fsg/fv2m9/+wdrb2u0X/7y5+4JVavZlw+/tBcvlxRHbs7P2b37b9vLV6/s8PjUAO7mcyV9ptnLkzY9MyZj662tA6tUm6yuPmHVeM0SzfUCrvHcJN3I/cR3LEgvCxz0A8Y69+/o9ERsTs/ZnQVBL0DodRrf5xUbGh5SvIGdwe/kTuPjY/L649yOJGiFeg4mu9TO5FU0G89r55Ij8wEQsYp9Bku54n6FeGRm0gEAhzxKm9jOYuNqUNKkXIB8yq8/NC3jPlDRUEGNy6rVNbAWiEOtkg5L1LvfWlN9XJKQ46MDNj42qDPwiy++tGIRydibQeLnUEANXo+mOewVmUbTfIUpz9CsI2Hd/R02MzFqpzs7NtDbrxhA3MjSL6mU7WRv35phfMRiahwODo/Y4eGJXZqbs403r61FCgpxxeD6RLO1dvVY1+i4bSyuavCbaO6wT/7wmZ2iXU9NLA9F6mAkJ2FhN4u1SD3hZWtQUvACVusQGVwAGXV1Fevv7ZXkWRt700rWiVR3R7c9evLMVte27ThTsPpEk3UPDNj+0bHX80hPIrMqzwf3R6P2j95N8lqSA/JnAaCVGCDAaxXViWYfkOu8ctAcMV/gAQYIyO4AtAwy2fSM6Isw3Idto6E9Pp/IUTLsP3fkeyioHCARchsfKsKsYp9izO5yhWIcIDdadt8qzhfuo9jaeF+em81NT9tZ6tRG+nrsYGvFbl6fs/WlZbt7fdoOdg9taGTQdra3gswmLFty5orl8+RHcfmu3nzruq2trdq99z+w3//LX+zGW9ft88+/tgcPbtmzJ2/sytxVe/3mhfUigZc/s1w+Zn3Dk/boxWvbPz213oF+OzxJiXXO+Z46OZV5PXVt/8CAALIC0SFdFRrf5JSSLkSWtd79o/ZhZ/T3q74iPpI3rq6sKldEYaCr089igDh6FpIrHNX+gg3DmSUQgkyloyFtUAQJfSD1hwL7QnXVeVXDBXJmKUjQrwsDJobN8v8JXlcyOOe8r6/z3A4AVamk/e/eCt6LcwnBnEBUDA71mfWsfTjMlwDKofHPdTuwgT6Zs6Si/porxDiw0/0JXcpN/ShyHNjhwUCcmlRMz8BwFntJjIqy9gT31K+3UYwcFAI0pJEEHXLxDh6WukAAX0smVvfae6gXrJIAFKUmoXdADc7Q4ujkSOAJPDrOJMNGP8Ql4fmMHjPJfN3oHjYTNWjEGFKOSF/qx0HFD87sH//3b+IOzLS2q2mmgirIwQwOguLPih1BI4KDBcQkRSeBTbr8NDRioH0Tmr5z0NAkxLzY0dve9CQZY4ODyFSzQpRNR4iSPAmVqOa6m2dHiHACmyaiXlYHGmhNyQCNaTVSgzyLgo4kjaCbnQvdw2eRKSTUciFJ69U4BV1K8ossUCQngXwBBa4X8TEfUtQ3WJ5JfLGooE8w0QHJ4Ym5V9qZEVECRkKmhl5To1CXvJSQZpKzcd8LPhONzQh1J0od8jnhnhBwCLaamiMNI9kMTAgd8SjNRdgo0l7Gy8AlfSINPSVzmDEGyqxEHdQg8mky95+AGwV/ISDCQUASoXt67jJV0sSMKHoE4UpZ90W0OBWVNBu90auDVL8jUeRyBiDlW5pc1oPhEM1Mkh0NKUBvxZzC69ITfCZ/1iQv52WnFvI+oN3VHA46iCSk/GJt0FwmaUPygXuNfjcJIAgZsrj2zg7XWQ8HKAVvJpsVugB6HahVn377QagrCU36qNnhjsCeJ3lR6/R1GuXcdz47PiQ6bMPza2iICdHW0dUtRJqeA4ydxjo7S6esoyVh0xMjVg7az9D20PKmcI7Mrju7e2QyyK4oFMuWyTmyTweekrg6UVPjsIuktyvSoxsDqkFbJ9YK6zYyiibxj3TM2W9cszdDQLEg6eKyXNyDaNjkkjw8i0iGCKkhDORh1LB+aOA6UlQ7VXL7Ppxw2Q2aMJ5kxKUh640yIYSKDOACciqOH0zJLl0alybq1tamYskvfvF3dvnqVaGaH337SIhBEh7WOdfOGgYRv7u74yhgfZ46Nd1dMoA1GzQgI5NQ7XXXmSd+8YAouhlI3L1713Z3d+3FixehaCPOqB2u580HJKGJaJ0wafz+elIjrXmK8eARQ5wDXcL+xyi7CZZALmvtra1CZRZyZzKZo+nFkI202lEzFL+uK84+1HOSW7tHRGesuQya7ve5J2MMyTBubEwgOVKCkiY/D6ESYSKVCtYA+glqK4V2eFYaXskDx5uYGtJW3CeHLw0F0NtEA7fe0e2sJaG0g5musxTOFIM1c4gTp73IYsgL8jdqBEhCSchglxEgGSTe5ZGmSDZLWoj7qfsakCjobsNkAZnN2sMzgrWFASADBdDbDEORrIBhQKwTmk9SAn6fGKZGklqkfKL6MkRtQzboxK5fmbV4kGPLMiSwmho1eFMQJDgPkCPhi8KdJlwbDDGQrLmcvVlc0b+1tzXbBGyu40N9PuIfe4amCIUcPhWp07Rtbe9IS1x8EJo7FGo082s1e+f2LcukjoUsJelH27QxgYzEohrHMmvs7lQTnHskY9FKVWgpkJsk4jwn1jWsl2iQTUFCE9hRqy6FEw1e5QsR9Fh5JipU+XfuE+y5c2SdvMHJHiSe4wnE0mQ44oNlBthNygmE4tY+4yxAYgJtWDSxHU3X0d7mzxPTvmSThoY0V1jrNED5frTIYRG8ePnGlpdXVbwVS3nrwBCveGbls5y9e+cta24ElY1UWl4I5XS+ZOmcy3lIVx5EUtnN6pBvgf3AwKUCQk0xjyYZ8gqhaZPN2dDQgKXR1VehVZF80eXLl3VtFIfEhmRru23ubNt+iN8g3mjg4i3FvUVPHiT2xua61hkx5/jQG67sZ2KvpL3yLoXHOkVeQB5cDKUL7oXDemb/cN1CEMMu4BnAtkSbV0CQmhtOE08jxGpzc2CyutcYXwAUaKZq+BhYCMlkkxf958jwNMtvIp9DxrJeBpWcU+Pjw4oxPC9yQK4ZdDTNcZf0c1lBPhPXA4qP2EJDkN8lF5NstLHJMTXA2X+sGSRwUsdpW3iz6Gjfhiatk+NUWgNeGBXsHQ26pAHmjArikWMKHWnqnh6OaBMLS+AH8r5idMB7Q43hQAPDdpCnfXb79rzt7e0E9iHyp/32zTdPLHWasa7OHtcZjtdsb39H7ByavWLWHRz6ALNyriYX7xudj6wnkJz8OZLKdNkSZyqwH30QwRAsSBYA0w2AHeUiMvANjESSypr7pjHk8/w3yHaqOHYTWr4irxMGG+TxeBYRo0qwZhJ+jmnwJrkkil6Pw1xLdG1CXtNsqqtXM6pmsDJoPDnjDY8FpUcClbAmy9bT02G9vd2WTp3a4MCgmpmuc41cm3+OKB4QOzg/GVBGuWpkbi9TcsBAofmpBn6lpOcJ4wng0/TUlN28+Zbu71//+qkQwEheFfK5MGAm5+X+VcxirAOXdb18eU5rfn/3QGwkoSmR5Gpy1jZNIbGUz6s2ONiv4TPPmkEQA5enT1/ajRvX7fbbb9sn//p7nYHOEDI/t0oYsiOndypW9ltv3ZT83Mrymm1u7dizZy/ci6kBXLbvWZhMnM/OmoElfK5BxUBvp/3m4weWSR9bb3enPf7qkQ0NDtvQ+Lgd7x/a9vaeff7wiY2OD9ul6VnbOzxyH6v6Oltb27FbN6+rAQ47FI8uhhOcV2owixEbs9GRUbHkaKqMjQ7ILwR2LkOUVBp982YNTjlzGVDMTl+yE6SkOttJizSIGR4esPN4SQ0U1SflmmWOUlbKlWx3a9MGBjEgX7YGYlp9q6RNjzOZwBjOW4l+P4NH5XTur8bzdiALqNekA0uC8SjyM6xTGslra+sabEQNLeIfA9B4rWq93d12eXpKuTZn6OLCkmoUwOe5QkmMCnLKnb09ST95PuvMQJdH/WGZ/4NBRcjB2Agxq1gjbPfGJvvw/fv2zVdfKmaylicvXdLzxFfkwYfv2u//7Y86fz784J4Gszffuqnm/OvXr+3ps+d2livaBx+8rdj39MUrKxZguZSEWr56ddruvnPTPv/ic2tswC8l4QAm/otXBIrwAaWjgKnrWbPEJoaVA/0D9urVK53ZUpcEpR3qaPeXI574Z2Sgy14jh4Ep8t13z7Q+2TezMzMaXBDvotzB7xKNO4xnY/Jwk5pBtWK7e7vBoNYbaTX8F6TD7g1HziRnmCHR401SAeuQU2mkrutQz0FNeTWuI6YFAElnE0vip+YgPbwQclmvwRsA1jTU2UAPsnEZMScHhwftT3/+s2UzVbtze86mJi+JNUw/gGa07h0s+WxWtR35ch3xrQ6D5Va7e2velp49s4nBEcXBZEeHNXZ16H1Otnesgil5oSgPB6SfYO+PTk7a4daWJTRIPrMsXkAoPCSbbWRy2tZXN62MF0my1f79k7+o9oNJyCDp4nxrYAAKoKam16SekjdDnF5J3Jl3dTG7cnlOg7Fksl7MDkBU4+P91tXeZDPT03Zeqtqnn39FV8UMiSlpmdUL0KS4gFysgFFnqklc/sZlDLkn5NORJyGfn7zINfS9ZmdoAbA10vVXLK/wLF1amB4IeXm0Z6mHyEOLRQfJKb8J8kJcjzdg3czeoeqhjgzMfgBa9JwEuuE+wCINoFgG4w5+hfUVpK6D79/VmVk72t21kf4eO9rbsLdv3bDN5QV7961rtrG6piH16tqq8kwY0f19PTKQR92Ctbu3u29Xrl6x1dUVe/e9+/anP35t87fm7cuHD+2jj+7Zw88e2Y3rN+2zzz638ZkRq9bFLJePW1vvkL1YWrLjdMb6hgblgcSggnokm06LtX14sK9YiR8IzXsGogL0kqPGHZTqJH6/F4C3AGJSI9DboJZCLm10bFS1MYwq7hGsGHKQCJAZAbCcDeNyuDxPcvWoB+e9BT/nI18EyZ1LhCKShvKaN+qhuEm3G5BTFzow2IG14Zu8vxcxDUK8IUcnZ2BQGF2bDyh8yMVXFJuj/hvXTj2pGIAsY2ubs42QypL3lfcn3P/WYwf5MvkF68wVIryfKOBwPV6kfo+kKpFwaWg3xMbzzCXpotflvPd16ueFszmdMS/QWThE9OfQu4h8kATYpr5HXq6TeiCmPcf9pQfL2b1/4FL75FCRcgvbgJwb6WNACdF7ibn746Dih4f2j///t3AHLiWaFbyY/tFMYwPSyCVYQdVDg5VDhyCJLIf0rLNZTXGjhg8DDA4f/h3UK00G0O1qQCV9KECDicDFe0hTPxTkbGL+3ht8HixEIywWXfNYhYYX32xmGkXeuAM5GBgfNCDEivCDjuKL4p7rJqDznmzwnq5uBTI10TibMQkV6oND0nWw1RwDiSTtfp+ISge4hBSFF2g0auTvIDSPMwh4P4Ifhqxu0B3TFJvmsDS2m5tFbdekOPhkiEotBBaT6HrR97g2EH00QtxPw4tVyewEveBIqzHSZ47QCjJ8DvqzkppCmxcdQxAhoZl9dHQiejv3UDJUDTQkXbNZ90koc//M7s3gJpzRQCI6HHk+/IzQZlADgxlzNeZGpjTJkpgKN4G2zdpAf5/uGQcQmp0UHZo4S4697JqF4TV4flFzncRDElOSaIpYF3VKpDThhkUTWA98VpAmoLKa21qVbILWBI17cHigBhyBnKTgzeJiGMzpiPl/bmUlh6Hrrva/D74c7e33MkLX0gjwpntRwwiKYb8vNFHi0pTngKFQaqqLWVdbs50cHCqBvnFtQgc5DVdoz27si7GqG9lSIMqsulSWfqnFGqytw58day2dywpVB7KUJA9PgkQTqMaEzJtJzDjAec5q3ATtYmdL0BCneYCMiiP1HUXAs3cJguiwjYaCF5JSwcQtks3iNVzGKwwQg78CzU0a0awhktFiCbRHUYeuo2Kcwiut2xI6vE12+/Yt293esqOjQw0b3nvvPV07ifne3oE9ff5MDXMaaUipgH7EkDaKI3ROImoozSR9hqBhqcYOZrkyP3c0l9hkgUbO99G0Aq28ubkj6jRrX82edEpFFl88b5orLk+D0WdShQn/TkMDXVc1DsN9BgEsJCyyOkjUlUu691wrhuTEP66TplatLq6mMkUHAxexoBRDMSuOTMvdSFSo27BnY7F6a8MwHuZGY9yl4AplyT+BzCK+8gtEV0uyUY0/GoDEUDUGmpCly4hxwPqm0Oe6NVgoV6yrp0sFMc0wil6XWmJgm7K2Vn7me/8BpPK4z6VyUY0jN85t0LUxdOTZ854klGwr1h+viYaF+nSxWNAPj6sRQbyTIW0JE8Jt/ZmmPBr8mLyyzvxMymm/4A1BQe60X/MGYpDJExsmgexGnVBvYgpBUc9C1++wvu52GxsetM62FiWIewf7knBjjdMc5FlxlvGc+Ts3hfQzbO7yrLRGQfCfnp7otS9fnlb85XlTbNOwh0UBap4EGEkLkE+rG9vS6j63OjXPWbs9nZ3W3YG2LGgaLxIYRO5srduNq9fs68ePrHd40AZHR6wFFgASi7v70rE/PT6x1kRSkjrLi4uuZUvzmEa12Gu+JjT4rfhe1wCagRrmwW0tYkOxvhItSLKc+tqv1SydTbvJbY2mjuk5iHJfcWPbvd1drQ0o5fw/RRJnImchBpcMWDGQr4JQl/58o2SNGKjQVKSpxpmI5BO5BfsNFPubN2v2+s2CNaMdnc9Ki7qUy1r6+Njmr81YTwfySB0Wr3NmE6asDCqE/AzMUIYSDLRB6IPgzp7ldZ5TlDtqE+8fCqyS5fMle/vuvD377pmGoSAsM9m0Tc/MCozA3k8k2jSUXlhZto3tPT9PKUaszhKNTRpAd/V26/OhB460CjFPhSJye1k31SM/cWmmiqQPmhrc3J6TSQ26oNUNk4q1JukivG1iMUf6BfYq10Rs/N5zI5iSB5NlGqjkFjybSCKBc5Pn29ePfrTHKKS6To5TGhqkT9PWznqwc5uanLBS6czKNZcSg9XhXiI+NK1UXPNc2sDxuiA9ktC9499pBh4eH9v1G1d0nrNPWlraNGRM1CcUe4l7yArIJwMz33TazoiPyFrSgKCpz9UEw+wYcgIUojS2QzGt4hBPKNh6+LYIZVl1tHUMNlaT9hUSfAzG529etbO8D51pLne0d9rxUcpev1q0ocExl8ZrrLftnU2xmHgtclvOLthUNIt8cO/NePk8BJN4DbA1uC4qHyOOseb5fjE2gyeP9qLqeWcyOCgC/Fws6Ll77uHnQIPnrmrmwUJ1M1JJchYwwC5eFMjRuc6AlZz3NJ3SvRVbN5hhOpLQ2Y3EWoZIkZlpZ1uHHR0fSmZKwxDkC7q6zaog3DHFLhhHY3NzQo29oaFeb/w31CvGLPT/sQAAIABJREFUeY7sDBHYQwz6kelk7RCD8G7R4BkmNx4Ure1iu9KkJF/zuJm8kAtBXo/ahDODuADQqLunxzY2NjUII79lf8ACcaYtjN+cmEC9PX06I0B8j49P2sOHD4WI5X6LZRMY0RKZCGbksJ36BwZ1ljBEffL4qS0uLFp3V49ySZi9PE/VUHhewQZAZzub1jASA1k+HzUBTffHT57JwLdUiVl7Z7diCv1hl5fLKP4UclnLpo9tbKTffvWLD2xh4bka7i+/e2mjI2M2ODZqKwvLhlF0OpO3oZExyTymMWRnWIg8F8CpegZVaa1L4gISkxgmR6hU4l0PcqBiW5LjVjRkYfi/trYpZOfc3BU1+BXXq1X72U8/svWVJTs9PrLhgWHLZXI2d23azsoZq1SLkuFaeLVgrQ2tKG3q33t7u+yskLXF5WUbmZyRkWw2X1KTFPmneEPCssjtgdKl8YTUoVW1313yxFHYajbB+OzqlE8U+eX27m5AwnrjFnCd4it5Wme73bh6le6WbW9vKuYjxXPGXgVFm0hYS1u73hsPK/m9AI7CIwjgW6gpvUD4QZ0Ao4M/SmoPIB05U5N98JN79tWXDwOj/dxGR0aUy+fOinbnrav25Zdfq6J48OH79vDhlzo72YuX5y4rN/off/iDEPAd3V328NvHli/AHmuQJGJdQ80+/vVP7fnz72x759CyGYbuJEAMHYpCK+dyZd2TmzevizmM7w/NawYHV69etU8++cSbkUgxMfgWsI21AgPQ2bXFvPs9sBcGBwYU53j2xFbuDbmvZBpBzgeJlR8i5dnn7Ked7W3JWm7t7Ih5xr4DjMWjcRa9M+ElwYsES8Kbr0IPB2YNf+Z8293b8+FyMIwmvvL3rG1nbTJI5sjB+LjV0in8oxpVW7Ymk9bRmrB4rWyXLo0JxfzZFw+VZ89OT8lDBlYtcRaPnFu3b130MPb39i2dOrZKOW/ZfNpmrlyyq7NTtrmwZG00DstV29jbs1vv3rW2znYfpOCLVyrb5198YVPTswJCkJPubqzLcJ1cA7ngrr4+6xsasbbOHjs4QE7bLJct2lffPDU5MdF/gA0IOERs3KTyMfyvpC4h2S5nF8hMW14N3ijd39u1s7OsAAbb21s2PTVmxwebduP6NevrHbS//OVza0xiXF+1AioSsTo1PGlQc/ZqUOXoPNVsNEVVS9XFVa/CTudc5Rzid+RYyWtolnvMPlaeQt6r/pKkrmsyfD46OFS9wfoBUMew35u5DgQFeMEZJNlgekVSo/DaNGqER6b2Om+DKgKDNNaSgAMB7MN5yTqgFlZ/KMR1vufGlauWOjq0yZFB21h6ZXduXrWD7Q177/a8rS4v2dDggKRdiTXZTMVGx/p0pmuYXKvpM04wZFpbses35+3Tvz63+VtX7NtvHtmvf/2RPfn2O7t2/bb9/t/+1SZnJ+wwlbdUtmCXrly3r55+Z/unKZufv2Yr6xs6lwCucXYDYkO1hHBTKBetu5fzFOb+iNYB4DbyZs4S7iG1NUxy6hqeFeerolUspkEH95fzlnvLNfNFThyBMjkLGC5RU7rEk3vGkn0qd5EBdTBuB0Aa2FnUamJKyNjbwaIuU+WKJJI8B6Qk5i7SkICdMLZHLjgjALFAJQE0obwp1HIyP5dflgN3fLrh4KZIxlrrIfgdcv0MDMr4/oVBjCSyOdeCvyvxkZ+PZO6VY1VrOuO4ZvUK61GP8DyS66TXoJ8J6iTk4T46dMCFM5OT2hPkY6wNzyUc3eoKHK4gIC/f0P8TAzrkavIC0xAngHAkn4bclPt+EOOIfwy0+Tmul1gYSZgKfBxD3aPTY+GPg4q/hdb8j5/hh3dgprXND5XgA8CGBHlC0kKzkOSWxMObGlC2k5rakiQSvGj2cfCj0wZqS9rTQfdfxjIyrTmX7qiQc5GkR9CBi+iANHwi48PoMInQdhEKiwaLDJhEg6eZ6qgMGjROLHQ0GwkfRTwB0BEcHuQ629oUTEiOiHkkRiDwJW11diakIwUFk16CAPeA/5cnAmZMFdf5JQkBtS70Cuaxavg6Yhfdz8j7gKROutoXbJW4CsgLkyFR7Pw1Kcp0yIiCDsLLm68q+ITCc91dGdYGSj7TdZkbgpamSEI3UP4THiCjabsmzaLtwQChEeaIcJISvofgJjQSDRQNYEj6HA3KTRW9DiS5BgnuLyBzaRlh+2GkIQpsl5gj7znEMFuiETMxNm4352/ImAo9Z3QXya/5fhrr7vEBmsZ9LiRbpQTF0YHcE9an0FXnnsCABkV+BemcasnXhJqIx8eSIuGAB0VLo5PAToDnMGEYtbO94wawyEoEPWs/B33yHulecxhQhHJvZKwbJBj0fEKywn1nj7BuipJXcS5GHchDBkBiHzSoidwQMyvm0tbZlrTG+Ln193Z78n50qKK3s6fbXny3YKVCxgaH+uW9gWQLmsQWbxQlGtqhI4FJRjArLlmeBk4DTAgTIpv+DetM5szBnDWS79LQpAyNsax17cMXR/ELSRHWF/uLPRL5T7g2oicmkYkbxXBkehahBlTsxmLaZyQn3sx1+i2oGO7lRcOfYU7QH+Xn5mZnJAWzSzO6BgrM9bbR9SeJoEBC3xq/CQY0bxbeiIrpiFBvGikJCQMCkiXt/8CeiJI4Sd7QkATpESTGon1A84T/Z2DBgIc1iAQB6ygqXnk9PhufEwQZ61HyFWGQGUlm8GcSQujWSGG0tHdYvlS4MCpnj7DW0UOlqQYTgHjJ840bsgJxIWChhWIQKvNp9lrY/5FvC4MIYllnR5tl8QgC5ijEcKNR5qJ6TZKqVOi8YoP9vRry0PjzuIHEnsuOaegUfiF6VherF6IoVh+zekm/OOqNoMsz4R6TJLvqqCOeQNarealmJTRZl4UjvqohKyNF9yngdyFf+L1SkUwW7BZ5wCBFkM8rAWN/8T4kbKw5niF/L5mJpMue8AwooN66dcuePX8h1CR7sa2tQ4w+EFwMBoh7xFKKL5gFzdLaTlszDfOuduvt7rBSIasmORIlL1++1vXzefjMrDHFDZ0vbhTvw6tuq4s3WHtnpx3uH9iz5y+laT8y0m8tLQnFHz4Tvj0gRIlXmIqqmNs7tK3dA9s9OJFeslgM8ZgQeDT6+axxGEGFkpXR0W+ot5bOdpuYnbG6ZKOtbm2qyaMYUAKNW7SNlXVLH59IvohUnz0idByAAbHQkEaoWWtgxrgPkYMJzkouCcSzIn5S8CDp9PjpUyXFSO5QgNPoBN3KgJZmgzxikGuK16kpyT0BgeaDpSnb2txWcYsvQDp9Is8gmnk0HjkPMDYHoctwTPufZmylbB1dvba8vGVff/tIa0roOIQXiC/lmv3k3evW1d5iKyuLQvdiYMpgF63nhYUFMTspoBkiyWDwJGXNyVYZzoIwB9nNPSb+RH4H7BfQbSBCoVhzJjNspelDIUXsRW0NxtL69pZt7lC8Y6jnZyfIN9V38pupyB8KwAVNIMyIYShw38RWohiv9yGEzvowvGRvkhtowCTPJJre7iNBXNAZivRWyGPkJdaIbAoDmO/PZ3IU8iI+A40sXg/WRld3l+IakgNIVG1uMSSqs4GBYdtY39JgCZ+GbDplrS1NYvrUN8asrafDhyyYGcL0q0eGzyVjGPzwWTjrOS+6e/rUnJAGemO9mAszczOSB6PZxPeenKTs+PDETjUcqVMRi2zB5199bfXoetc3aF8gqaVchT2nYTxnng/JNfgNQ3wnSsaEQFTTJZi/skadSejo03w+ZyMjgzZ3ZcbSKZdwpDgkbg/0DWtQkc0ieQITqGTHp5gSd6kpQM6rwdzevjdRgwQBDRcfRBT9DA1IQoY+Ua4UsTAicI78miol5Sz87rEF/zGQ5cH/i6GLvCFc6lN5Wx0yaTRUgwRTkMvk5937wgeUytVpZDDACOajytMCo47rwJsh+hmxdGGCNbdoL9JMZyCCnJvrgiMJ1aFcg8/IXn7vvXtWq5U1WGB/iJ3F0I7mv6CUMQ0XuH7WDnk4Gvoe66OzI6ch0db2roZJ1Bcu61rnMjZIJCKNJMRnvdjcxHZk8UAwc8ZzP4RURDKhBpstaXW1mJ0r33VpLdbe7MxlPeulpUWdK2DTuV8gG1OnJxcAHTS/0ZpnL7LPTo5PtKYwEh8ZGrHe7h7r7GIg36j1JBka5bfO1nEJjLLQ8jyDQqEsZtibpXWrBJk7gEHELM554nE+m7FyMWcTo/320YN7ljrds/6+Xnv+5LnAP8hhAtxARqpA/luP2WuLlc9r8pzhnCOOA3hAQov6a2xsVMhxwB2cX8j3jI4OKwbDtNBws1qyVOrErl27YV988ZWGjfPzN+3pk+/07Ev5gt2+eV1SiYX8mS2/XrTxsXEbGOm19BnDh5RNjI/beali22t71tHcaaeHpy5v1QBwp9Eq8TrL5PO2trlnQJTQbq9Dai7eYGeFooY/MLIddFLW8AHzV7wMiDfEVMBOknOKgegGCACD1D2BWE/a/1azzrZW6+/qsnw2LQAJ/04ekUUSmPwLWc22Duvu65W8KPmfS254bRTltf/zoIJznBqFeCiPipgpF3r//jv25RdfKrZzjiAzCEADZtb09Ji9evlG9dH9+/fs0aNHAiwcHB4pF3rw4H09m53dHVtaWbaz86qlMnmrFNGBB2l8YvPzM8qjP/v0kcXryEk8L6MB1gBDrFKz1rZmuzQ5aRvr6zLlJlYAshgZHrEXz1/oo4gNrpwfeWKXMNHZxTkUpImpfdnrXK9ytvo6samifcBrEDMilLzrscOOxQvHfZioMTDTpgZiqKmYE/M6VSaxmCprf+OZ4awr7i33X+dd5VzXDiAmYmRFSGuBsGA0BzAeco+UH7Bq+dySLqQHQSNfmXDZrl6dtZGRUXv06IneY7C/3yZGR2xlaVHAusXFNfv1xz8XeIR+hpqDhYKdHu9bV1+7zV2blczz7sKi1YqoDLRa6ixn53UxsWuHhgeUW+WQA5bnUMx2d/c0FD3c3bZWQE35M/lPVGP1NjI+YfVNLba5tWuNYlg1WDpb0L/BIOQZIe3FPY4Mjflc6okoVwm/yMnVuCX2xKyzs91Sp8e2srykfHxwsNdOj7att7vP5ufn7bf//DuL1SesUDFr7+qxppZgYo6hcWDUbO3tKY6Pjo6o58Ngh+cHI40hmEtENmm/ArTjDKaZzvcyyGK9MHwGAMJzZPjNoAIGFHkKwAieD+uE/SoJRZ49/o5qUCPV483oSMZQeXcAcETofPaazpkA5FRdhAya+hMKI6FPRJ/E83jAPLOXpixzcmSXRoZtfeml3b5xxTZWFu3Dd96ytaVFGx4ZscWFBdUBx8c56x/oUvxnOIWxNtc9Ojqu/HD2ymX74tMXdvXGZfvii2/tn/7pp/bNl49tamrOnjx5ZJOzk7a5e2CVWpMNjF+yp29e2e7BvnX391kmixy4n/XEWCSBBQRGihy/v3bY9+zvRqHsWwBaMWDUnzMOvlRtERODFXCbwF5Z721Fyg/4mEXAWveL8h6Re56i2BCBGT2nk9IC0k1BSlqAP/wuxaCPCYyqIQK5BsDekE9EvRH2rwAdGkyktT+I266i4UBQSV7iNyomDK8PCxf2pj6CMxUuPCr8uaoXQeCPmWRaOcu5V/QKGjhDwuemBoXF7+wJH/bxPsoBNfDmtZCjcokpsc8Cez8agIitFGQDI9Cykk/yM+SvJBfvORbnJ1/ewwrng04hN+KmQ0mPgrycYc8P2XqKbUFWkxgbAXXJ8yPACPeanF9DspPjC5NxKUwEjzTdtx8HFT82+f/W7sDlNm8ScMBFyHoMFCnCmNRSqBCUOHhApqPrfHCwL+YExTRNIumZ5/MyPhMtTjrp3tShgSb60j70tjafGlJMBuNul/IJckNBgy6a3vr8FNkSp+8H76ULRgbPIpIZoSCNvp+DUTRAGus0/0KAoilF85HEB4QcmpR8rzcdHeXhw446JbtMfb2gZSKKRI1PeB2h54msmvkqyCpiTIC60/tDv21pFWLP7YQcoaUmKSAYZAyCphyB3eloThVzTT2XHCL5oyiSvp0SMv97TXOZ7EonHDMiZEny+h6KNdHQ1Fh2Wq0mvEHPlYaF094CfS0cNn4sBAZHoORFUgIaUqHlDxMieBZEKPoLrT4NLDjcMDADmVOwSxNjwH2k5U7jAe14hkI0M0CQc0iUpVXshyK/HGzqhlpcY4TG8AGGS0uJXgcLBipstWb9fX2S4+KQo/mytbsrLWIZeEq3vUmIlNXVdRmD8nc8C2nmq5ntB2MkG+GQguDToEQJKSyX4uGeeGPUGTwyqZXkApIfjugQWycg4GmscdbiR8Gx1YTZXHertdC4LSOP1iEk9vsffmDd7e32L7/9b9baklTSghEaSTzLjHmbCl3QYKKnn0vaB4Pdc5AjjVDBObQaAxvJzci5ZtZx5CnBcCeiczpuwuW8fAAWGXk6jTrap44UjWSdaMyX3YQe+Q2ovbBo1Kj3JERNFBglYSjm/jKBIeRZp9axhl3n5yryxsdGZe4l5EHxTEMAbwBxXyvWjLGi6OmgiXxwyrWzZmiiREm7mCKikLuES9Qc4rpgJihBCw0aDS9C04d1RsHnchy+392oDWSP6Zn4cItBIE0wBBx84YjFERB3NFhJzPh7JXXBTwWWiyS15MMSU9HCfQA9JOSvdOJ9fdHUcmNYp+17keB+Do7+aLyI17w+z4I1xr1BP1ODRhmYc8/9Z/gs/FtvD81JjG29EGevRU3QTpl1O5KRIpzEiESX54F8BteqhBIEcQHkHU0oX4u+V13OTdqgJIhB/ov7BbKG+BHpyup1iQWB7UEc7unqDGwKlx/LZDBO79bwhuEUeqsMK8UAq693GaWQVNNsQpaFOL67vy8ZL2jvXBeoLsW2gNBkuChJFhXKDIZoelfs0sSotbUkLJ06spbmpA+oJF3iTTXQXlHjCaYYCDLOSu41z4lmCehemgkkyLvb27a7s6v9gIwQxRpofyFGg8n40NCgzhsK03yxIiQrsk6YM7rhqz9XijdiDqaq7967az39vXbeELeTs6wdn55qMErhXClWjC5Mc1PSvnv81M/PmAnpir4tZzqNYGKoe/C42Vs0QBSqWtJCFEqwd2AdgjzKq5EtqTwa5wwkC3nr7u6VSTTr9s2rBZuZvqTijfU2NjqqQaI8rtrbxIzieylY9w529Z6sDZrnHW2tYvSwDijAWpvbLhopNEaPTrP275/8UfcWmShkQPBkaayP2+jIgE2MjViyCa1Z93vC9yCXK8iPpV0JvtnxyakNDg3ZhgYmFA2YW3rzUpKQOaTHEn6vg3Ys3Vg1/hscDED4It9gKHOGaWBrmzebYIwQV6qc734m0FiHfk6simjoxAcaknwReyJ/oAh8ISCGABfe2CSPSQVgCEXp/v6e9GkZ+DiyHAR5oySyQGWz1kCCoi/O8GB/j0YueugMgfdtampCrCDYC3fu3rE3r9/Y/sGxffD+uzIMbkrADpqz7757LmNH1uqzZ9/Z1blZvef6+qp19/do7xHfV5fXtObJiZDDunbtmp4hjEYKWHIS9ohyHyTT8OJqbLSZmWmZynJOs9Zgrqyvb2hf0pij4fnVoyeGDOLu/oGVA+CEs1gADpi0yoOIpt/LlkR73FuVjsNT3BG4xfM1YhhyGeRMgAJu3LgqnxVyQ5exAhRyrqYJMoA0xGlYc+08AxnXhi69Ykhg8jGQks+DmFaeTzlzgYarS/vI9FIMWY/nFPySMZSR/bka+5zK3pzyARXnGWtULMFgFqrzT9vQ5Rd1bul9nJHhcqEBkRh05zXYwm8IEAwsz0Y3jidP5ysCZTi7laF/XPJ/MCXIDZCTGBiAHWtq1LMGvEFBPlV02Sea7W3NlkllNOiNPL5outE8Yegj5hDDfRpYknVys2eeJ6hSYo3OwTrYNQ4KYJ2TkwhglHHpVQfNeH5GLOJcAxna0YnpNQhzl6MTAyfkJ7CJlL/J06BZwyakJl0O0tm9SBbyXCOQDvdCzYNwjor9VCq5/wFMxeaE9cLAbGiww8N9+WaxN3hv/CGmp2YFbuJ6aaIiPbe3f2zpbN6OTg7VWARdLOP6tlZLn55YMZ+zyzOj9tOfvmfVsgOjnnz5rfV099rk1LSGFMiGvHq1bDNzl629rdN29g/s4OhU8jf7e0d27dqcEJkbG+t27/59++brr21ocFDMge2tXZuduWTTM9P28vlzxeaWJJITKXv33fu2tLKmnYUPzssXb+xgf88a4w12dW5KZuY/ffDA/vW3/2JNjQmbuzprLR1NljtL616/evHKhgdGrLMNTx6XfdncXFPT9e0PH9if/vKprh3pmfRZUQOb+sakzjHOUQZFAJyIj9SeND+RYmEdwgIFiATLDWASgZ2mcqQTHtVVyJTRNAegxrMitqvJC0utWrPTdPr/Zu89e+vMsj2/RZ7AnHMmRZGUROVUqtBdne5gfMe+nhn4tQ1/NL8wDNgGLgz49sy1u/t2V1epS6ou5UCKEnPO8QSeQOP3X3tT8h1/ATeKjYLUInnOc55n77VX+Ac1xjq7eiSbJHBAYImxbiIq9v+z5g95k/ZaMF7FOPxnX9y3b795GEznzQaGR2xza0eSeP39Pfb6zbQMl2/cumEvnr+wO3fviJ3DcIK1M3FpQiyMucUFDgcNt9hnrMOGBkyn8RXLaGgveRKYe5IKoXakwZuSf05k58WGI/uYvc7+53MCWKAxSaz0gbb/G+eug/sc/gfrlbMbnyEiKddIzoO/FntIfjnRry40H8mbGOaDCifaAgZwyVePUZwT50PSEIuJLdTkkuyhPpa0q0uxOZPbm6LkJo60TjpbnIY/YDq8iswBJMQ34hTPGpBXOlFhzY21AoBdvjQu0AKMW/YAOVF7a4vNvX8vfy2GxONj4/aH3/9BDXq83srFvHV1NFp7R4uAYtnMsS2/n7VGWP35gtjJ1fW1quNoKGu9MZSBMUB8TLPGM7Y9Ny9jbpjGBe5HImmjFyesVKywlbVNg4dZIUAa3oTUxyBtKmVCLAanfNjwrguediWvlTlXWV/eLTmz61cnxdxsaW2yrc111eQ16aS9n3ptrS3d9rNfPLB//Mf/03b2M5Y5PbOm1iYbGBqxqal3Ome6Ojp1z/FAg+1GvJBvh0zsz2xocEj5NeuenxMgQJ4TZ/IH4Tkha8rwkLisXDf4WDKwIneRckW4Xhgf5DnEH85+4pw3jB086ed3GNYzqNS/+f84DyRDxXAjyMbxfXo4fBFn5SvKgQWZWGAtpEyTdmV8wnY2Nmy4t8dW5mbt1rUrNjs9Y7/6+ra9fPZUTJunT17Y9RvXbHNj28jTqT/w4CL/ZKjZCmNhb9faOzvF+O3r77MXz97a1WtjNvuBoXC71ByqGPzj0YffDix47h3gJ1QmkADOnxp9N2RG1bMAcMQglHM9yT2stQsjFxQbMclG5jAylzBoZ+8ARCJGsr4YaBArVfPjkZCmpqxUns33WEucj+Ss5GIRbCXVBYE7vFaPjE8NDFQ/OQjHGZ+xd+d7lK8IaCb/A0TImcrzBxBMPwxVAdX98l714QFnv4NeiV9JAaL0/BNe/8aehJ/L3rchl2L9EPt0RgdQBXUzZyg1lvxVo0qEFEUcbMm1KycBZVSRUG2pYUiQYZW/alDRiNJN3uv7yLik3+HSncGrMawpz7d8+BNrX9ZdBGh7Te8sZwfe0qNwmXUNYdQfZF17D0z5X5Bkl7dYwmNoBGBq3eseulE36/unQcXfWpf+p89jE40tGiKcTxArKlwP++BQhUSkRLFRKeBB79GIpxlN8kCywGGPbBGbh4PaG6KYCoMEZEJeVJMHNLsa+tI/RsOe4tH17GWshyyLJsce9PyaKJh8wssmjqgNIX8DzV7BiC2KVmUZOYVjIfzUgMAgSPR6U5CmKKMw4SAVVU6NakceamARJrkkaAQ7NSdAiijBgAEASq1su7tIVtBkDRp0MAgkZYScAMyCCh1ONGlACxO0+cwUYTqg1Tx01JvLCnhS5g3hKMsTDJ0lXYVRkNPQdIAHvXTdI5rQwVDMkXje4I9GcE5x8+YyxZOekyRxvPGu+/pJUcxrxP+EoA9myNw/EqUYYCNy3XX9/Jm5/jmo6BMhryi2NlZXJYMFkgP0IaaE6C5yOJ9heBUm8hrAcFgJVeGeHOcyX1DamIDL8NOklSzpDXTUSyWtweWllcCSOZaJIAF8fXPDGhuaVDjS+EO3tb2jQ4kRBTXNJv7O4SfmkIpln6wLURVihDegeLZuAsdaI+GOBp8gY9U8xghM8h2gbWq1T/hhmSCBDgHffmZWm6qQ+aM8RtDfpZl3krcijcj6pJLnk6NDJcUVQq/7/QWV4LrPBdH7q2rr7ABaLuQX9gjFBOuOhAhIuXSsnRUUzdtpdrBB4yHOZ1QSzCAlyOXwe6xJP9D9WbCGQC1E+R75iQQ9dxIF7ldMPOJwjIaepILQn6WZzYEajYmDKRZoA1CMNL0ppniNyMYQSig0e/g9Ne+qql2DMnw2R185wkISGGF4wvN0WSvXN9UeyONb4B4watKbU8tBWEs/Ei/zIO0lWaXAXuF7SEqAjgPBgMwFaAwNkaKGp1CssDpC4SzNaUzlvOkTkWBRa1KFlwa6Lv3kQc/3AHEp6qxG0255bYQkVqbGDMLCIIg9WV9XL0QNa4mE5pxNEhhT8g6orlL806BVEiOg8NAxLku7GgQ8xWdDHahi2CU+YCqW+HmXJTlvnstXhvch1tJEP1Why3vwc/ki6Ehkojx2RdQ3GuM0otiTjjr2feY6+wwskWpyXxEkaFpbOoVCpcl6lEFCjCGLCe2GnIn0bU/zOrNoetHIAjlOEgpStKUF3fKsBnju0eONYG9cBshVqWgN9bXW09VmtdU08SlIT1Sg43UDalb031JZskrsA0fy+GNjj7h0IENEPFRSQuHDnKA5BwrcpVfQAAAgAElEQVSX2Mcaxj8BRgHP2OUKTOuql6ZtQ7Oum+IX9sL65q7lTkn2Uxr4EhsvDg/Yr379tZ2c5m03c2SrW1tW0LC/QkgxNIhTlTTzTuzVq9fW09kpRGlHW7uG7wALGFho4BR0br3p6WcS8Y/4y1okkcbPhEKTUuXgyA3NOcPZaweS9Wi1ocFhnaEMGkFzcu/IE4j7DMdAPHd1tsubQYzHkyMbujBsI8NDTt2nKNMZHjwWEi4pgFQEQ1kV4sm0/eM//h+KacS/lqZ6yayAOurr7ba+3i4xWPASQPKguqpGgyUKM/TWMfFE8gOPpK3NbZ3PfIkVpIYHhSFDBi9yodgP9PXb1Nu3+lMDlONjm5yc1HvihVSJ9EHQ1YV95MwrH47T0Cb+0yCjySrt7VP3emLfiQ5eU217eztaj8TM1RV8EhLW3z9gc7PzQsrVN9TZu3fvxCRjj3M9NFEoMBfm5oWIpvB7+eqlXb9xQ/vs7dSMfBeIO+/ezdjk1SuS4uDsQFcZtC3nIJJUb968Fqrv5z//yn788ani6+jomP34419tZGREheaPT5/ZpfELGrStrq3q/UBSooH8ww8/SMKEZwWA5dKVyxq8w7qVcT3FZbEgSSXJfsjjpGy9PTR5kcpkeNVpS8uYae8q3lSnUnbn1m178eqV7e4fWe60aLkigzOaUmk7PNo/Z7PJr0oowrAZhQllAEtocVCMBnGB9elFt8tHMSSrb6ix/j6at+6lQHNraWnFjgAAwJRNwNZ02QI+l9hNoNuaAfkcuFF98C+TljDxR95QMEGIrwB3vEiOrL/ISlV+EQYLDmLxPUje6oOx4JsQYjgxiyYq+88lBpytGJEWGp6ocS86pJueBy81AUwU650VG025uR/xvHaUoZuX+lAuFPCnyLr5MEreQjUuyURTkJwY5CznKPsoVZWQpBdMKZow5NLkWjUM11IAK44UO7nfQlaDJgVpCDAlNEwZzEWQDWckTRi++FmaYbNzs4r13E+k/ZBzQ5ee+EZcZfBLQ9fZzOQ6gDd8fbD+/Kh1JC6DMs4JXs/XDYCivBhbgIR4JmJhq0YIe7lYkF/DnVs3Fd/Y3zs7W3rmsM+od7gnxC0atqC4Ga5wnvkjr7DW9m4bHBqx/+1//1/tJHuic4pzhUEsUqGlQt5Gh3vtqy9uWzazL1bu8ycvbGR41Dq6un0osb1vv/v9I7t6bcL6B4bERHnxalqDWxhTt27fkNQRw/Jf/uoX9t1330qKiuc0N7to4xeH/CzKYV5fa40NNH8PNXyF3UAjjWcMq5CYmTirtP/m3/3GVhYXLHvs0qN7e0fWBBOxrdmKhbzt7R7ayPCg9Xb3KkcSA7qmyvYP92x+cd6KFWk1abe296zEAPoooybWccbZpmLxVpoaxzCnYfwjV8ZZT94ngFHOfUDw0MD3R1Jo8vdwaT+WLYa0Lc2ez7A/8VrgTHKQlPvCsFejjj2xki/Wj/sBRVRvSMxCLaDnpy3n0mxJWO3FM+vraLT/+A9/bx9mZuztmynb3Dmxi+MXbGt3T0yX3r5em5qaVr6HDBMD0Pv374vRwzDAa8eiXb9+Tftlc3vL5f1kkl1lF0ZGhPKenp7S+QAAhToy1oNey7knIvuC9cZwzpUFYNxUS1aRgQSfjwqaxmGUZtMA/l/VPfiawL6FFcC9RQ5lbOyiTb97ZwUa6WEt86fy1TNHziMZtb29JaTv4sqqgyLEyvCamdqb92P9cL3eQPVGtbwmQk7NZ+N3ffjrSPuYF6u5GYbFyvEr3RePWHJ8jD8WgAO8ZgARJi13cmCXr4yLJcl5yvoYHxuTLM7rFwA6ijY0PGjjF8fsz39+qM/R399lsx/e2RcPJgUs48yVxOY8flMNtrW5qyb+0FC/dfZ0qylNvVZZrrDDXM4GLl/S2oTxVNjft53VFdWwO0cHlqyqsQvDo1bMlW19c8dOTqltkzY1M2sHhyd2dFLQ/SOfEEMq5PzUkYprKfd04XmKYSE5VrMHD+7bu3dT1lhfY/X1tdbS3GAV1BTkgORhvX322//r/7bd/WPL4QeZTNnY2CXV5fC42T/UQM7Y8AEW910+PUgcozBAfYvXUUCQa08G2SH2AzGD8wHgiZq2sJDlO0E8BW3u5wyfhXVCncYzdw9Qb+xGX4DY61ET3LzmQl2AvgoKEeoNFf0e6NhDnijIPHk9Rt1UsETaAV3egK8U8GJ1YdEmx8ZsYfq93b1105bn5+zevUl7+fKZJNDfvnprAwODOlfI7zlH8JVDajmbL1lNXdqOsjlr7Wqx4in+CPViVSv3KxQUs8gBOFvYf5lcxto6u6ykBreD/6jZ3k3P2PT0jO655zPUyl6jMhzjc8Lq++z+ZzojYLRwz1eXVyQNCrADrw48Zfidjs4O9Sl4Xs58haHmjX3kYxn+EgN5/0PihDCPXsumkrDxEsp3tR+DlxHrjzNebIoSQJ2s6mnuJzWqGBehYULM5Wc54zVohNXJ8CgA7VgLgKXo0fDs5ceKTx0+KAdIyxblGcU6F4DKSQz6bFHO2c+JCqlqCKABG4xhbADEaIiFEkcARcvbQrWfDyoEYqmskO8I7y8gghGTTs794rQmASuHNS/AGOBH3RMAqS4JHgcR0bMnAny9xk5oz388NxwM7Pmb56LsMe6dpKc0jHPwlPKOMDThugSUVd3twGNisq4xDDoEwvyJUfHJSf3TX/8m7sBka4eSdIKBdGAxdiRJzWTU8CLIsIFJpEBPoXG6tbOlwM0GockL8g36NY2jKFnkTUSfpuMfwdQ8siKEqsBsmcFFcLJXI0/NxoC2VvPHm3h80TAU6yFddc6cIODEgoNiEl1KRysV1PB000I3M6yocK8FITXrmfondYiibwv6gmABKieismkmKFgGE1sSRpJI0Pgcii6pAxrUEWtiYwQjZjVrRVE0oTKJsCRBKoBAk+AdAaU9Nr1JmGvceJvmEk1Q7jPSRlwrxV68ByRkFG58LoI6qOUo4RSD+KfJo6MzvaFIIuGMkJTuP89XxajkuHwiq/sZWC4egH1yLQpfdc35NP3TwluFfzih8OqoSiWtq71dDALkFJAp4VgAPUmTdG5+UbIZdOiOMafi0AqyYOc+B6CkYMCcHOvZc53cZxKVADfQcybJlNY9RlRCQZmtra/rvfYO9nWo4rNC0s/9olhlEEdyxCFJ41dTcTFZ3ESPe6Wpu1iNrkUYKYFOOZRTsCNZit7YA21OYkFySxLGoSKZGJrmEIADjZEGrKR7QGDX1QhljhwI79PX0y3pHvTy8RKA6l9AO3drUyg7CliuE3kNEgsSjDQoddgh5Qrdy3JlUneIxlw6WeXo9TDUY9+xxsVcyaNJ7zI/3FsOddYUiRWfHTSGZCJCg5+mtQ/Q3FiKv/vnZiDpBtxqNktD1pvkQlqdgYo/0tqOxUyUjlLfgLWP/BAU8zAwZHBGUifGSFh7vHgcKsloURIAyJY5wybqZsqEXckeTUPXdwQVyzXHBqRQmnkSG2eogKSWXwu6zjGmBAmNbAYpEMwnXeqI4UA1QwoZfZIkxOTYh2qhhFXsooElWbYwOPSE2mUruGYaJPJUYUgWhomuXw/awu+xCoSGRg2CVbwFrxbFgZJLAnAd7GkaI0LEBaQGfxIvz5O4pBd8JF54BLght+97mF8tTU1qdHtC58mXTMrQ+W2sNyowfl+yacdo1noDzhlQPqTkTxpUosMi0xa0h9GpjsNQH3ZUiIEnWZKIchHCD4YM8a5s+3v7ajQkk9WWzRZsfR35pmpdS1UtjS1kUAqiDkOFlTZ7LmdoioP488ExpmPuP4DkHG9Aw1rDoExexabOILb1GWdftdVWp6ypoVbNFdY9RbQbl9Vpb8D4oQm0sQ6Do01SA+x3l28paECj5DxfsKrq2jCwqNIwYubdjLT/e/o6ra+v1w4P9627t12a7Eh99XT2qJhqQ2qkqkpG2yDdtrf3LZsp2cRIjzU11kkyqLO/z5L1dba5v68hJUdkLoO3UcoW5hYVUyk6QSTj45ClCUYhiMZ3U7NtrK07GyygdiKbTBJ/okefyZRd91gJe1LIKM7F2vo6IRMpeDg/OEtJqtE3BlEMe4L1SkO9keeVhCq/rX1KvtDZ0ykzY4pZjGMZkvEcGKJkMuiE19g+w0MNP6tsZxcT5gb7z//8zxoAE7N78RJpalQTc3VlyTraW2xu7oOKtSNJFdUrJmM4i+9HBYPr9U27OD4hrwtkNjjHeaZHx0dWw74unVmdWGwp290+sBvXLtmzp880ROKL9QpqjrXGmmtsa9ZrEEuRLgJ9LCmg06INDPbLdJRGLhIwNJhYQx3tnTb9blr50OTkhD1+/EjPaXDIpUHYx8gr/Mu/fGsDA73W0dlur1+/1jCAvITh0/j4mPbis2cv7cb1qz5M+PFHu3n7lvY0zMV79+5Kd31qetZuXr+iGDc3t2DXr1+VXCf50NzcnL5fla6wL7/8yh4+fKgh/5XLV+zHH59ogMDZ83bqjRgQBCDyJdYIn4n7hBb37Vu3bWV1RTJJY+NjASF54GdIRYWajTx7zjuQiORm29u7an7IeJNmVX2d8qCToyPJAF6emLB/+eOfbHv3wNI1dXaczavhx9nA84roPUk/wKwJcoiSPwseYgwqNPwKrELJUwZWKrKOFPeViTPLnNAwB8FJA+VMxS/5KVJ7ff09wUy6Qs0/BhS8Jo0Azj5kL4hnNLGIP2JfqkBlH/k5JXS2bDO8AUCecC6nKA1uhgj8rLMFI4JUZ2ZAmPJc2VPkLMozzmU3HbgSEXmc7WLgViFF5PKlsbkU8z3ugZs/gtDzIb/nP369XDtnoRqeyKiaqRE8MjSks4hnyTWwHmg0UBsMD49oQHF84qwLWEYM4hjOwcoiHnFPYSHFfNblEJCD8eaMGwHXBKnOJjFkBSoQShb9aGfBMpSioXx44KatDAJ4nsjUEYcWF+bFjgFdyrUSy8ibXPrJmU8aVGvoCfihRtJCIEzl3yNJzyDJCuNZ8jkwcc1qqtK2t7Mt1DLgjgsjwzY3N6szC0bb8PCAckzWB4M76ivyFPI84s/de/ecjV00Sf+8nX6rxvTW1oZeH0Q6OSBMscGBTvv5V/eskD+UH9vrF69seOSidQ4O27s3b21v/8jqG1s0HIBNKw+B9g4xMFlygHMYbNFoHhsft7dv36rhBfBlcX7exi6O6pki3UWTDQnEes475BGrqm11Y1OMuXfT07a8tGbV6Uq7ND5m7fjvZTL29u07S1aB6D1RLtzejrRX3u7de2B1tTAjDtwvJJeV/CGSfS9eT0neZnB4xO5+9rn9T//z/2JJACrpatva2da6Ys2yDhhEM9gS0yaf1/nj+9lrBvZbHGTxjKkHyC9pwskHDI+qk4zAI/xJ/ssa4T65txvP1r2a+GKPsWckoRMYrV7oxyFoLPsdD64hAMlD6czam+rsv/sPf2/NjXUCMzz8yyMrGkzAI8sXzqyzu9M+zM7pbGQA/PLVG3vw4J78P8i3WXOs5StXJtVoxc+DWCG5kgCCuXz5inIVkN2SyrEKnZecw8Q2clVyzpvXr2ugLa+GRELD7OamFnvy7Ok5IEGwKZXbjpQWS12SWgDZGLabZL/IWxaXlpSnsTbxd3k7NR3AQXEg7HU7slEMjsgBXfopaRvbWxpM8vs8L49J+CH6YMiHrpXK76kD4r2OzT7FM8CKYWjqQ2GXY3YWqDPK1NB1JRoHatF8pXFnZWuorbJERdEmr0zIn+nxo8fKKW/cuCL5sxdPnyk/uXnrhpg6xDEYdn19ffb0r0/tN7++bW1dnXa4taV9vb26rv2ytb4TVBpqrKev17X4Ey59/HJq2savTwpE0t/da0nibblkr189syIM47pGDR0po9bXti0bWNlT72Ytky1YJl+yisqkziDWBWu1RN0PQxMAGd6TSAGqlgFVzp5I2a1bt2x66o1VVpQl80rvgz9TZyUbHOy3vcNje/joB6tIVUlyraq6zuYXlm3kwqgPt+jFAKRE+rK1RfkMcVxgqmCgLHkbhuaZE+VjLqftfkU0w8Wy10Ax656Y9BHKZscnWW/yImsoGe28bWysK66LGRSAqbGH48Aib+hTG8HwBeTgtU0435LulcE9ogahTo5MDEmbSU4M75JayXZRk7AWqXcSEFvOynayf2JtTdQC1GaAbVk7zhpvbMRkvcE21ndsaLjP1tbpdTXavQcPVHvVN9VL0q7yzP00GZRxzkiyUyAb9xg7zlBzmSVQxjBqqzoNbRyoCwizbH/4wx8kC4g8HUOmKHnF98g5e3p61O+A1XL79m3t+7dvXmuAjsQhtcr7D+/V36CHRH6ChyMxI3r/9PUN6BxeXF5WDiZZospKSSwLLCAAoU8cqPfVDwq5BtfkoAZTr0CSYGI3evNfjfnKSg1YGWry2hEEgXcotTbrVCoJRcBh9efy6wXkqmHQ0Vtkb4faFpaEMxvY3M6oEONKgKLg65n2OOADMa7fjbCp2fGKi70Or6HJF30IRBxhMMCN5v5wPe6PcqYBNz8vBqyekedfPjh1Nr6rTnjfjC8NsENu+BGMVKN16wBNr7ljHa/BSajXJS0V2Byn9KEky+WxnzOKnisxHqAgXzKnl/qDg3h1TpDK/TSoOH8eP/3lb+QOwKigsfupFn1vT4+S961NGg5Oy+cApmgFzUShgnkSgZHf6+joVEMHejxshkgf4/doxkFbJFGWIz3arehkB2S/gmeNS4JEKpjLOVVoGuwIbze7VtAMgYMgwAEkhBg0rGoMiN3gmyDrNDH6Um40VSi6ZIf/HshGR8Zz/SSuFKlxMOGNP/S7vUASyuwT82dp7hPsQKwH6RlNVCNKO6CiY7Nb0hqloppijsTx5JD7IO1ODI3RRm6oV6IJijcaeRN0Sbg9Ic06YjtKSAWzIe6hU+c+HgDnaLjATPHJNJrdnmxwbed+BCAVQqPec28v7BV4gxyX7gkDn0/WfZwei0YstCDN5oSlEhU2PDhgr188t442qLMfdQ5JwpEoQVaCRhwUSH7b0TY00bwAEIoonfbkVUwHR+JEvxAhUMN1w55hDVAUifqLnnThVPe0obFJBwHa9VBOhfo7BnV3eu5rEgdMsZEsiaME03I9rXA/HGkviRvx8lz3mnOPYlXa/ZIKgG5ereuggeVm8E4tFANFZOgzwyuVwhqkOLIBrA+Q5pJRo9mMyXQyad2dHSwe25bOa4WKOGl4YqiG8fJJTjq72ULJTtBtRpJCKEDM5pHI+ojWD6VVQBM4W0lDA0xOMXlKVKqhGxsVrj8eqJ40qAMCABkYCgA9Cw5g5GmCdJR8FQJKS4f7uUGoo14djeDsgpow4CARIJmg4cGwSVJnov76Ho5r0aVaQEh4s0fU0GJZtO/I/HJ2gw/OaJ64JJPLCEX6Ju/Pa7lxljNplACEZIUFGOnv/B5FFc0RnqtMooOUzTlFPhjVi65bLgthDpqY63Bjxvy5/JQPcBN6HeIBn4PCksRLSYwQoC71IS3wSho3zgSjQc51RGaG2CkhESbOiSYaEE5xcKhBQKCtCjEuBgnDVlB3FKZuZKghIBJq7Uj4+BAu7m/iMPrZyZTHTrkDcN+TNOYdeU8z24tG98ugqNJ1590fxn120JrG+MsHoLGBRiOXwlgmvw2+dykY2F/dnT12csLw2ZTA0/RAsi+RCvrzAY2L8TUJM2cQDSeQz9wfGlUkdqKHq/kOOtEbGMQt1h0FFc2nXA5d+hYZaedzDB6SksliyC6j10xWa0DJbxXNtLzt7jLQA8GLJ4JHR84VXp9mez7PYCov2TsNlM1sb39X6FQoxzU1Kesb7NL+w1i9o6VdMh3IEyHdA6KO319eWra9zW0xrWpq8NpI2dbBoa3h7YAUzikDzFqrPKO48mcbz1O8MY4PD/UarCEKgosXRsWkRM9VqK0wrFZDV4PAgtPDkUXTmYoMDj5NgU1EURwSeC8IGH4XxaCgwUdTzwdQgBUAF5yJlYK5Oo0zSdUkKDJgGzIAZMDCffMGsIyTk7Db0IDFC+PM6ppa7cnTZzoPWTsudQgCa9+q0hS+lZaWNmxReQiSYRiDzs4uWFtnJ1xEST8NX7hgMzMfVNTx2oAB2F/e7PYzjsY/zaa21jblIcRiN/J0GUGKGWL+cfZEa4Om7PLypt28gYnpgiQpbt2+Ze/fz+o67967Y09+fKKi/tLEJXv2/KnOItbFs2dPZSQ+NDQok0ukmSgm//Tnh3bxwrAQ2gxLhkeG9XM//PDELsnjoV7/DgKXGIXmOU3Qnb0dm50FGXhX7AeYSBOXxoTyJr7jAcKa4DODYqNRwP69ODam4RvnKc3J5eUlPRsWM+crDXoKVaG+U0mXdIDlJgaJqTBmiMH+IkcRMi3H/s+rKKdhq8GB8g9Yc1nJKfl5WXJ2mMATCWttarRb12/YG0lFZm3/6ETSGOwZqn1eU88BDzDOlRQDemcBRKSiyzV6nqiBrM4LlxLg7GKgd3yMKSwUfgpO1mTCSgXYhMQDzvWypauR9mEv462QkRk8zxFpK1CXDJvdZNGLXfYQ8Ua5YRj66p5QRBfYQwymg9dGkA9l/4m9FHyDnMnmTFoHjvggWDIW4b0c0ecxJ+Z+kjDAy03sQM9JfRDhbEc1CASawbPG826++Pl4lpAzcD3nclkMnYOkFecVnjlq9gN+ycPMIn4k7OaN67reg8M9O8kc671k/soAk4FgQCZyCrkclPt6ODjAmXtcAw0ZGrdejFe57GE6JZALwIPG5kaZTvNzNLJgwPB7MGdjrsA9I846ewl5nFo1iMQepREX2Ix8DxZERHA7yzqvNSz5B3x7qqqV1wIYWFtbkbExA1bAJDQOYQrBxsMsGlkcnhuSd8j3cT0MtcljBWwpl+3C8AU906bGFqsoV9hZJXvlyDa3NtX05Llmjg6F1J+4OGi//tWXlj3ekV79zKs31tTUYv1DF2xpadU2kBUq44fB8vP7WN+Aqa8zefDEoplFfCL3ZrgqD6LMsZgeSC021tdJLogBBdMTBvvkeEsrm16TNDTYi5ev7XDvQIP8vq5Oxdkbk1ft4fePraKqVvl1Q2Ot1dQyJFqyyko3TGefE0MwOQfMI98QS1g276yIgZELdloq2fFJTmtsZW3VByaZEw1QWBNcO2tRUkO5rNZu3BusEepK7jNrUvLCFejdO1OzMjTcxCriFOJe0YUUGcGbQC6V5n8nnnEWERdBe0sa9Rxk9LH4cQlYl4NlUGqFkjU31NrNyVE72t+3O3cwZE7am6n39ubdrBjPDU2NtrqGJG2DfD3eTr2z+/fu2MLigqEfH30FYVtk8zlbWFgS2549TdOP8+bSpcv6uYcPHys/cclNl1chFwfkRoxAtgb5LR/almxkeES56I9PnvgAVgb3ZTdqJlZJvtSZFjSlxX4ulez69evKZefm5/VZGbL0Dw7a9PS78Nohtxb7naabmy13drRJopC4sLG19VHKLrCb/Z4nfZhkpnPDwWDO8v+UgUw9ED1sNBNCYlTePV7DS+894aw9JG6o3WHyyBND5tMJq6tJWbKyrEEFgxgYE/QvMJcmX3329Knyu7t3b9vshw82PDKkfQ1Yrrmp2kaGum15cd4WF9bsF7/+mW2vLFtTfYMtzi9IZg2A5vjkFVv88EHPAo+wtZ0da+vv0zrr7+kVu42zY3V+1rqGB21tfdPaewasdIxk4p5qN5gCz56/lr/aaZlzzgGaXoy7/A5AHhD9NHIZ7nmp7nUJdRl74PjowDraWhS3kD0dGx206sSZTU5eEVPq4aO/SoKoIpmWxw2xg/UaexrEbPaBmyU7SyUap7NHqK3LkszxuA2rRMbaaa/LkZbk/wO249xnEI38JnGV3JwY3NHZqTxKHhb0f3T2uwSQS/y6ZC1ngDf7nfEqCe6kI9nTada7D0I5c8lPvEntUrrcHBj2nm86Mp5/OzrcV+5PXlfM5eWrVsjhWdJhB4e7trq67oj5ygrLZegvVVlXV6eGp+ub25KvvnHjmoA43b3dtrO9qfMIwAm5gfxyZOZMfeVSvfz/hsY6m19atnczc5bJUuMw6IeRCVOwUb5J1KsfPsxqz9FX46u6zuWMqVnkZZZKh3ys3iYmxu3d9JTyXvJi4ktVbbX2Fs+ffyN+IH8HaIC8jucHCAyWCPcTKa/Vzc1zrz/qFq2FMBT0Wt5BbYDo1IvDglC5mMuxsQ7dW6GsM4f7oHoQwGbsBch31YFI5IfksFyTBk0CpCLXiMyZM2T5Pc8ZqTc9p2JfM9Ry8K9LyuFhJbBGiGOsFUll4qFSX3/ex/L+m8cX5R9BepnBk4ZaYoqc6Fno2QFOkkSlDz24VtYnOSv5jHpl0RA89NAcHOPg05JgpBVar8TZyLxgfCpgSPD78PsaclX2uBRUXALNc8kKDYX4ApjnQ1x/bw0oYNEGL7SfBhWfNCl/+uvfxh2YaG4VspIvTfPKZ5rakpxQlHiQBVmUViEpZFM6JaQgXxxgXZ0dgeKNXAjMA+SO/GcJlmw2KJFxYqjme40fsFGeJDbUaAroQKTwFL3K6WIEpCi9AfJOzf9A7ZIeegJEPUbeAfEu4+1geBp042iKyIsDlK8kgxyJTMHMoUSiG5t9sdEfm62u4U3zBz18n+Sfo9XlU+CyT0oZggmUS1YxKHEqIsUuySCHjQJfdY0K70h7B23kevtpNz7M5c+HOtw7AjivR0BWIgfbVYV4LDK94ejX4H96Y9Q1+blPakoF+p3LGflwI6Kd9b1gyuUTAy8qXS8vHPSxGapC0v06CJoUJKf5jPV2dQgN+erFU0mBkSjyvPS5auuUbDPN39s/tEp8CDSICoh7mgjoewc9UibzrjGM8omvRQHxP9EKpnDmC4oy94kml5oBku0K0gmYJLa02ML8gtYvqJpcPqtnGpGNQhNSfASEMQg5X0MMptxoimSBJJjEUEMxCm7o1hrGOKl4K6gAACAASURBVKLeTTVBVbhfB8/em/+kmQw5uJcqgVzaKhxImKCmE5XSsC1g9neat/bWZiF/ARoxrCCBaG9tVfIlOSMJICYsXyzbyWlB7BTMtaW9XuEJDUlgTPZEH5TxZj6gDwIqKazRmMzFIZY00hnoySgPqSeXseKA5RocfRNl2hxVEWWMvDHMz3szgCRSTZNAF/ehJQguGE8uMaGCMzQKSBq4r1ESwumhUH4dfcqXxw2XrlLxI18EZ1lQmLFnZBBfiZ8NknTOSuAfYjIcaefRrI9iyOXNGM6xHjwJilra+uzFopIl9rIQFmi18jy41yT5xDCSCT6ukKvRrN4HhsQRDQc+kQ5iLSjhRrtUOpyu0ekyZaBa0cnEjMz3KP+JY6TGWEooHxrnrufr6801LB05GtlxNBxB2TCgEPIpyIEg+8QepvnLzzM4ovCUnrAaYmXtGz4zjQBHedF0c1YHSTzri33w0RfHJQNp0nOPuPlu3uaoFYoFJXsktDXQ292Mm+Efz6mttcOOjnKSl4BmT3EmeZBiXhJn3F+Z0IFuLcB4axLjBTaGEHzo4SfT56wSKNSsER/2OApNjCqkEEqn1tXRas1N9Vam0Elyd4t2Vi6KMk+TTD5DpwUNDPmMFEkM4mX0K+kyvCc8gQWN5c80Lw8dzgxQ6FLKPTuztbVVafKna9PW2tKkxldLQ5PMtkGF4ePAfenr7VHDJXdyLBQrA5XKqpQdZPO2uLFlBUtYvsB5CHE/4TJXlQmrrau2S5cmbGllRWaeywtLgX3kxR/oPsn/qbHpzRs1E7VufZCpBp70rSlCOdPdXA75JzUAZabYoAIMCRG0xSlwaW5RNLN20CpGF5hmWJRPZB2XyqeK6+wXMZR0PS4LoP1ZOpNEYF1dg7wPpmfnJW/FfqDoogne3d0huaCTowMNCOtqHdnnhtKOuIa9J2Ri8cyqJCHjEpNqRiJnIWS4yTDYm9lIRdToXjfWI+XEWe/nAv+1trV6k/3kSLR+7gPINCj2yCmtrKA3XqVmx8L8ooZlGA3/5S/f675PXp60v/74Vw3crk5esm+//bMMG0Gqfv/oRxsa7NeQ5dnT53qvto52+/D+vfSHuZ+Li4uS1iAezX6YFbsCJhXSS9xj1gwNSQaSkouA2l4DW9QBFvwezxt0cltbm3sZgGCuqXWmZYFcxdlOKpKJRwEQQnxjIEjDiv1MjhjlnVjnvJ48TUol+WfQyCYOworBE8PlLqv1PqwhmuVbW9vaOzS8WYMqLMsl++z+PXvy9LmADaBAc2Kxua56bGKA+1SIlTSZ55NRl9nzRm03R76JheaeQTznVCIdTHMZnHOWFcJZFmJ+YMAxqEB+i9eB1dXd3Xkui+TNU5dR84GeIwUjuCUiO2OOJY+Jc8aDSywoFgafKPIGzjZ+n/vqr+eIWmI8NygO192Xwu+ZBsjBZ4ZzKKL2/IxxdCHngw/k/NzWoIezIkgoENskvSnPLh92uDm855v8J6ZxoaC17mekn3/82/37n+lntncAVSRUCxD7nanl18q+qWto0O8y8OJ9YD9HRge/z3pVPAqAH/Yqci2SpUD24+RY5zhnG2tRTF+aVkn3NVlfX1cTktdA/okmdW09A2ze1yVkaBiiNU4OjM8ewCXJRkqCwVmZJGnOrnANdPL4ru5O297YVI6SIkxqGEPdVLR8IeevK31s9ynjvQCCcS7xujTl0OAmL6uvabDWpmYxBDG+ZQ1jfE1Ta3drU0jw8dEB++LzW7a1saTB9au/PrH29k4bmLhs0y9e297Bsb2ZWbP+nlZrbe9QbgqaPIIjkArd3N4W4/3uvfv2zTff2OVLlzQIwFtm8sqYnmnm5EifScbQlWYXRsckR8MeJ+7jpyCfnkSlXRgatCKNrqYGm3o/Z4WKlNhoDPyQN2KYnMnSTManx6VDGCTT6JL0aSXDb0cj0cZBZopGKesFoIoYs4VTeTrJL6ngDPYoMRuNrnmWn+4L1g3rDnAcA2kGEuSQyFgSj72BXVSTETan4pfY6meqUchbWZcADzQwEjDHwWj/BaMisIaFzg7ShV1tjXZLDLmn1trQYJPXx5hf2OLKhh0wiCmd6TnAKmOQxTAZj6C3b984qtmDm127dlXXCfsCho+D+fBSqrDJq5P6/29eT3lertw0oHQr3YMNibaLo6NiwbhnZFmyUeyTZ89fKL9k3yt/DQ1gnlH0sZM3YJmYU7Ib16/LqwCQg+STa2ttaGTIZt69D/I95A3uh8g+IBwBwOnp7pTUIGtne5emdZV7ShwfnwPOeB7sE64lMtAVOyPDNtS5nMehaLBUkBHSewWPNfLhRIohtj9/4hr5KXkptUmKnoX6eqd2/dplnT9//OP31tZaZzdv3tC5gHcLOdPk5GV7/fKV3bx1XdKLGxu7dvXyoN2+dcmeP3kipsNnP//ctj58cI+UrU2tc6QuL1+7aqsLCw4AyuZsfm3NOgf7xXbt6u62/eV1gfhSNVXW3N0lJlKpImn7a3t2cHCiWg5WFAxCjNKRRaO+lHy21BCQoEMCO6c9Lqlg9nqe+hOMvg+3+YLtxV4tlx1wNH5xxN6+fGE3bk5aT9+A/fHb7+wke2rlikprANBxWlKNQbzjnKAep4FOrtvd063nw7qjQUu+BgOYNUteTE6yuram9YSnB4BRSf/U1egsh03JOdTU2CxJvvmFRQ1FqGvT1dW2vLLkcTjUApwlMdcSoCz4JrB+iP+19bWKk3yvublVcpaRXeX9GYbjsIkbNQzx+lUTDq0f2DJ48mxv7QhEQ9rB5wcwiI8Mr/nyxQv1X2AeM1iBWSJvpXJZMTwvj8+ChsJDAz2SMGUNYCZOHkU+pvpAQFeeDcBUGudpa2pttc3tfZt6O62BH/KRgKn4zNwP7gugEc4MpPKIDzTgtaZlDO1nFAGU+3v79i3LZk/s8qUJsVI5UwulU8kNaZ/IYN3Bb6xV8hjOKIBKm5tb+vn2rm7D+n17Z08ygUiB8vr01KJyAOcooEB/PgmrSsEY8f8fp2nODig6uycqSsgvlljqvrEatqSIs4AMkGh08B17NQJoJZep88KHxT4ocEUPAUmDjyu1hdeU3OGPPT/fM96TEQM75EFRpkmgDAa15DKZqH7hvQrWbux78JrUbT5Y9SEKXRwHOADicR/TyP766Fnr1ykfNcAqUgtwMCDXLkkqeip6Ng7e1NA7yrSHQQX1EjGXGAkgxq/De40+XNcVWEdbp1iZ1ME/DSr+NnrzP32KT+7ASE29CkpJglCkl0oKziACReOr8cMGVBAHBUbFbC6CnKhSDQ062EhAkH+ggGHzc1CQIMnXoEiyvqZEQProQp05lYsNR9Ls+sDesIASGIur2IyMgxQhsWtq9NokfARuEAaSWslwgIMEpXjyIMJhQvCQ3n6FIyX5YuOD4tUUV1qHlQri0ezbI4CbZcfEiT/VgAzavXEgI/ZFyY2ynZrlen+gUgmgJBgY08rfAl3qWqQ7SNzNNjd3VARznwnwJJMUZgRPPgPXB8KJexO9O2Kx5ci6kEaHIlUFXkj0lF6HTmhEkUt3UubANNw8MXfPhWDc868YFRpUxOayJtdexKrxHSSZHO10qgDf2lRv1VVJGx7ol5H2b//pn6yxvlbFuXxDMLGavGpt7Z32+z/80Y5ozCKpEib3XJPLcXjSVZVKa33FwQuJdUTDx8KZNJnmjQ4G0f+z1tzaoj95JiB8aDyhBUuxNTo+pgRZhq+BiifNZBk9nemAZO3w3DxhCuZIYY3J3Bb7XQ0q3KhTuu7hfmgApwKNot+LVRVpgUnA2qAAqUY3NQv9sUaHFQluPpvhBYWcTlVW2jHavKDa6tI20N9j76EFYxbZ1KBrZ69UIM+QzQt1yupLV9WIZUGTjufHQcvz4fB3aqEPr6KkhIycNN/zRj9rjWa6PBFyOTUDHBHi1NbIXhAClCRF2rgubUbjkQKQBIRmJe/R1NKsNYncifRagymWD+VSavrCdlldcYNAZ6qwTt0cj6+oXcxapRCiEPVBg6dISKAhreDoWZofSDU0KdkmHlDA8zyIUXyx17hu1hZoLDXrgtYp3/emPr4ynuBFrUniXBvmzmq05fUszhGoQcZOknOnp158CrFRVOODdevoDEf1koiCbGFNOp35o8k5iSXPQs36ttZguAbV3wehznD6iPLm84D+xvAuonklZRUGvmJkIOMUGkEUb2JVgNZwVRI1d/iszS1oVuf0syRJFL/sodIZBvIMGPx+gfbiPSmUSOoJE3zm2EQEUUmciNqjzh4J9Flo3zL9drSP+wOcybSbzy6WjBLrGkmxrK9vE33kFQTKEHkRPAaIzuw7CvmY5GIOOj+/oCILlHxsuEevFtHQRSUPBpTJpIzNKe6IVRSTueyJmyueZqy1tVGF0djFi3pWUHAp3FjzNJJBW5HYPn70g7W2t+uZoyHNzymGq+kGldgbWMR7DPAwfOVzT828s8X5JUnk/ZtffW2bINyRpEihMZ+xgf4+6+vp0RAzhz/Nac4OcxmzdLV9WFq3qQ+L1tU7aIkEQwM0gSv1GjV1INWLXuRkTlWAsP7ZV0rEg8GmtGk1+EaL3w3wkqmKc6Q77JE4eJMxskzdEhpa6WysrLTlpQUrn51q8NTT12Otzc26V+5T5cgyNUhgfVVY0Hp3U8U4LHbt+ArFlIZGkGl1tri4bN99/72tr+/ZKdIeLQ02PDQo42jW06VLY/bm1Ruitd25c1lnZW9fl4YXoO22aLYRy/D94Fyh8aam+b7+3RFh7iMlGcVTNzpnjx7u71tne4do9EgJ8toUvHxuzuut7U0hx5HxmJ56p3MLI+m5uXk1ZB88eGBPn720dCph9+7dtoffPdTevXf/gX3//fd69hdGhuz9h3c6n4iXm+ubiulIdayvbWi4vn+0r3VDXFaBFND6oNa4ViSuaH4ycKHx7w0bN2eOyGNHlbsXE+uWNcvgjWfig2fXK6YQY6DLZ+QeUlxxv/GxAKnX3d2l+y52EHIKtbUaooyMjGqfr65s2OTVS5LUJK9kKMJ1wvahSMtkvfEG05H3wrulpbXV2QIMVYKkZarizNrk41K0dE2tLa1tqHhGy55GvvSrJbNA3C+5DIbYnz5ocoQaZ7APaFnzQjgG5pz0lCtp6vDv5EKZ0JRnq3LeJ+3gCHPtBuW8oN3xPdne2tXzBulI7svZilwG+SWFd5SuID4qP2BoRl4rhKA302nQ83eXGvTGkvJBDWCdNSrWnQyqvWnD+cj3VSgHuUXutyMW0+dnRRz0SzqjCgaBS7JEmRXP6atdojUgVnl/vx+e63EOxhyB1xBiOeSA7Bv5DjGsB4Ah0IprONJcoSmwt78jv4bevn6xIYgpAE5gXssjQOAJl3Xlerh/UR6E85R9eXSEdNGZpNJgwHLPl5dXtP77+3ptbnFWDVoYNZJZCkNnnvPY2Jiknzo62nUP2avHGXTeq3WfqT9Yl6B+WR9CKoZz1nXvK+SJ4PHtzA3DE8jeHVtrE1rkeTEpOK+Teo6Yu2fULOW+01DgdThv2Zc8P54Va4D7h+waecf2+raaZ2UrqbnMPiSGcNauLi3K72F0pNc+v3/LZj+8sSvjY/bmxUu7MHrR6ptabPbDgtDQz1++tv7BYTXYNja29e+DQ/0aGMIkQ6oEBshv/u439tvf/tYmxselz7+ztWuXJkatt6dbjJCd7S0NIGGV4dFSXVcvn5am5hZ78eK17WxtWXdXu/38yy9saX7e1lcBG51YqTJliaogKciwGvnaukZbX9uSrAw5O33C/CkDTFDYTHgSyk3QS6cZSy1Hjkd+BeeChgzAFge9AH6h2ePeUnFoFo1IBaJLI1EG4rRCA2AYG6rH8FGsouarEAJ5F2Nn9rf2G4wCZ+Cmk24IrCavBmUeYz5+/b+lnzQgQIpGspFnVsmZ39Fk//bXX9v76Tf2buq9JZJpG7owaJWpGkvX1NvM/KIkKfmsDKYXFubts88+k/wejAJAKpUVSZu8elk51dLKqhrSAKUiWxW2BWvkw4cPYnMrvxKALWG1DTXy7qGWmRgblw8Dco+c8/0Dg4oh09PTOueIt+wLl6YF6MPgwoeQcUBNTXjr1k2bn19U/ON+Nbc0ySgbTX32jn5W8koO5OKsa6yvV160u7OtuHtwsKfvsSc8D60N4CWkcRk48tzxQwOp7yhmxaRQo0Q5WcU2GvZC8bt/jlhKys+dBS9DdGrvAsMxR0DXVaWttiYl6aebN67qc/7+d99YXW3Krl67qljw+NH3GsgD7Hj86IkkGelxcD71drXaL7/+zN68eikgxoP797QXyBn3YVYFzykkpA739hz9Xyzby+l31jXYa5XptPUOXbDs2oYGGJlC1lL19TY6edUsWW2Hq9t2eJi1EwanCdiytfLjyp0WlLPQfIQBgARRXW3adndgXmVkul2Vdvng0zxDfPI8hgslsfPF5KepWmHW2d5qcx+mFaPHJi7ZP//+9xpEMhzp7O61XKGghj9Mnu6eXh9kpVJ67oAPABlw78nVYQ0g80i9RezlWaCwQQ7FUIPYto+vzP6e7inX5E1Z1+Dv7u7VOUyOgPcGZyzrYGtrxwYG+jXwiEoKeP9QPzG45M/FRcAqZTGnkfvjOlHruH37jnpN3373nYYo6vXUVFtvf498tIaHhqwO6T98GtS7KNjrN6/sh78+tVMAi3jc5As2NDJoFWeVtru9q/uBn6GY5p2dWo/kvusbm4rhPb3d8vqiNkAuls/xxedf2NDwsG1t4ulCA52mNKAb95EgDsNoGRm9aK0okRwc2sLisljQGuSdZKy/vz8wyE6DHHnJnrx4blNvpwIzr2wtzYB+AljvNK8B+e3bN3VdUl0oF1Qj8XfyI9r4nGHqu0kNpGSN9T6QevLkic0vLeoeXLlyVfuPvtRJNiupQo+HZwL8wJgjVxUwpAQotOheFin3WPPz1c2xxZCKnhL4z+KpqHq/3iVyz428uaaYAzkTQmAL+AiSnfIaj30LMI58hpyK2CWPSIFSXa5O+Qq9rODPQRwh/jvYLqHzNjIl1XvMZsReiOBH9UFDTRAZqMQYB2VgZl8Q81uDL9dHCUBezxO4r8qlg6qDBgqpjx4qXA9xy8GpLqVMDu/AEAeLEcwiyDmqEfAMJJccfFLotalHWirp/jPcAqArtuhP0k+fnNs//fVv4g5cam4NVDxHCbMZerq7FSw4qDG5ZffQ8EOT2mU1drzxGWhJND9ArnJ4qBAJxso0zWhW0dQB7e6FdF3QtK1RsSSTnQrT313uxaeEkYqtAy5IMNG4igkMQYTAoECDiVOKog8JIDausx30eaC8y8THlTkoKghoHJjSEVezPqkkUSa3XE+gB0Y2Ak3cKEclCqQMkl2ayE2pXVIgIsPVdBMD302Iy8GckEKXhk9dTa0MPblWDhuaMkLwpLiOnA9OJH2ENntOTR1v1Hsyfa4tDKJOzTY3L5esR5B6ifctBsYYWGleiCIaEnUdJmgzh+ZxlC+JPhUgXD9N2OOz5fei9jMHhmsBpq1czAqd3NXZandu3lRisQTKhOLzOKOmBAnLnfv3bWFh2Va3tyxV7YhrNYiDt4HkrkBEavASKKA0ugL6kEXC50XPOsoWcIhxP6Ch1zc1ng9kkFPi3yRT1tmp+856jKyH2LyIgzm0ayVZFMzEKEZocvvgxxvF0lSGXhwOizMZwDkN2gcmVUr6WCP+LLywJ5mDbolOM5IgQt4FVoUa8tAgQaDSEKtGLx9TPPSKTU06mgQ00PjcaA2zx1JVNVaZSstUe+/oxDK5U8sXHLkmyQYovkHCyQdkLskQ1wh/RiYJQzJRCWUc7s0o0eHVgHbElOQjYjMoRXGSUtLKgUsM4HNGqiTIkuwpBvJmnZ2YOOcVD6KECgmjo+IcOUOy6oMhl6OJjQU3Iyfpo7kYUagu9eE+Gz4YgsrrUmA0VwLTQoZXTiGV/FCgmrphsOvwE3/0vAOVk991ZK7oO0pHSKApEqGI+x73wZ3HDxBceHJYMBDm+eblFyLmVWA2cY2scT4b94p9H314uGaxDjRcdMos1yUvH5naMfj0JEnSUBqCOZLWUXKe4JEk8bNi/zCkVdIIM8Bporwv0ko0eWTwhjG0KMAlDUWcgeL6mIoPwbsF6THpYVqlitw4GPamoD8T5BK0xoSo8eEBhTNxms8d45OaDUoQnT3G+UFjnWsoFpGSYX/XKoG3s6RkLqwSn4NdNVlpxpahBn+i4U7c5L0pnlh37rPkyZsGZHr+iYD0CUhs4qrYWe4nBPUb6SJ4zZwbucyR1dPwl9xAUo0zYjDsEVgbyI3s7jNsblShRGMK9Bs6/JyXPC8a9kj2SP+3XNKZCBKPe40UUhbUaD5vi+9n7eTwQE3+9rYma21rkYcFzTBkMBpra4RkTdfV2Fmi0jb2Dm37MGuZUzPdJpgVuYIGeRsbq3aSxUQ6K/3ZBky6HXqte8CwTVrRyCIEvXw1UysrJJvU2OSIep37jS0qsDR0bPShIwUry5TBDE2Pw8NdsRkoUtnf2lewXwQ8SIWh0Ec2FkgoYpdQay2tdnh4HCT7XF4KVsLzly90lhfLNMQZ1CPvlJJ/wvramq2ubtq1q5ckyXBwmLGbNybERkEayw1+W+zo8ESosTSyWMmkCq++/n4ZItIQ5DwhJrNXTws5NbcZ2InZmYEh0CI5JBgxDB9S1WkNEVhbmD8zcELuhcZe5iSrtcez58v9pbyIi5KTvD7nDk+LIhz0LpJJNGZ1DiRpcNbahQuj9vTpM98/DUih+OtIZmpzU+uRNbW4sKj40dnZJXYOOswMsWfn5mxkZFjXgZk2hTYxApQt0k/EChC9yPUQg6am39mVK5dVCK6trdvlS5clGYE++Vdffmk//PUHnT0XLgxL0oN9xn+sld2dPQO5TV7Es8c4nc/I3zlP2HcDaPG/nXYz0rJ7AxHricV1DegUH3tTI5uVF0bCyra5vmYdXT1iCC6vrrsJZ5DucWBF0K0OJtSc22IyFNnvICXdmys2tMSmpemHzCRNtXSNZbIMmsmraKB5wUjMqKpyvzIKZYpzyYIx4NqDudOm+8/PtrS0CTlM7CE2SpYiILEjEzDmaLFwj+eQfNdC4erxE2awn9nOPHHJC36f6+X+xsatcuLzPmoA1ahwT0n6KTIVIlrRDSWRCPL9yN7mZ3ldFdXkWOFMiyw/B6SkFfe49k+Zp2V80mgQBKNLP2ud0UYcZ696/u2eEzwHycrAIj4tBMbFiSM+QTyLbWdq5BOPWJP8m3yrAsOXoTjxk8EXA21ihxrfAUnMzzp6kjO4RTGDnISzBY+T/UP0152Vy55F3kPofYZZDPaQKJSvkd8LsUGlP32mHEzefcjW8WnOSsrrmxsbJKUHTJXhGxIoNF0Z0rV3dKqB5IjflAoQ2EN8XtUOubzVVnF9WTWAOde4vlM+V+FUciJIP/3m11/a8vKcdTY32tPHf7Wx8Qlr7+23uQ/ztrK6YY0tbZbLAbhiYEWs9SYRjZ3N3T2bX1hQXXH9xk179OiR9hdDyM2tHbt6eczqa2uFyJVsa5KhC8yQJns9Na3hR1tHp715+8ZyJ7DITu0XX9yxpro6O9jbtUc/vLTG1harq69WbCR/mV9aU5M+mYIxHrTFYT5Vel6REmO0KMYD8k9IWrEmqOOIdWocBukxr/ecFSYw0Wlezyw2nojzILYZPHDWEmdpdlcm3QdQfjjIjUou1T2rGIa6rGGKuWZgvXuzjC/lDbDPA5DB96h/LwK/YkEJ+Ihc/axYss6Wevv3/+43VpOqsI2NDXv18pVV1dTb6saedfX12THDh6UVoZ5Zy3PzC/bgwWc2M/NOa09a+mby2KIxNT+/LK8Q3ps9RMy7fOWy4tLz5y90Vql+UH6JzFzOklVJ+UQAqpiemnb2QmWlDfQP6tm8//DBZRND3U2+dZ67BfkmDe+Va1banTt3NBSRXE+xYM2tzdbX2yvjXwAQ3Mc4bCWGIAGJ31RzM+fUhtY9uZ9AZbWYtTcqLrAPyBWIQzwTeV3xepJP/gjY0b0P2kdR1o7zTqjyMLgSExuT5SqY1twvpP0YTCTlCUlN0FBXZYX8sV29ekmf69s/P7aW5jq7du2aehrffvOd9v2dO9clpwhzZXVlTc9xoKfd/u3f/Uy+D8gy3/3snq3Pz1tTY72tr66BorKW5nobGr9oWwuLftYXCrYCe6a1WfUZedPu8qo11tXaYebETgEvpqps8uoN21jesp2dA0tV1Un6aXZxxTK5gp1JdqkkGbxS6dTu3L5u9+/ftnIxL1kqZMTwfDg9LYm9y5mVZXgBYxH5MnwS0/Q43Hh6c31D62fy2lX7lz9+Y4sr65Zn3Xb3WLoaSaMNDTeHh4fUl+CzoQKB9CS5jySZQs8HgBUN25gHKJ9X7u6yhp/dv6ua4vH3sEidCcifyVSVJK8kS4QPUEO9BojkTfSanj57Zm/fTikew3gl7+L77AnWDpKZ0zMf7PjoUD0D9j31CmsJ7zD2FeARZO0Y/mGUjCTdzRs3bKC313IwBcpnknqVvGM+b3MLc7Z/dCDpSCQqs8c5DeLYF5FdqCFbZPqpl4znRZ3WFzmc9x4q5KnDoBypNYYJxFLWCVJc1JHcT0mfBmNpgEX0rbi/MCbIubiXMHOpN+XxgKIJPZLTgs28f6/BIbmV+3+5twwxjb1OjT08Mqh7cVZR1l5kyBMH6uTj9FTYU3mxySrkaUT8QdZwdn5B50ZTc6tiOPUMHig08wEbM3DnbEd+OpWqVk4dpSwjo5S+lXtFuBQ294qBCLkEANyorBLZmlHhQ/VhABBrSInXiEA05FrOAmedEy9ivcq/k6sD/hKTPLDBYs4H6KOemi2AA3UGBG9Oah1nRrtfI4Aql6NDGcQVAOJQXCBP9RYAk7rqQexFRsZp7DF4THXgtxjFSY+nyuNCbewMW2ezO5MC4QV8HwAAIABJREFUoDT3ypGXYvoH4Djvo7wyyGarDxNiIkMZ5TBFzlJq6LqfBhV+VP/09bd0By61ttvG+roP8gLVEokBmlcEleq0N2n8QKJobnDDvGNvurC5mADz/2lekHCQCAlVTGIDsjKXVbOAjUow4oBg+kwSKcNZFT2RzvZJVvivbjTJCUGboCH2hVBqID/TQaUIU2QvNCPC2/NL1x4lEAWmvJoiQrAEIxwSJkdSuu4lwYwCB1QGQVfFWzAR5jXVHA/SAi6N9LFB5wMXzkMmyooyarzSyOJ9aHZxD2QWDPW1gDZo3hvY2cw5ylnBMvhCEOh5Dt5cjsbXnllrEhtQ4PwZUZSu7+h054ikJ7C54ZPLtYjBEv4ek0INi6QFyBDjU6Mgb16e09yC/BKfXSwCPnMxK+QvveGBvl6hMafevBGyjtciUcGwtKOrW9JXhzR/0H8OhuFcOwePKHoEatDoMr9yJg1INw5nDXSCMTjIAArcOCigAKLpAJUVNEjm+Fg/D5uHBuanhyj33RtHEZEjsV+hwGIzJHoceAHvVET+c5kS0Ak015xRoOeh++LFvctIMdV3A1+ts1rXP3YvB0/+2C8USnxeksoqDrTiqbWgHYwpVe6EMZVQnSQ+6OBy4PP+IHCLSMNIIuPEjtEMr0iqsRMlh3hmPOe4FqKGo4ZsIcnUZwkSEhoSIS/EoRsQll4IwuKgCGSQ5EyGQt4NyrQGQU6l0yrUhc6WbrgjJNHopUCneAf1QkLEa9Cs5jVJLrkeFU4BQadmUSimeE5RN5u9S7IL8oZnIskMiq8w5FTSiFaoDC+9qaRGVcllhuIwgOdT10BjBImoMCj1ilT3y5MqHxJKIoFBTmAZxcTDZeg8xvAe7inhzCtfV+xZp3ySEGpYm3MDUprXkdkShyNRokWkzjNYDXVC2hQKNEQcxRG11iPThPcGSUgB48Zh0eDeWTKiidKQSafUxBFzJyRL55JlZ6DQ0mp80kQhMYORxn3kvd24iyaey3lIcoO1E4zUXaseRIwjW2pr64NpqbOKomyIf96yEkKuW8/x+ERNg3QV+5+hUUmSPzvbe5ZK19j87JIKMRBNUJSRflKREjoIscnGmqOBSzxwFlFJrJXIBNOglXWrM8oHbxgHkswzgOju6pDpoRtON9pZmcGuoxKJfVwriT7v4w3+kiSDSHhBUu3ubUvqiNjNNdBEw0BODcEzBvJZGc0y7Gc90ODN5ouS8qksl21tccn2d/a0bvv6OqW5XFdTbd1dnZYiQYf5USpYNQbH72dtY/fIGlu7bHPn0IoFjGmrneGwsmgpZAKQs1Ez0L0XiJkkwcRCzmpiHHqsq2sbVt/gSEfYGEPDAwIdHB0c2PDgsPZvc2OTDDmJdawZ5JiQE1leXrSaamSATmx7a0sm4dDuPzYifO1HpKYG9Gi9asBGHEkoPi+vrOk11zZ2gsEez8dZQXwOw+epsd5GRy/a2uqa5Kxu3rxq87MfZOL89c8+s1evXllbe7OeUVtbhwYgK6vr2hvQ9clDYLvMLSxYb3eXkKsAB46ODxxtVgn6Eumzkh3tH4lBAHqwq6NTe2/i8oQ+B00CZGXYqxTgIF/JFYjjNJtBVCbT3jyjcKZxw8CKNYnJLM1JYhmSAodHoBVPNcDq7urVtYLmxoB+bh75j6zNzs4qhjEkefvmrd4T9Nz83LxeG4Tuy1dvJU3DGkaLHGYRhTvsDQp9msSvX7+yC6Oj2ncvnr+1O3evqzH3/v2M3b17Tw0pkOt3bt+TVjfn460bN+zV61eKHcNDA2rG4q9BGKXI29zY1DUTqze3dq2np1PSVRTdMZ/q7x+0qekZ5W+gtNUATzH4zck40tFxsF5ydvnyJcuduE/TISyK+kZbWlnTOqZAlgSQgBZFl77DP0wIO4o7B594QRpABZUwZdzUm0Eqv0/TmVyRNZtKnMnoN58D9e65HmuS3IwcFlkz7jfxDSkVzi+dbWL9nblet8AazoYl1tCg4H7hCRaLSv95PFEwvOXc92G32Begu4MWuDcOXZIx+lPEhkk8x7xwBXvuRpexqNbPxbyD84NcSF4UPqCBjcZ1ycNCyakbYLr2tQ8tNORAjxn0YDCc1tA9MByVRwRpQpeFcAnV+NkYlpHj0Nznuvg+TWZHRCNTgsYzw2bX6I7NUuIpf+ceSgouyO7w/8njWCuS1Uw7u0HDxFxen08yQxUJNbt4D+IECFaXnipboWx2ksPDwFGkcZgP08MHQrAwPVd23WrQwzVqqLK/lpdWZLpLrockHOuOZhdshLPAKGbwBfuUWog99fUvf2Ed7R1uzJz0NfHtd99qzfkaqxA7hJgLq5OcRmhzABCJhL149qNNjA3ZV5/fsUSqbPnMiaSfurq6rXtgyFaWVm11Y0uglLa2Tknb8R5b27ta/8S27t5e+T4cHB7bjRs37OXLl/K6Yc8W8lmx9Xq6u+wvDx+qsUYeXlNTZaNjY/bqzZQ1tbRq4PLixQsBNM6KZzZ+cUiNWFjT3337veIdEngt7W3W2d1tz15N6bwpGzloUg0vBn3sV8BblUKYer4olDWo2E/kZ5EFVI4Aw1ksbva0N+U8v3aQg+PW3PCXcx6WiHu8VGn4BHMDJh/DK3IWeeGUykI0cx7RCD06cTPgijNqRmdUUCOwF/kZ1qxqx8Cu8JwYYBh5VUrDKuqeCs6b5nq7e53YdWCff/7A1ra27c3Lt7a4vCVwQbKqRucbeR+x/sPsrH3x+ed6JooNoX64cvmy7R0c2MLiiu6PZIOVayBddF1n4xudAfgoRobtmRXKDNp8UHHx4phNTU0FKTuzifEJrfu5+VnFNQcd4fGIhr77Ukn6K+RFktFKJOzmzZsaeuNvRAxpamm0nt5eNXIBQqlODEazxJ6qVEoD+A4Q/HOz+qw8I/lTBlAJDUekoxnkc008B+oF4o0Q07o+ByYpfz4HGJ26FHTQu/d827/PoAJAIeUWcV2ebYYPEesob23NaM6f2N07NxSPv/mGQUW13bhxU/XKD4/x/EjbjevX7OHDv9idO7dtfn5e5+HYhX772YPb9u2f/2S506J9hfTTyrJ1trXZ+tqqy/rkMnb9zm1bX5iX1BiN9D2k75D0bGgSu3NnYUmAriL/g7Fd32AXRydsZ2vf9veOrKa2yTa2d+yvT15YZbpazCQGbijdHx9lrb+vzb784o4N9XdbVUODnWZOhOaHRXV4xKCRBjGNT2ev8HA4U9krwJfEbhPDNWUz7z/Y7v6BmKaWSFpza5vWPNJG5/c+oNwjk1To8DAMVE8kIMLV+0AlAFnS4EnHToWNWk3+Wud5JeuM+PRu5oOe8RmDppTLMJPndrS3yZuNtTk/N6c8gx4U59zk5KRdvTopFvXh4YHiMmwX6rGjw2PFANYs/4ZnCDGb6xJYR5J2CQEAAVGqp4CRc2Oj2JKqL5E1T7i/T2b/2L5/+BfFD8kXixnpfRWdQcE/k3MsShC5zKTX//KQhPnX3ydJKMBPDXWcUQk7PNjTWk2kWN/O3izjU6TzoNLNrwN4L4IlJZ1XXavroXbk5xiiIbfFEJE8XjUweagAhCaJ7a7uVknA8d7IFsKiV23D6VdytqLkpxlchryFfbO/f2irq2u2ubktWWn5btTV2cbWpmoCvg6R6ctkNajQ8B+DcPpJACjkU+mMTnImhs+uyoCvBOoS7kulfMwxFmGQ7MomLpdJL89zgDiQVH1Zdh8Ml+CmV8cQJGftba3yzpWEUohh5M0wY2F4uS+Xy0xGuXOGDbAfYY5w9hODI1NL1wYTMvhoALLQQAXVhuDxxWeIXrYOTvG+QuyjUgtwr6kDHMTizFQH+HruF3uH8ZxRTcpAQyovLt0cVV4igJCYLzar6nGYndGrqKSB1k+Min/VOP7p//7//w5cbGgW2pxNFxvc0IiY2MpUpqFBwwg8Jtpa2mSmTbBCt5JJHkEDT4utrU0FNBJDDjoOJA4+kH4EEn+PpH5eibkYDpUqZkTf1CZ25LPMisPE8NM77Aeio4NjUKF5TSPu5PhIv4dMhQ4LNGdpTCohJni4rl00Y2IowUFFsIvSSqDsSWgjDcwHAK7VGwu6iDbT94JRW2QjuIQFZju0ZykEo+YecNeytZIsBfNe0MJo/JNUczCoUKewqqsNk/IKKxUc1R8R7aBLGxvQl+b1z3QYRnaEdHyhf+E9EJrm3C81W8OfOpAD9T1OiAnaGlAENI0zAvzAVfAMCaN/xo8SAQrYAZ0rQ2ZJ53AQFq2pvlZFHjTYK1cuqUH55vVrlwiQXFGNGoxoT5MkneRzmpqTlhKAVRxjhgTaFQRq2hOE3r4+rcnD4yMfMJXR266z2mo3+IySUKCFMImj6BPKXLQ6mlxNasjQyAQxBloUOuOn4wdvdnijgCatmDiamrgkgjMKfDDDISiWi+jTrDV+xwsLkkVR04WKcT8DPkcswH3SDkrS5XcoeGT4B1NHdMaSpGAKpzl9RlDdlVa048MjJd31aAJTaB0dq9FT39xiB8cZ2z08tpr6Rjs8Zurvpq+SdQheJhy8kjQLOtUUDVFXW54MMtKV84WuiwYDA0hooRp8pWDGHKuoo1kQNa3dU6SoZ03hx3sTMyRRJFYJCJkq/T5NNVCHJCxIe1HUk3yC0KcxJjQbzeNPzNNVkMjjwwcGNLswQNO1aM+5XJC8TISWS4hiKtPbT+TQolRN1EB1uRs+c1FJohAsAXGqpmPQwpRsEhIYmKupIe/JBmvBpaVcD5TdxOdnACtZMDG0XNvS0b2OxuF6aQwouQqCzSBI3HPGB5yscV63oxOfhmMh9XmOEX0Rdb01IJIXAKgb1/2MTAuuUUNRDSSTalS5BjQUVhpxRSVp7qUCeth1YFmPopQHvyFJ6EG5rm9QY44EWyyUEB+5T87cQG4ByjKyPhQDTfoMrHcSRp/3oq3aoHXGs5ZkFSgV9GITlZbJHInOKwZJBQ3wU9vY2FGspAg4PDmwdNqNdRmSqHkXhjCs0YGBQTWLGKgTN1jjnG88KwxDKfRpYHFdYhwFrx4KKjRsYTQcIf2hoqCkRiWFJ8MKlzc8VjHOPQSBRkOYhrIHUgbBGetoa1dcOD46UUMduQ2Q+a1tzedyZNKY56zMl6ypodF6u7qstbFJzA4ayguLi9bV3aYhxtjIiIYGuCzW1NdYU0e7PX763E6gXp8y9OQ8gHqdtoO9fSuVC3Z0cmhNLU3SQJ95P2udNNsxd93atp6ebltZXtF5CgqaBv7F8Ys627d3+D4NtjPJGlwcHZOx9N7OjgpjEPmcC8srKzLWpMAk9mNozlml100mbPTCqGJEZAFxtnKPOUvqGxuZckpPfvrde1tcXpG5IGtCzMu6eg3t2Tc0zojhyHPwWrAAeA/OAgY4sCsYMo6Pjeqc7e7pUpOkr7dfDbqXr16pkc7hjwQcaDVphSOnmARZ77KQUSrJTYZLut8MWxy9XqH7hA7//PycLa2u2MrysmIz/y4Zo7096+8fkvY9n4v7hPwFDTQkJlZXVjWQuzh60RaXFhQDKb4pOHd3D+zv//7fWN/gkGIAP4d2+8nBgS2vLNt//k//SdeNBM7rV681KAK59/zZSzWFhoaH7IfHP9iQDLfb7dHjxxqcYWb53XcPbXx8XE2jH398JlQp9/nlqxm7f++6hlCv3szaZ/euy2uD6/z5z7+26Xczam4gdQHSEUm4sYsjanKyT3kWDKS+/e4v8tfg3Fta3pAOOIAWJLO2t7a15/lcU2/fCfVNcUdcJgeiSSUNazVqPWfEtDJ3fGytzU22ubNrDU0tMnukSSQvArFROWuLGuIxnGW4ynlCnCb3IzYgv8h7Dw4MqDEWQSA06BicMAxfWl604aE++/nPv7Q/f/NnFehIBbjPjBerpTP3h1Ajp+BePMQbkNGg8slVXGM4ce69Rs7LtUiOpFgM8nfuSUGjWmjNwGpUMy74n+h9Q0x1KVbPsyQVoFzNczOXW+Io9z+dveGFNuhuIfMwZZTcgt+b+BWHC56/kZP7+aCcMjAL/LXdY4aYERuXjoD2IQnXzHkCkzaebXwuQEjoY5OL07iinnB/CZd+kTyXPgumm4dCympwwBAPje3ymWRB4j3k7ANxG9kRvMfW9rZiuPKagBDl/EZznDyMPeEa0u5rkUhV29LqutaKZCFO8zY2Nm6v37zR+bq/d+hyaxvrOpsxV2cIgdExr8v5RGOVe8E5DHuSQQjyZMQcMRxTDDbwSStrrcFQwjSZhgjPkvXOgJLX495zXmdyWfv+EU0xagU3BJfGfS5v3z/8s924fsluXJuww71N6+nusOlXb2x4eMTq6pFf2bDltQ1LpKqsu6dP/lSLSyu2sLCm61rZ2Lavv/5Ksix41ly7fkMyH6Ojo2qw7u1sq5EFoGhpaUFoYBm1phkOV9kJjLuwF148fyX5Gcy///0//Fe2t7Vlcx/e29HBkWIzgBU8o5DX2jvKmiWrbHvn0Gprm4TGhblZOiPXLss8mzjgwB08+9ygNDZ4gvrFubdbU2OTUN54XzhMA0CMs5754rmxT9ZWV1zqrYqcEnacn/k0pxjSKh9DmkPxnDWIdIazeavS3gBnrzKocNaqA+HULpcRmzflVR9peCE0muo8PHVgVNy5ftkeP35uI/2t9sVXP7O3Ux9sc2ffNvHMSiS1rpFWvn37tuRq2W9LyyuKwZw15FuSd8rnbebDnK7R6wkkzKp1jiDDg3+Co26dNQaKmUGF5qtlkzwT5xR5NOynkQsXdEYtLS17EwzZKgHwPKZEFQHPR5y1wvO5dfOWBirkBdwPfFJggcLSQ/qT5yiUPX9yRqeSYooSu2k20y9gAEytTV5M7KfOZgAgiWkAjkiMHQNazDo4puzguwjA8/vvfn6SPoVZjW+hAC/u5+MNTbOqaq7DDWf5+RSsE9hOddVm5VO7cf2K7hvrmXuArj/N3+//8r3y3atXr+jvt27fspmZGeVv46P99vnda/btt99YNluyr3/5wFYAOvR02urykgbqZ8WiXb5zy+ZfvrSWlmbLkvdlM1bb0mKNzS1Wk0zb8c6upSoqbW1rw86qqzRsGBu7ZPvbyH5RQyZteX3zfFAh+TKxFNyQubW5xtpb8UTotkuXxiUdyqAhc3Qi9k0mj3xXveIX5x9gCXJMaj7WFn2O/cNDSSW1tHWIVcM+57/N7S2tNcCV+LdQl3CCRGUDSUkG+Rkxz6g3qqo0TGDvcg/ZO9RxgH7wYsseHVPuy08M7xpy3D1JSLknEzX4qfT7kdOsVW7129/+k5jImLgfMJDY3HKz7QBkldx1hUlGkPyPM5znTw3Je6iWQdYMj898TvJMntcnLRmMlslfZqamlfuOTYzbwNCgGOKHJ4Bt62z69Vv75k9/Cn0cX2te84QhaQlwHWwm4gfDPkAp+LcFNDyAr6oa7fW6mirraGsVIxrQZg0/lzhTLIyMjUQireY+ta36DopRHhcji7Kpuc2BveRIpwXFN3IoQCXkjzFXqK11jysk7dLVCbt/9471dHWLUSGuPT0J7gNSSoHxrr2kIaLnneR1DK6Q5VtaXpaXBvU/wyJiArkU+fPh8YnOcSQ0YRqx7+hzuGxlUs/WzbW9J0JNyD5HXYPciP2uui0AMpQXBINsemlIJikXCsxMsTLzBVcZUI7uYA4AQ8Sc7R1qxLSmldTA0dPB5d69PnWQsftgqRcG8whVCvkyutKE9+9c3SMyTx1gyLCowjLHzgpxT0JADj50/zhYRerWe0extyRQXRxO0PsKCiLEXh/EMphwVqr7qX1UMnFvWAfWMTCR7yr1ShieOJAc6dG8Bkc/DSo+7Rr/9Pe/iTtwqaVNRTW7xAPGmbWDQudQ29/XRmSDK1Gvq9NhTrKJQZxv/AobHBwQRdJNWjFj9GKGLzX4yiV9n4YRDR6SmqjvLhS0pqcuJeTIGgLUf/nlEiQu6cLfGaLwBRKJIlL95EqXHSHwx2SMQsIHIz6oCHmPAihNEQ68yBiJXhkcFjRWNXARut5B2Cr4eH81HR2NLokUtIXDNFTBFt3SIJPjohxmdfVo2Ll5Nj8Lq+PkBBRVjeVO82pgCTlDEV4EgYwpExT4pJqumKK2cLhL2981+mIBSYDjfhBk+Tf+zuuA4lQg08DCm5YqEGIgVf5Nk8snuDFIO2rFp8NK1TWk8EZRnB77UMqb95pWc3gbTeaSkFrZkyNN7ievXNKgCnM4/BPOVAA76mmXw7fgciU8fxpbbtIUzW4dncCbIEm2ur6mZ01iQe3ANTB4ANlIQuba3I4i5pCUjndVWj4rNLVBsKOfShNcDYPzA6TSEQE0LpERUvPYG1QgwWSuGOR7XFJCq8gPYXlaePPAZZFcMoikQybBFLoyZK2whgbQlAxhvOkspH2QIyLBBMmLhibJHvstmahQ4zKdrrTe7k5JvyAPA9MCM0N+FzkTTLTrG1tsZWPLahubpG+aTLrXC/uUgkCJQUCEeQLhVlWsSf5OsumSGGmhINQYkKE70i5HSppYS6xX7ifNpYMjZ7hQXSih0F4oCU3COkH+inscafvs92iwqn0emyvlsm1sbOp5OVrWC3mKSkc6u+m4mlGg2mGk5PNKyiRlVPLEjs8ldEeQQ+NaPG58lNlweTnXhIwDQiG8pRGOFIxTKfUaZ6zJnAod1oXT2F1qLcojRaSfkKHQzJHnOnB0hw/4nPIpwy/0NdGKD4a9rsnt7Bu+eA9J5pR8gMBXlMTTa2D2FczH4pDSUbYuOSLjX9FLHZkah4m8fpT3wJiU5nyUxopsM4r5qFkMshJza5IovmjsoF9NXEW2jOd/AgslSFthKE1zmqYXz0vyJaUz7VMaNaCvSLI0qA4+JhpQhwGdDNShXedzkqUCEeumZrUy0S4UyhrIkYglU6B+9qQfGxsOXCP7RpJajeiP7yjGYbwH6pYPS3ziuXEdPGMliRjYQUk+OtZnYm21NDap4KJpg1cDgUbyJ4oNSRVexHaeC81/UFs00rjvx8cHGpq73AmDd4+NS4vL+jea2hROxAJvYhYsc5LT+qyrrrX25hYbvXBB33v6/Jm9nZq2fK5oP/vyvlWUyvJxaWlvtWR1lc0vr1i2UBIjg+EkNRz7Vw3CXEaJe0Nzg86xxcUF6+7scrTyaUENtJWVZcWwgcEBe/r8ufYsDYXdvR1pOTOcobjd3dpTY477w1AYzeT1jQ2r5f/rvHIGG8+YNYlkJI1z4h9mzwdHWevrabfbd+7oNdj/6PzSCBc9/5TiE8ZhvZo5FKaxaRqLC+IhA3AG9eQQ7Gv5qLB+KjAe77BshrMjqbhOsxukL142bggLjd5zEwpy9gkIN9a+73fXCM6f5nSPeE5nRZBsGHMihzBsY+PjolYzFGHA/PTJE/vDH7+zzx/cVvH/fmZRXhQ0oGDMPPj8gRpKyHx9/cuf24f3H+xg/8A+u39fg3ti6pdffW7PXzwT6OEf/tv/WjJbFFgaGlbXqqmDJMM3f/zO2jtabHT0gr188VKx98b1G/aX73+wvp4uNfIePXqsRhL5GFrNNLxgx/7ud7+TxAWF1eMfntud21d1354/n7IHn9/W2fDmzZR9+eXnatTz3y9/8St78/qNnu3dO7ftT9/8Sedsf1+3BjIaRotZVyW09fjEJVtdXVFj58rVqxo+sO7JIWnwVtXW2evXb9XYImbQWKNZxV6kAJTcoOQWQd/WCv2YRUaqo1PIT5qmmNFKjofvZTKSRXSGinuKKJ5J6s4ldDxVq9Q9ezfzzj0hhDAtac0TFxaX5m1ifNT+h//xv7fHDx/aH/7wL1YqgE6k0XGqddna3qLGDfF4G83y7m7lVkJqS8JqS/Eb6QYKdTEk4sCtvk5o5FgIM8mO+SvDAcnfERNl7siZ482Q2MSQHEzIdyPIIRbEAvDBqRBj19luys2CbIByRHkJnZ57PXk+jvcUzA+XNuAuiTGiRhSIxepw9rgGMq+nhkSQgCTWci7QDFCxLAmFjBofPDv+g2WGtwH5Gecdw2FdDzloYLASH2gKw1wjtyDH5XzlC4YaQ0C+z5qACeEIQ4ZQ/nkYkhDjaZjB7iMn52wBXYtWPihLZDaUPyL7trVjRweHWo+sQc5aZNRozOFTQTMXOT8+P/G/raVZe08eSsFvjz1LTkZO1N7WIrAEXhKOhDVbXFpWw4dcmToKeTl8a8hn41lHvDnY3xciH9m3mQ8zYlUxuITZSUOP3PbVixd2dfKCff3VfVtfWxBA5cWTZ3Zl8po1dXbZy6cv5L3BAK+6GnlIs/WNLZ07xFmKnZb2Dg3Ruf/37t23P3/zjXTqDw/2bWFxze7dviqWHrGQGIhXBWuOXHl1fdNa2toFLmI4yrkHe3ZksNeG+/tte3PD5mbmbWJsUOtwD9lfpI42d8xSNHWqDIA8cZjmHPJS5AIMYDlHyfXJi9mH3jDnbHagiNeADsaCMX/t6lV79PiRN6hhdUuqg3wnq6a8S5dQkzKUSqkpz2uw52XaHgZ7DB/ZszTepBGObApehcVTqw0MT3wsHBl7nuaf17OxKhUy1sdzMiCvZEDe1miT4xftzcvnBhkkkUrbpckxK5Yrbe/w2Da3nSlIUw19fc4Yrv/d9Ds18MRKTyZldr69u6v7TzPZ2aAuWTYxMaHcBkYyLD72MM07KQ3ARElWqtkKuIHXhVfA2kUKij0DM48v2Ow0QxVBiKleICsfj01hfu7WrVs2835G+4JYwNmLHA8gBd7fUc34k4R6vzqtWo7/qGfFbK5lgMjQ0nXWZ+ccNCGU9vqG8ixem6E4a42c33NhgEIwgf2avN7ynNyZsc7SJAdk/ZGqSpJF/47EjTOjaQ7X16YtlSjbg8/uSr5vZua9Xpf7STz64fEjDdcZ4j17+tzu3r9r01NTOhsnRgfsqwc37fGjv2jw+qu/+43tbqyLZYyHIEbsAGsuXrhgq0tLyidgH62s71rXULeGiGfUFydZK+T3g+N4AAAgAElEQVRytrGzaeWqlJUTSbv94Cs7WN+xw6OMDOj3jzM29W7WzhL4vlRrD5PLlYo5q6tGqq9kNalKa2lptIsXhq21td1qWjtse23DFhZW7ewsYUd4oYkNANuoVT0M8nOeEHGV/CiXp+YjB2UfZgSqYT3StFUtG9QWJIcMgAu5a0UWnifyRSf/D3dvHiN5et73PV1dZ9/3OffZc/dce8xeXotci4RIQw5t0xYihYpA2BJMYA2ETiyHhpQoQug/CNCQrAhCBBNgTAcKVmIkimRILanlXrOzu7MzO3dPH9PT1/R9VdfRXRV8vs/79gyXpGRCQSCygcHMdFdX/X7v7z2e43uIXUjzLNZQFK9n8CPKq3lZn0upiaOmV8gbmTtuZO/+RIBjeIb4tBADOKLdzzJ5z+B9wPlIHg5bvZ76U43ibf52piD+A27GrXqMJHH93EulEjK55h7EKFbRN6EYc2R4RIV4zvK+HTt0vlC/msObZH5RLE32+UKRdUUDzXMoFZWVf4Y6jCVsg5wAUCIAS2oxDQ0u91tTI5lm1kFfV6ft27PHuns7LZlGgrioGEPFd+Sai2U1Z5i7zjx0sBb3tLAE4IfPBlzmsQ17I+oRrprhXjaKDfBASPP8NyXbiTxhBXWTxkY9H+ZmBBnzWW2trYpRKHJxpjP+eTFCXT6T2OXGjRs2OjaqzwSYxXOfeTCr+JoYldhHDUKBBJOqEwrEgMSXAArOaKVW4iwCj/VYx3rWmbSlk2ntuVyTVAs4Z7dconJr02srzDnGhrOT9Qt7fW2dGKJZeYkAHDUJ9/tYW3MGimZukNIMfltRnYTzB9ZOlFxmv9GeEgyvBV4SY8EVXwRaCnKEXBfPQwzNANrltTLQDtLLghSrmeNNLOYOeXKUTRdjIsRWYrMCghX4xOtvPGhXw0CO2Otx3FMEizLn3KvM80zAuT9FjYrD9s///a/bv35hr/U0eTHEiqs2ffOS/eH/9kX73EuT8TwOf/fZP/nsZ+xffvKcDfZ6cdhf/5r9L//qc/Yf3vvAy7/wn63882Z/+Ol/bJ/+5gd+tv3fX7erUx83+8rjduJFs99/5U371IEf9dpHvj/0VUs981uPfOPj9tX3ft0+sv4Ne+HC5+zlH/kW/yX3/Av2zVufseeb/vrrWHr1i9b5iS//9S/8W/4KST/NzIQF4Y0KEFBs0BQc2EhYvEKH6W/3DkCvTpTLalVayATwbJgUi/l5pJBGNBfvRRFIhfKtTSW7MXjkYJFerxoJ0Kt+xKCFjqMaAqAyGxv0QpIbdYsl++LBo+KmgHxRlyEoSm0X1ZGO2vKGCvRsNlXv5nrAJf1YtFtFNycZdJKH00w9RI3UfaHQCk4N41BVoybQUBlH0dJra3RISmtPaCI3rCRIAiGjMcD4FNQ6Bpc1CV2D61wHL4OgGS/aPogfXVdlu+srxLs6w06xZzOOBelonCgWR/AQYRPWwRaKaWpKhGenYCVsoK7b72OoRgUbLWMt3T+XlRETgbcq54XMam9ttYZ6dNwXbeeOHaLuc9hR9AVJy3EFanZpdU0JjsynQzfdzVvR1XQ6njbgbFbvMQ+9GwkcPqtSFc2WIFgBsw4DR/kpWFXzChR1vVDQMoDlIEbHFk+UYHApuiH0Q4IMday92SWeoZowzmDxAyqg3r1KIIkIguSH0mVIOTjSniQdhKTGJiAcCVhIxPgeTaQo2UDAyCcIHagDjQAdpFJSwQGJNwiOTDJhWxR1SYarjg7GrHp4ZMxK1Rorlrcsma0TogJUB5/Lgc0fJVdhfsd/R4NWHYA5inAVrXUKiKBrQLPxOwRzBLx8xUZDS1uTirgwIWB3qJEQGgw+d9CZZF4HZkkoHsVD1YvFTuUkcJyfwzeExAvtfDdAVSNFh7XrdPNMhZTD3Ct4gPAeLnfk4y4j0Bo3aEQfmiQifqaaDwH9oOJ+slbFgvn5RQWToAkJQCk4uTyGfy7jw7gQyEsrd/vLkXXR/J3g2+XivAAlOYHAvhFTJOwRKswHamyUGODzXJoLiSFvEPMchEKnSFQgGKxoj2VchKijABLGXJ4tJCHSq3XqN0ERwaOQsZiwBh8RkkIZDcJ8kLxJk/YpAmUKP1EOjL2CMVJwKLPDgpBwNHZ8H4r6zwntX5Llyzq6iH2RdcY4s5YlOReaMmqOhCaomzsitZCysgJB9rGkkOitzUjjEIBypjjzJZ2jELHmwZx8RLzRTdBHs9zHlYRswwYGjti98XuaU9wLybM3U1yOyBlj4czYgjHSoD0uCQKLfTuNgZ4HwtwbY6pgX14umHu6tjnoMJeLcBaN5qSKza7PzvnG/Z44edKapKdasByU6OVFe+edS9JRhj1GYxd5pWw9+1St3R4aUuNBhbJsvZqWKshWNy2Zzdk8iTJGxUIWV6TLzJ5IgY9EYzUPSgyUeSEwbTAm3FQRkOcPOoo9ZH5pxXbv7legu7i0YJUtkrCkVcqgk7tkQqjiJiaPxaLt3LNHUm4UGFZWV2zi/pQK8Ugk0djHtwCz6aamFhWS0DmGPUkzkgSHwi9rS1rj8s0JVGv0xUMTR8UTzjJJgUFVzzqVvaFR78XvU0TkWSwtLagwiSE6zdOd/Tu0DxDQs7dKP7eCFEBByTuFFgqRzl6qcSkmzhA8OyR15r4hFOfRc/8Hn/iEPKRAOvMaxnr03j370z/7up0/N6hm8cjImD355JM2NjqmmOrpp5+xoaEhm56esr/z/HN259YdSWP9neeelQ4zY4AUxfvXrtrg6dOSoUDzGNSr9rGKKcZBauiVV17V+tm9e6d997uvWXdXq5on77z9rlgNFENf+d6rdujQQevsbFdj4dix42JBwBQ4NXhKc/Lq1esCDjCe12/csuPHj2jvHRsbt3Pnzojuj8nw44/RZBnR88Xw++7dIckpSJ84FBHYF9k7kdvau3efS4WtrocmVVnzQsV41nRADosZl3D9aS9QYp7uLFDmOM1RadCzLqtVGVySNOPB5EbTXjCISGbMsDl7xNBUwdERthRqSO4oXdPEQcZDZ0vwM4OJw/MtFPPW2tJo/9U/+Pu2vLJqf/Z//7nkI6qVhEwh2WcptHEWcpazP4JOFXOjvOlylEtIL4QknfhA8ZADECgWMAYUd5Ss69qCVGhIgGPDQAy9YPTLWRH9LrzA7ey6GJPxee4NFBo8oXEfDSNVpA3NcX7H5XP8/HFpz+iBEVkajhyNnkkk1M669MJgjCdjjKkmIfsbzDQ1SHxeMBelFw1jNJh30qxW7BgQ7hGNTlzLmLgnlTeM/fmklHuAmuVz2bNZ8zx7zjNiLZqwAiMJPOONAfZ39KiJr7LppLxa2Cc4S2vTGVvLF8QWIr5m/4Mdg/67N05qJANCg01x/8aGABCYyXKmAMzC18KbNS5NyP4h4AnxBRKW6ZxNTFIs9AIDZx2AgOPHj6vBSoGIA4R4lPuShGIVk9KCzOqXVlwPnGbwwQP7bQXvo1zKnnnqvK2vzVt1s2yXL71ru3bvtd5du+32rSE1KYipQeViwgvKnc/lzF/L5621vV2MNeYOe8C3vvVtO3furI3fG7PZuSU7f/aECrl4EHl8V7Wmhjrp1r/2xlu2H2345ha7dOltFfxSiZQ1N9ZZW3Oj7ezrt3cuXrRnL5yV9NPQyKgVNqs2Pj1nyWyjFbcoqgHQAjQFI9MZ6sD+Y8NJyNlQ7JHPS5CpVVFLEm9IwyB92ClfBvcE87UQ87SBIwOKM/CKYV47WMlzKeIYzk+epYNRYLug5Q1oTNQZPTsa8ZIvramx1RXY+W4UH8E8kZXvTcIgTRIk1mA11VQr1k8jefcOu3H1fZ1VSHK1dnTYemHTWtrbta/OPJiz/fv2qLjF+qJQTpOP+SwJ5pqE8mn2s6G7I5KmApDh6ydphw8ftIWFRbHa1NAkZhJbFiaBM1Qp4vb39drQ7SHFRpxVeAtRZh66O6R7pLGHPw+o5SjxK2Y10rMUPoMR7sCRI8HsG2nEqvtndbbb8MiotwXDeHhM7r5eysly6MkXNI7IW0YAGI1rxUnyrnH1AEequzSRZHaJl8LzfShD5IU70Nj8ggMavc5A7si9l2DAE/urPoB2P1rzRYEXcjBmtor21NNP2PzsvFDi3A8eHOwpF998UzEcbCUYmGfPnZXxOHPhyMFd9tjgEbv01huWSCXtZ372Bc2VxZlpGaLjUVIuFoQ4H7s7LF+ArWLZhkYnrKO/03bv2Wc1NGUfzGkNr6yvWKa50VaLRTt28rQ9mJi19Y2SbRS2rCaVtbWNkgzY4bVThGSPyq8tWrq2as2NOfkVbpY2rK25WbFNT98OW8uX7O7IuG1xbpVdgoezWPlBaLpRJCambmhoUh1meRk1C8/xlPtu4km2ISAfz45YG+ABTX0aq1GmmDw8yoaSPzijwX14yHmJu/ErA8XPODkP3plv8qWocxYquS8FddY9ezhzg5ytt7fP9uzdK2AP8RCxbASBcTZIKUBnmYMmBUoIxWA+z1kXUSK3rOY1i5l6BfOa/IZ8hPiX96HQjr8X0sOAETraOqS0gC/WRn5V3njsJ37Wet0hekuynbGrYUYuiVXmYzptq+vuKaYGC8AFmCPKgwCiAYqkyQcAIDLCHQSrBq2Xl77vC39AV/EIhSz5dvr+5L5W7oHA+2pMRAs0e+HDH1JOg4yegDliDbjEFL8L4IMx59koV5TsFMAjGAveEGEu8JyJ0ziLx8bGQp5XJ+8zqTqQvy8uCiTKnGL82EfUUAh3oiYjzPtwPrF/sZ5jnUryv6G2JtC0dKFC8xG2BWz65dVtCUqNLfKfiYTACbB7iDMBRPCeAH5oGAFgi2BcgTmILQMjlPyAnFl1syCNqxjSPGdV80mSdK6Awdi6JLvHIgKGBFYIoBsGLNb3vNniNVJqbXEgJH0V/E8cDOky694g8VqCyz35xOX3o0SX19lcxpsmDtfi9Tzi6JIUHX46GhV7f8G++cefseeb5+3yX3zV/vevjdiSmbUcfN5++ZNP2WDbqr38279iL/xubFZcsM//yb+xFx9rtNGLL9t/+uqrdmPZbM/gz9o//YcXbCAzaS/921+zf/QfH2lu0Kj45B6zhUv22Z/7NftCUEX4/qX3/Y2KwRf+nh15tEFw5B/aF391j9383X9nv3vjkd9cGbX/9M1bD7/x4h/Y6r88YdnkvP35ix+1j3/l+z9F//svvmez5z92wno8LvCvF/6ZfeljZi/9i9+zlx75dmHqqr306gcbOj/ks/+Wf+tgS6sKhEoegqEeiFuSPiULGCOCPJqd1eFCEATyh0RcyNBkUugJp3C65h1foFgo6In1UFMjAyC62wTnHEBshnTlY3PAkRGOoid5/WFfjmLxRRsNfGKXVgY5FARFp0+qxuwF5nhYxs3fUbQcmNrYQ+GSA8TZBHRuKY4UlUz7Bp7UwcOX/46fg9Dn2CCioZMMC9W8CXrDFOwC3U7IL8zmAtKfgg8oLsylMeHkUKGZwYbIHwo7GwEVFMcTiS0aQjwb9Ge9w+5FRKHPgylx9O+IXhaRqskmSJJFwUWbZ9FluuJ9xeJ1/DsiAvi5514B3RdQ1jIBEs0v3HO5ZJlaCiyblknWWntbq7r0UH+fevppFWYuvvUuoaS6720dnUKQgFIkEY+bN+MobUMCPlC6FIy6XLZExQ+Mq0WHBtUHK2VduvskORSmae5wUNPAYhzXV9AMXpemN0FJ9BRwupzL1/DMI1rLddxd2oeEVIWRwMhhLKSzuBV0UCkQoo8aGgBeeHHarSPeHS3k0lre/CGYQkuZIFTzVxqYrhXJa8XqkQGtN8Z4RCRZyURVOpOpmqql5XvhzBz0wFPZnC2v5216dsFqkmkmk4qKJEH84XUk6KxL6UmHeU+BmsBNPhSVqi3OL4RD0pt9jCXzn4IESC6eNfNLuvspcd4VjBHQM64UCqTbnsluB8ksZ6H5RadMO2OjvkFjxnUQVPB8hu4M6T1cQzqiY11yw5sKSX0W+4wCZQVpXqCNDTo9K30OATGNijUF5ZJJCwVkNR8CWkuJjRpvyMY5MoVgm/tjzep+066lzr8J5qV3GRplTp93KQD2Mi4cxJAkLgjyMEMkea7xhoESBxX4a1QwZQ/g8/iK9E8hi5SAuWY7eyhzXIGfAvOAuKWYtE0T9aKvmkpibaVUeIjG6E6Vd2YJc4qCCHtupOB2dXdta2uzFhln0OW+v7ksAkUX9rfIEiFw1NiGRgamYd7EcbSrpLOClBXjoyZMYLfwfZnAFf0zWDNobGvrJ5hOgmwpSm6wWKJg5p4YrH08HuoacjIGjrWP2DBgblIYc3P0qn34wx+yv3j5O4FdAjoYphzyM14g8WajJzXy3UilrT5X7whA1id62hVH7VJY5W+apr63ck9epOK5gIokcCfgbqz3Z8a6JfmXCbdkJjKWX1uVSbMby9NQoIkN9jER9o2y1SRT1rtjh7351iVra+/UXi15BxX2aAqVrbmtxbZYW0mXlGAPnH8wbz3dvcGMlgId0gwYpwMg8PxnbWXNdu3eJemgmzduqhBLcgUTgH2TsT06cEh+BNNT0yxER1XLVyQr8+vmrk4hz5bXVuzdy+/Z0sKyzTxY1L7PeB46fNi6e7pVnIFdRKEPRgwFKs4VDMtlKg+dG+k00PKhBMR65HXSwZfZqTfI4/mAR8UkUlHreUk30AyfnpyUbMP09KTQ0BTd2U8nJiZFjeecJTEEAbZv/z4VrluamgJwwKWfaMSAtEWOLhwS2p+QTTp9+owkmNh3hD5saZFMDQh85g2IMmQKzp49Z2Nj98SweOLxxyXfhSzm0888pUbO0vy8PfvM03b16hXtoxcuPCEPin0HD4p1yR5Mos8FoL0sT5SaqmKxCCTgMzkfkEd4842LYo/AGqCZcXjgkLW1YUr5nu3dt1fzfGR4WL4crGMQ5G3t7ZqvvCcNOMaJa0QyjaRz9sGcGg9cB/MbGQ+SOeadEGyw82A01HmTkzOC70laTUhuTFWzaoLF4nimvl5ocxpG8ujZcCQ1xQoVsbYbIK5xzjpFhm11bUPyFxRfcvVhX0UmiGYJTXsSvFLJPvXLv2Rf+9qfBoYnMY0XsWnaIoXFZ7nRqsdMSLvRiOvp7pDJ7/PPPWstbW126/2b9sd/8udCw6+srAvRDHqQQgHXDOOLGJj7Iw5TgTAwDrxY70AHFaKzyOfkNf+Jeb3Q4PErSSWxiyT4SDplCB5YmYqzKNxTIClvI0X5/Yh81vuoyeqIaBktik2SUjNE+z9FwAA2Yf+PSXocc/ejcrkovuK5wb2x9xEXxXNEBVuK6vL78Sa4GvcUr1V48AYRaHGkd4hx+L8YLkgslGGx+TW4RxNyn+53lFZTvaqGHI1Mmh3yIQMpGNi6vH+UxuHMJHzZKBQVGyLvwl6OrB+nk1hXDfUyhsbsnucEcINGhRDc4Rzl+mlYguxmv2ddyFdIMbwX2CUvggdKOu0s3gSIT2Q7OKMFibIkknQqkKTt/sSkCjvss8hQ0WBhLNjfKfYxr1kjXDeoYuYlHlmLS/PaU/bu2af53NfTazmBJlatr7vdrJJX7HHlrXds794Dip2HRu7Z5NQDGxmbtKNHj1ljU4vMkpFcam9rtpmZWbvw1AW7duOG1ubBQwft5e+8YufOnbYH09OSPj1+7Iikuq6+d9nlqxjHhpztP3DYbg3dlecEcoKvvXFRBdmUCm8l62prleTXg8lJe/zsgPKpBwsLlq5vtveu37HVwqZVEznLZBusKpQqaw+2NwCkrIPUQkwQ56MQ/SHxkz48aOFMxtpam6yvp9MuX37PY6zwxTqmSE+BmOfGfia/t5RLsopxrjwC+dJ6zV1ibthwNOd5zuiTM885jziPmZ/sbdtG2iG2c4k1l+7ki2xZ60nFPxoVW9bf3W67+/ts6NYNFUUxUcZE+9bdMUkPEhrhUYEnCHs/OTSmzTDLaKbCWgAAiBQmzIvJBw+C1Ifna8QtsORg642OjmndikWpWNbPXRmzt7QIMEDDnOvgFjjvidfYk9mBGFe8k/AG8Bvyhp/08GUyDCAiYbt27RKoUMAMpH0T5Bv4agG0yYUi9cZ2bIpfB58DK1YMd/lLuckyBWgQ7B3tHcpJ2Ef4GbENcRJFcuJHxxP7lzMqHsqsBgTiNvLe5wOa7g4Yk5eIYnFALGSaNZIHbMF/y8p2+vRJNS/x2CDHPHnyhMb2vcvvKW6HVYVx/LGjx+wWTJeVVTt5fL89PnjYXnv1FYHCzl14QiAxzuAiwKG5Obt/b8wODQzY7WvXrRPZnHxBMk6N7a3Wje8ChsD5DeMqJ6YnLNvcaFvJpA0MHLPp+zO2vlG2jVLVltY2bHF53SoUxzerqjvk8/jxrFtjXcp6OlqtpalOviip2hqxIXL1zbawuGrDo5NiLsJQJZ4ipiNmk29BbY3l6tO2sLRoDXUN1t7eoWeRTKSsq9vjtIjixwh6cZlnXtD3kO+mQS9DehhO2ew2WIDnJilENStWvYnEWQDDvw6p1pLOcS+CO+Oe3AxPsaaWBrFEqbPwJUAYz79S0Zro6e2RZCpMF+IM4mruhRhb55HYhy7XozmC1CE5t0B95jEwxeQQ+G4DCEKjntwBNi7FdxjkzMn74+M2+2DeOru7rH/HDlteXbNLb79r63nOenJqcmf3teO8l+cIbxQAeaUgx7bxiNE3F8o1SF4pyC5TafKswxn3vn69lhN9GrxJKkiaAyW0HrxRypxnC42+kg4CcD8D8iQVxmvMnnn6aQFHqRU4i74q2bwoxe7KG95A5jMEbN1y8C8NXp4FYBnGRjU221JdhrW9MLsgPztymmMnTuiMAYR08xayWoBMqzY7vyAwEWuLa6LZwfnPvblvaUJSndQQeUySoo5NJ5QUaNAob3bwKGw3zlma/irWK57IKlYiBypvmc5zzcOgUsDnh/6HAC7ukeFsLcA1eQCPQWEigi1V8wqFL9VKAmhKNYvgT8u1x/2Ja2L/pbEWc+5YM1IdTawIj7OoKzwqF8X8Vfyl8wQgjktJRxBwnOsCcodaHPvq7p27NAZ4CMWmuwCzyZ7HfpgizfbB+bf/Hxfs91/5X+1TbVfsc//01+y3P8iEsD578Y/+wP519uv2sZ/7or1hZi9+5Vv2+SdK9uef/xX7+HbzIt7pBfvit37T/vmBSfvC879on40NCRoVH2u3pWSjZd//Qzvxc79noz8wON/fqPiBH3/6d2z2Nw7bu//2Q/bC7/+oke2zL37rJfvU+pftpc5fsOdHfst2/sJXP/DiH/+ev+8N1HQx+8Pef2yf/tv/gH/sKzzU3GpzFCcj68DQ/+vUomFTEBU8TVCTF42ZTYtAXIyIUJyFgSF6UjolaR02Dzq2Mr3R+9YocedAExtCqCSCExBwmN84vdN1dR2Z9vDLt/PtjSNo6UUTbCFVsSuAIh8CLi8wOqJMqOwgcSPEf7hPUQzF3vBGhApXCWhUXtR1zwyC3WCSDUJeiDYPmjDH0gEYGjNsMFRa6NAKEU9xj+JHsaCAXvT9YFxYLHiiQ4GZ4j3NINAtLn/gesB8fg5EfECqcJ+iYQYDYg5JycaEBF8SLaF4ysZKMs17KdgPRkGiWZecFhqZCtLhCyhuIVNAJAQNYh2RwUw4NjTic3FUgVPhvDnkyQic5872lmDetWR79+yyB9Mz8oc4OThod0fGbGllVbJPWeiBUPk2PSGJRUwS2tgsEVIuoAFBPYDmAYGmJB7D30RyW7oDBA2JR0QMCqEnY25PxhlLkgHGSSZayD+tr7ssQ5h/KjzqXKKYDXvEiyHS0A2HhA6ZUPDgQFGRIaDshRwJbAKQBWLXBN8LFd8olKajSbPPEZDPKoRTdFezzSnNBEHyLVACgR53TkaO9SQXm5vW192lIh1BQW//DtsolW29WLKJqWmZaRGsE0jyvpK/wT+hzuUaouQVY5RN57RWN5BJSCZd25HOflg/BDNCqYexhR7NAU/iBCJVKEw1A9xYS40NIbbyeg8+kwIgY0pxgXGgAABSmaQdORSuk8/RPpFzaaSIqhOSMuWBBUECBQbdQzCwig1HIViCpwrjp6KNkpaHEmnx58xxR4/AACA42nIpiU0CMQzbVrcR/yV8ATJJN7vPb5iC0Fo3WIzBjJJsGWaT6FOI8yaUGixCvuI3QmEmSBcEbXACQIIzR+s4Kyx6Zojay16apemT0N4SUaoKLitVl1MKutw+702JdgzcI1UVvVGhBs1sR3+/5iha+pJlqpob846O6DpBtTorxdEdcQ+IciHeAHO6KeslFui2PTDSSWttaRbyj8/lM2lSq/kXTMXZ4kFm5vNFK6E1yl5cdXM9mpBCYRsyhG1aHzQAmWcguPlz4MBeJZqX374s3VuXoXEzVBJ1fsYc4Y/mXyqp5J2/mceOiPamk6j6GwV5LUm+rOrrjzkN2p/KH3ONBJfmK/ORYhJzkcIL+wpeBOxhLnmDX4qfJzzDXK5e6xRUJ+MOMn1lZUk/X15GwgoJxYolxNZAfogmeZ01tbTZraEhSXrk6up9nw0yYjTSYEsgGcjaorCBFu398ftqktCIwniQL9g1xMjsX+z3+bU1sRyYz7du37b5JZfgASnHq5DA2L93l84XGqqS7kkjqUYzvKxiNp4FzEcMqiemONvr9HOkIthbaXAMDQ8rIaJYzPnnxprsb1DBkTPwRr9o1mIiBiNbKPs06lIwyVIq5MuMu+Tm0ySvFGHwkDhy5Ki01jFuPnRov2SWeOYUfmSSW63Yg5lZLzxJztCbSpynNCZZo/zN3KJgKpk5ZPs2S9ba3KL76du1SwUfvDBAiqkoXNmy/p07tIZgs3HOYMJ56OBhFUNn5+fs7OBpyWvNzc/a008/bbdv35Y81YXHH7OLF9/UOnziicf1XhRBI0of/d+t4MUgX6SES5yALORsfOP113WmM18ZZ/xGmPecbTRx8TAB2c3P1fjYyGseRu7P2SoAACAASURBVJ8iYjKZJZe8WUnchp8ETB72btC93V09kmbhPXfv2qnxoVmBufj4+LiSR94f8Mr169elE4+8GNrJyDmw/7kBc0WFXnSw746MqLhFw4j5zPOgQEIjAHYh5wlVAO6hualBLFXOc0wba5MZIbGdDu9NJZmebyFxaPbLn/pv7C9fec3u3x93nd4EchCO1ARQwnN1mYpGW15d1VhXyxtiUyzMz9qTTz4mFDtn5re++Rf21ttXNV+JKll/zEUBPUrO9iP5dSbegq6XJgZFjOiDwXlGwR1QD2NM04CNgb3cfXMCa7ZY1O8L/BC8KYhH2Fdc0oQmHTIRziTcPr8UY4QmKzGEpOloYHu8wtnHM8Bvg/eT5Nvmpu6JmFTzX3sgyG6fD2LRBZNvb4DTgCjrPbQGaTqH2FDxuExrY+MdnXFnCtAoQ3rHEYiOumZ8KI7hcdPR1aU8QWeNgCI8c5hci0L3sndLwx5D1DB/ufeBw4cl/ckUYI1EGQ4YNZrHSYpgSckxwT6lYcEezr6dq2u0+YVFxRVqQOjcdekwGmOLi8u6BhrmXiz15jnPnL2VcwIGtApAnLEbbuDa1dmmc4oCDM+K4h/PUrrYQQ5VWQJjsL6uHAC0e09Pr3Ik6bwvLwk174WJpMAivGd7S7M11MMuApGbt7pMWufduceesHR9o71/5ZotLa/Ze+8N2bHjh6y5td3u35+0mdlZq29olpzUuXPn7MZ1zK0TdvTYUXv99dclA4Tc7/SDeTt1/JD19XTb/CwxepPOCOZKIwzCSlWMZ5hMI6Njksxpg0VXKNqFx8/Y3ds3bX56Xo2K/p2d9rVvvG7dOzptbHreajONNj27YvVNLVYM85IYC/lF8gziPzZacj3OIYBXdIEkrRhyQvJDYqO2tmbbv3e3vfbqaypaUthkrrNHs664HwrKrL0Y5yo2Cblf1DinAcBcZy9jjvG8MCuWbyHNKPIMvNeCCbw327yhEr1gNO8DK0xMJ4EdaEBWbGdPh+3Z0W9X371qddlagQ36d++1d6/etG5kWzfLOu8BqOzYsUN7K03/4eG72tfxRSAOIbZmj5pfWnIfhs1NN51Op+zAgQNaG3fvjngsH5p9jBnvD7AKuT9ijfGxcYHZ2NOQzSWOw4tA/kBBAq4ibrvrncexp2DJuiM23Ld333ac7QzIWp3/xKHkkzB4iHdB3kcvDYrDnNcUImtB0APcCecB+xeIYJkuF92TShKnKAjAcgdpHsE/gTUm5muQHfaY2tmRPBfFt672IgCB2C3sgZuObFZ5eKusWLMum5RHBQy4qYkprX9MxzlXkVPEiBZGIqyTQ4cO2y1Yj8urdubUgD1+9qh95y++bV3dHbZn3x5bmJ3Wa2FYpBvqrbCwqHN8+M4dZ0wVSjY5NWM9/f3ylZodn7TS6ppM1xdXl6ypo82qyaQdOHzEJu9P2/Jy3mrTdTYx9cBuDY3ZxiasCJOEL+wIFEh7upolpwQzpDGXU/4HCxlG7d3R+3ZneNwaW9tsk/gVbyPzmJnznT81iYpyZ2JMgGLMI/fWSanmA9DCZca8PE7+681xz03EZgisO/8/Z5hL9XAW8XNiS9Z2qtbE5GVONsCcyaNM4c9W8q+AbaRoURHgo7u3R+9NXM3f3V3dAlgwOYnlkN2sb2zU+iD3cJCVM1+JkSIIza+ZPNvjNECT8lsUex9fzLL2dd4DUBL7LWxmziNiJArmvOa7r3xP5wU+XzSvxu6Nax9dW6Mxjmx3TmxjyWOLtcLYli3BGJAfqgnnaHnVTgLTI01RWgd38IVRQ5WYJvhhScnBK14ChkoCG0U0CuTcV5C0FGAseD0FIKByZClJoE7i70EjrlSE4VLn0u2ZtECHxLPEFKxDAeRIPgTW8ufDs2Wsxa5ij8lmtM5pmvGc2cfrM+ThZbtz57YYSr39fbZ79x55jNAcJ85jLeJ/xzxkz+G6OEfZRMVSwI+TphbgQ8zeA6iQ2If5kcm6tJ1yruKm/JaQp2IvYu0Tp5DX8m+8c/BsoRFNjRKmCHsQuYsDPLwZFkHRnLfLqysuBRyUXnyue0PIz2Nvhruvl68FYif2/QgclIx6OOM5lzj7VTvEI1cgFgcWOkg1+IgFKUL3NgPsGgCG+PhKzYFYzMEfOoNCThlrq+y9xJKAzTivJycntyWhf+IbFXt+40t29dMd9vKPYh58sMz93G/ana/8PbM/etEO/ovXfngRHLbC1z9jT978PWv8+3/or6G4/9E5++xXGu03P73XRr/yr+zEix/8/f8PGhW6vnN248WP2meOf8nufLJknzvwK/bbj1zpj33PH7zLn/JGxUBLm5DSocavxQTigcAFlAqbt5oQKh67FAGoQg53IUkTtUq4o0lrpIgLVQYNtdkNnheXlra9EzjInObuByIFWf+XB4EeGHqRj2BZBbbAh4soL9dbp4Ds5nYUDr2x4B4XfMVOaDSC9kfrkiNe5IzdeG+mUOhi45DeXwje2DSiwXMsbBEkxeI8BTTei69ohMThEhSVFARGfkhMLBlTklUSJBI4FSJrHQFIwCUUbjAQEn0sGCELQR719eXp4YdaHC/9fvg0dXiDcZAMgYMpm+szaXT0TGma8Pvq9srA2FHPakAErwB/Lg97tBHZGa8n3iBoG7mWVEA9t1t+bVnvCZV8fm7R9h88JA3SPA0qaMoUW1VMQJbAC+oETlGqJiIWhfTAuFaocmi+LtuiYiLzUpu5y2AJVRT09SkoQJvlwCIhZI6ShIDs4RCQQVZoPG2PYSicRUpebHqokBAZJWqoBcmsoPEqCZqgmRojDZmGBYQ7SYA3OAL7PZg0w2hgnfhh5IU0NUuCzFb0DMAWgyQEQzAqJ0hjEChQSKSoDiNDBXfWTY1Jtx7ZDOaXfBiQkBIlnuaOz1c1IxLeQGBSKKgLpsiu44+ET42CHArqHMCgWnb09esQzlAogt0h6YBF62jvlJkkBRoaFdwXa5+iEogc//ySglHp/9d6E0Ov2fDEUQEJTZpwffzbkTAwN3yN8EUh2+W5fJ1H6S++r+QxmIG7xBfj6QMfp/HDJkJCBRGn+4PccDZB3Ev4OzZAhCQKclTIHHEPsREYxzMmXk519+YEyVNE0+t+mD8O0FPQw5hwzdFDQoi0IBfG6ym8E+ipgSDNci9GOTrJ/Tz4Q4FoZYWmESwU2B0U/p2Sr2ZlMEtnDy9s5BX0co2SRmhqttnZOUdLhyTeR9qDZcZQiBcYBw0U3pE7ech88/3Om7j8Gz+L/OqakqwQh7t8ScmLFTxLtLhX866PK/QJeyhsECW6zE0vfsVmE3sY/0fndt/+vXbr5m2dXTxTkN6x4BYbexElQ6JP45bxooDP/YtVk8JMrShkfgw6QbwKrZ3JCD3IXTEmrM/l5SVr7+hQYBt9SXhvCqHsK6CG0JZOSeva2Ssk4dyXmnj6f0bFQhljq5iyCczK0pmk6NmYuEpnvbXNGptaZfoIepZ1TTJEEiWzvM1gfC8WHQV2fqdV0iY0Frgv0MpiU6WgIFesIVdvacbVaqy7u8d2IQeRToq2TlEalsLE+H3r6+q2hozL5MDq2Hdgn57TwuysTYxP2K2bt+QZwr4Myh3kG6g85ixNR1gEkp4Sc8tNh9nTuZaI8FOSq+aBAgBHawWzYJrxjLev/SALBnrJYHRkVLDEyBrT8FMnT4hNsbS8aHv37Bbjbnp63s6dO6W1PHF/0ouwoaHOMwcVz7qry/reo2I261qSQlvW1FRvp04eV+Gyqa1NZ1rFUiqmc95LWjDhTCyK52raprNqVPB8AXEsLszb4MlTapxwbefPn7PR4btWKK7bwOEDNjY6qmIliQaFEwpweFZJf9+qkphDogTqfCblZoAuAVmjJg1f7Mcgs4mf+FzmKRIs+LLMqvHQoqQQpgx7F+PAc2btkUzevnPX+vq6tb7Hxids184+yV6B2IWdgw8MDMUTp07atfff156/b/9+u3r1fWusb5JRJUnv3TtD1tPT475my2j97woeZPngKZG0mmrChodHBUqgCYdEgprpm5u6L9fq9bVPkRb5IM4WCsaYBCMXaVVHENPwNKTPaiuK/ZCt/pX/9pdsemLCLl1+31byJWtoatezEdCh1gEpfE4ynbNqbVpNvHQF35Oc0KpbW0V7/vlnZf4KEv3L/8cfiSWTyTVaIpmVTnUmzX6BDJGzRoj7SJpp2MUYkCZxRIi71JTHLjHmjFrHis2CJJOKQSrcuPwpe05zc4sKmkNDd9wzKzQTKO5FzyNJQYWieASlPCqZIn3s9XXJ+kU2xbbhJ4kwSP8Ql3j44RKVxKawPWiCyocirJcQPgczdC/YU2yXPNi+vYo1QInTzC0WQaq7HJPLdcDSgI3hjXHOMYqvFIxz+D+lkTak+UuBMWMrSwAhaNCz/ktiaSCzpLFOJpSDuEym0Dk6ByXdmKoVoIqCDHO+VKABhjxVjfwcaDrUop0SznXkPoSS3dwS8nl2YU77OMjjppYmW5ibl54/khMgiymAOKAI2a+0dXS06nwXWEq+ZGVLCbDhPnCxOax9P1unecK6VcGDZrfDczWWxKO6X2SBtspWzK/ZoYE9tm9Pry3NT1pdJmuXL75rJ04OWkNbu73//jXodLaRJ86ikYK5bsLKMpTGH8LlRiZgn+U3VAh/9dXX7MD+fWJQLS2t2tGBfYoXYDByLhNLsmfDQLvy/nU1tGFDvXnxbRW8QUfD6D138piV8is2OjRszz93VGP85sUralCMTMxZpqnN1koV26pJqhmg/R1GXirtYASrSDdfMZdkxkBysb7dLw9BFZf1cO+p/r5+ScyhUR91uXkfCm27d+/WebO0sOjPlTOjWFTsgdwNc5ozkmIY108RmdhcUh1CxXLOO1COOMcN3/0rMo89zXoY70jfH8AXGuoB9XtwV691d7TZzfeva11gLH58cNBeefU1a25vk1QHEls0hOSNkHRzedh9sK6IrbgXADs0KiqsX4qyJfepoIjKeuEaaUg1NNBIdSYuGTSFYfYfGA/EdMTqmmuKddLaC+7fvx9Q3J4nkNNwBsbY1sFA3rAkJjp08JCumbOF8575zjqbmprR+BC30wjlGuW7lUiIwcYeSROa+Qj7QrFOKKBullzKjjxESgYBOU6xmMKm/BWiQW0AL3r87zWBmHdGJpgX/5xRwfken9kmXkPsC4xNFpDHpp2HTTQ7bzeu3RQTEWkr5g6eUcTAyBQj+XT69KBdu3ZdksH4o/R1d9hfvvyXNnjmgO3a2WPzMxPyYAR8B6ySmI7GQH59RecnDY652QXr6eywfbt22/LsvJXWN1TLGB0bt5bOdjUqBk6cEIusWKjIqBtfkqHRcUuk62xlfd0KZZfmw2Ogt6fders6LM18g/3JekxlrK2r2+7eu2/jkzO2xdgZjNtQCIcBJrabNySYP8TQAu7hZSAZtSANG4yLXeff2fwUqQXiDB5tUbVBhdTgK+osCI/9kRhdX9uwXDbpnnBV87+Vo3leG+NeGB/VCiA/b4DXNTRbR7tLt1ZBMonBmxE4gLna0d1p+/cf1P7AnGfusSYjWzDmH5w9XBNNNeYkRvcAGjmfBHLDOKfqnlDaa4KJONdFzWGjCJPPpXbvjU8ovkOGECbK7Py8GKfku5IMFMLePUAB7ZSos1C3AuCg+nLYMzj0AkhLzccgK+31nNj8JA71gngECXB/7jdCjcBrMu6hSXPI5ZBiUisGewCrUS9gHI4cO+ZqAwHgx3qDbQjoRwV1NaYZF+p7W6Ep4TLOkn3c3veqOp8AJXudRZujrokYkGcxNz+n/J/xwJ/KDc2L2geojbk/Sl7nq7MpAZ84M833B2foRwBTBeUM7d8uL0zDgmtlnySe4Dqcze8ND81lySFHmWjAvfgcej7x6P7N58k8XE0vr3vEGqPWW8iVI+CR2IzXkRMAroh1BhrpjD97WQR9cP7zjJWHsk5gIqkBD6jGwdNeP6TB5g1iV2rwnJ770PwP5w0/J3aVgXjwwnBAiQN8o9rDtozxTzqj4vPfetNezHzVDj7zWz+E4bC9h2z/45/8x6/Zl56a/IHi/wdf+fzvvmTf/NiqfWHnL9pn+WFsVBz+LbM/+pJ9/imzl/+nX3xETooX/c0bFZ/68tfs9w9esRce++/tZfuUvTL0zyz7lZ+38//moSTTj3vPPzAKP+WNiqNtnY5CC3q3LIDYqJB2G+auJLhCodVZW0ebCjYEVnyxiDo62oWyYGNiI2Qzigs96r+CLGRRg8Aj6OHAI8hk02U9SstYFPZQBN5Wq3PT2siSUGE0mPHpYGJjp3NZAbnuyFdP+kh8qYt7qyAW8KPuG2wIXusbsmv/0agggUYXnu6xuvShrk9xFQQdCRJJBxtHNMXmRUoUQ4Hx4YboCcjDRok3Grg2uvh8+SFb0gHq2qpusMSXy6a4DvyjBVa+5wXT8P6hWxzv0pPm6HfghVZ/n4QzPEjgSl4c5wCPgR2fQUDM9UtqSN3uH24YEsdZfhU0iwJzoCENrXvTWpsbrKE+I5RGX2+XLS2sqkhR19hseSRlglHSFo2e0KjwjjdyN44+9Ot6mBxwzYxfCQmHoHlMWYPENBY5aUgIEdrdo0OKsaYIxFzmOinmE5zE/ysQCE0i7tUlDBgXtKb93mLRORbM9XBCYh9pyhzYKh4LgYmxtI8b/3bJG++ob39JWsf1mAkYhW4M98fBw7pgPvJvFTdqKd9URL8n4KlhbldrFHTQOCCAggmRTLv+d52Qo3n9Pocrmv5u2u2f6cEpgSLPznWNSdacJUChqMF1toOOPMEDCDDQlXv37LEHD2aso6vDGpoapOktI/GqKYgTCiNozDIvaEbIoLaladtLgHsjECSZwmjbaceYa655cSsEry6/5bI8kjqTDFWdErLIvNLzC/OEgi6MDJ67koetSthnHF3rgVf4m2A2GAEKsRWKoryGa/B1S7GfYsDGQ1SEGoDO+HA0UdCRlJlrReagKxTpJbNE8w9tZEdyq88E8s2QfmrVfqI5KAQGZlg+VtqbAtOLYjeSBZFBEhEujuz2OcWa9mAP1I3LO+naZRbvHjPRuIznATKG8aEISFEMOi7MBLwFSOBJfLUGgodD9LPBM0VeGJIQI9D0ZJ69hWax9p0K5p5eJJIMH3MXgzN8TBLIWRTltyAJDeYiAScNSOnHprVGuX5nMrmsCfcOqhcJB/YIPt/HA71lfH6WQmDoBpEU6WEhxTUdpdbYW5HBoUCl9alAkqaS75FCE9G8yWadbaU9ENYeibAXBUhEmK9Cl2GuSiBJEA41nSQjE6RcIsW4BvkwR1Bz7kjuJXhbMH5IH9XV56Q7XGPQ5rdsz6490jxfXl7TnKKZsF5Ydy8WnVU0zQI6Rwli2fbt3Wt37tzxwDycGzzjZAY0eFWyURura1baKEii6OiJ45bIYtqY1nOgQLaytKwguYlkERZEU6Ndu3nN3nrrks3NLVpZSPY66+vutZ7ePjWbl/CeePBAaGnOahKXiADiWjlHKVICOohNFQwHuX765pKUQJouIDEpWNJMYMzkZUDjniKuUM05O3niuI1LUmneTh47IrQm8xm5Hp7Lytqq9ff1Ce25vrruBUDAFpm0GltCws/NW39vr3RtedbsLRaK2W2tjfbscxcMA29+1trRbaVS1daWliVfxb5T31gnFh2rDzQwBcz74xOa26zjpfkF27lrh/SJaVa0trUosSsWYaY2SMoA1CbjRBEUXWgKE+7pU3EmgYqyKWtt7dC+ODIybEcHjtjly1clvwJSk6IHrIIjh4/InBwk+c49O+3ajZsaD6R4bly/Yb19/bZz5w67fPmy0LzEULzm0MEDQlteuXbdzg6eVDGLfQMAABJa3Gtff7+MFFmXoHXvDg+rkQGij/NWzRIQhUHLmD0aCRLGATYF64RmC4UfCihIvMGSKpGwJWodwNJQL4kO6f1XK4YUHU0XzjWYiQuLK5bNAOwoSiKNHlFTA1rV65ZJbdkv/deftM1S0a7fGra/+N5leRIw3ziH63MP2YC1qYxt8PnJtNUlq9bV0WI93e02OnLXHjt/2gaODqio973vvWaX3r5ipXKNFUoVea1QsCfOpGDI3sP9gkTF2DYmkLGQE2O0GAtyXjGXHAVYdVN59LzXvZjI9xmroEUnGS7Oh0tvX5J0DQcHMbfL+3mSLW1iSUlFreoQ+wYvC8adz1X8J5NyZzzQvObc4rNoarJ3CrQCO0wayf5MxIjG9yyZdAR8KNxyniBTxM+iXEiMV11PH08xGsdeCGW/oGHGnu1FDhpIzo7h/3jisJ4o4lGMoMi6MLeo8SJWW1pZ1lhk62gYbQTWz4JLiajB7dI9bhCaUgOgo6ND0kvEGczP2kTW7t+ftuJmWY3ATC6rZvDYyIiac8zzTuTsFhd09sncM5uyudk5a23rkK59H3HW7JzmKoyK9o5W27mjTwWxYrng+UswepdvUpBZJG7iXjgjGC9JClaRpKEBsuy+L5sug4VOPo2FDM+oULTHzh+1J58YtOLGkuKraxcv2579B1UIujt2T2y2uQcr1tfbp0LrynpeDIZKwr3auto7bHJiwjbLW3bsxHGdDxRoafSWSgXr6eq0vt5uefwQU7LPworasXOHJE+QjytXE/b+tZsqKoEITtVU7MShA7YyP2OF9RV7/tnjypmGR6cs29BuN4buW7EmZYWtGkvVNxoxvlhNwZhdbFaMnBMwBWHdA4SQivg261IMTIqYhkxqmzU3NAnpngysSfI0j2dLKvrTIJ+ZmXYATGDe8hzxLRAyFvkpZMIStWp8cI5zLtXAGqp4s9+9R6rOXAsx7I9qVFDodLZDSYVj5s+hPX3W1dpqt6/fVJyM7OKJwdP28it/aU1tLTor2VM5k2UGXDUbwDh7bl4NBNYcxSj2ZyTE5mB/B8Ng2EEH9h9QfKe4iDM/yMaxRpTnBrYBwAt9DxbusgMGyAGmZx6oiE4xkC/k2Fyq2It4itmD7Bz3TZH42JGjdu3Gde1TfG/Xrh0aK/yYtn3jQBzzesAdeDzV12t/AySGzw+NCuWkwUeGeEr5UABx8X9JYuYfxjdRQz4C82I8E/dTsf0FakMCkEau1w/4fC86StVdDFQk1ADLWbVoZ86cEuv02jWa9B0af0BKNCcABO3Y0S8ZqPPnz6s5v7S4KgPu1uZG++53XrPHzu+3vbt7bXlhRutn54H9tjA5rfhp94EDytHI6zCUHrkzLKnegf0H7cHEpIAvxDn37t23HJK6MDhOnrTRu8NmVdQoCja7uGz37k/ZVgJkPntVQLaBGG+qs9amep3xPe1tVlvesrW1PHQ/m5xdsPGpWUvDYsCrcBNPGLN01tl0Kt7KwD5vfb2wa7zAjCea8lWeidQbaNh5kV4ytTJHZr8OJsMBjBeLsJ4rufeCS9+iUpC35sYG389Btmcz2suYL7EgLCAVTQRyE+QLYTuoSY2fCI3JPvl58L6cKTUpahdFyWF29/TJk4s8hMK1gF+R3S3fAE/QBTotFy2b9oaJYvZkiJuJd0ueJ3Hd5N7yEU17QRl5Qc5EGo40xycnpuQdxv/bOzp1frKe8BxjjGgu0ljM46lEo5najcBKLr0mVQXJuwo/5vllOGtZzzQ6HITgBufyNgz1IRmbb1ET8nVKXYuYTfJykrD1WpLXsRxEu2U8t4T8hdj7AHcR81G7ktF3AEfkMhln7G6sKv+PLBrmgK9RB/N63ozsMj5IDrygQc/vS4IpAPOoJ7GPkQ9Q+yEuZD/jWU1MTtndu8POaEeWmXg3vDd7kktUe76q3HrTYxVyM77W1zd0PvD55AWMF/VEnhfnJ3EZ8TnXTHw6MTmhfFEAZJoFUmWgpsN4et7OemDc/HNjfcZlA6PXhI+775PebHPAo2Iw4rHIktDPXZ5TjaRQO4mNCZcrd8ZPGFD3zsCTDSChedOYPSsCt9jnWAMCz4l55r59Md705owzlWIj5CecUeFG0Ufe+Jzt/KVvPCyY/RX/ksF18cuW+tAX/+rXf+ILNv7vT9iNKNO03aj4NfuCBemlriv22Z991K/ib9qo8MZEzzd/zQ7+6iVd34t/9C37fN9rj5hq//j3/AM3+tPeqGjvFOIuIubZnNjUWNSgMykCu/4gmsQ5/eHsBHnD99h8QSFIYocNGDmMghdDVfQW6qTiBf5ggsRrWXQENMhL8T5RMy5uUtEIzWU00CAMndJAP+RgcdRwVYVrDt4o9SKavDwP3HjR1QEffqmAF1DXbryN/nqtd3gTMCsyokaDBGUjS6Xp1rrusHTe1YF1aZzY2Y4aoSqMIZQXkMjf97nIqUivddO72oGCC2oDzTlpnge9QDfw9eCAjdoLto6Cj8EaAVE8QCIiWWmb5KocsRJRJ4w5exwbuifGLmklg6zAROCz2fh0zMuI1xMo///DjnQszPL9iIzRdYhNAdqfwuum7ezrlpwQFMDGhmZRzaGkFnhPAutaGiIUAf1wiqh4f15RBseNbxWgS4+SjdllWfjsMuaDuZySDw4AxoprplhHgkvwyRwA5cqhxnuBkPD56RJMvF5d/FCsVpE8IHhkTulxz/Y4cBA+yjDxH/s1SoJMybMXeYUWDQVF/7k3NIQqY27Sdd/cUlLAtUNfZ/4xlvyuF0/T0uaXRBfXCIoESZCqCRXMp+/es9cmpyYdiUvBqKHRmppaNV7efDKZCqtIwZgH0y7mmc8vtNHXxJKQtAVyFoUNFRhj80Z0SEsoIGA8s3UZae+SbFNMXV1Z1+9R9Oa1LsEDtbRWSYsOdiS7grQZ+qgKrIQyqChwoYHEoa1ghMZhQD5EVA+HsUvQOJpS8hIqxjvDApQzBzvJpjwNCGICi0GNpNBcYMyY7+wj+GqI/aF9y82CQfbyc4pdfPF/0CTQgQnQkIhyKryvUz4/SpRRbCBY5/MksYJOK54ZwRRbRalyWQEjQbBkQBLeHIzoiZLGfgAAIABJREFUIF5DAUWG4ciiUQABESwpohrtw4vzyAZhyOkUUw8k67fRcSTFzEQ0XSmYMpfZ1xzVCwXXDV6RfKF4BIqP4JICE4UaXhOL9wTxkoGKZmHo/0LXZ6yCtBw4IlFnzen8jo2mEF/SnJSKgjJM/5t1u0RTuLnJdu7ZrQCWJhNzBikBEO4kgJI+KRYllQfKm7FEdubtt991fxZ45oGi4oXwimjE7IHu95IW6n9iYsoN36tVFRj5FcaVAqwaVoFFR2DJeXXq1Cnr6Oq0P/6Tl0JAjNwE44hB/brLH0hWxxMh1juSTKWKF52Qe2IeMI+jNEvcm7l/0ccpBOZg1MEMRD4mYZVyyU6eOGnLS2t26dJ70tPONtTLS4LEE8k7jGCj/CJFBO5h185d9t6Vq7azn6JVk5IRrmts4p6lsrVWWzVrzNZZY12D7uf44Enr7u8zBI9rky5/NzszY6NDQ3bpzbfs0OFDtpJft/dvUGCukaHpgb37raWpWVR55ECGx+4J9SrzOQqbwRCeggtLh3XFvEsnSYgSAjyINSNkLWOuLM51vtWTdkNBNRlVxFzR/eNzJNPKcslOD560oTt3bKu8pUIhe/fa2ooXGufmdD5jsIq2+pX3rmo+UVgFJc2aROYMSSrp83IWE4csLKhQTrOksSFn5x8/a0uL89LCrW9oUhGhvb1TTQn2h7X8qjU0ewGZJiJ7HZJP7OUkgxS1hQxUwkOzC8P6RpufnZWUgftDtMhjgnX7sx/5iI2Mjlp7V4diDtdSL9I61n5KTPHWW2/a4YOH1ZwoFfJ24ckn7dJb7whZS7P6xvXr1tPbq0bFq6+/Jp8JxpD75zxhbyABFyhCBVWXbwPF6obxLcEjpSADdRr97B/s8fMLcyoK8Fr21YX5eaGtkT/gWilGEB8Ry/X19drquntWiMFBXCPmGAzDhKVz9ZKnQRaO/YLPfuzcedwu7eKbl6yxPmtogXf39eq5MMEmJ0HwUhjEUBRfJYyTk1bI06As2c//3Ecsm0za5IM5++M/+7YVKrX6HOYASGrQhRPjU0LHM6ZKxCtlq8+mbc/uHZbNsm+U7fT5s5KIW18r2P/10ldtdGzSsrAqUpxJBWuCTba0pEK45JxCkiq5C8mUFTTP2dvYD9SIZhQjUyEYyMosMgRa8hQLTD3FjQBKmO+hCMG5QMzGfKjP+ZnBOSAwDUUReXw4u48//J7Hpd78FtpPMZEDVOSzgGdazhGPrAMBU/CSCPNWgBrYWqm0ZO1iI99RgGUxyyhMgsxnnXNOaQ+toQHP3uMSSvK1QeIom9OaZ+3LNJPYNkgmtLS1WKlcCKbkNdZUTyMIdP+KN83w+shvuOxnYUPxnBq4OoM9cSeel0SMVbS3g+KVgBNsxjJyDA22spq3haUlMSpAZPKFVIli+0JR8iOLK0vW2NwkGSrYNcjWES/Nzy1Is5z4DKhsqQzjac2euvCENLJTmaStbuBp4pKAbS1tWuMU6mCVE5tSTKfx8WAGxlKz9fd02/CdISuUuX6znbt3aG+9cuV9a6DZu1W0x84ds9ODR6xYXLFsKmXvv/WeHRw4Yi1dXUL7Tk/P2ndfuWZPP35KgJwrV6/bIrJa3F9N1Q7u3y+TZs6jXbt325UrV+S5MzU5YRsb63boIPt5k42Pj6mRAOqVRj7xKAVmmHtrhaKNjt5X0ZnYsy5Va2dPHLX7I3esZqtkH/7wWclVXbp0zWpS9Ta/UrANS1qhkpCEDUwJYhnenz2H+QZbZ6Owbpm6nJqWFFwrFfzPcipGEXZvbtIsS1l7a5sKXUgJEkOpsBq8yJjPSLNwHnEeIgOm2LxitpZfF3PDGdgUrUVhVKGPuA/pWQE9iEtVSHepXOZdZEh9kEm+nc99X6OCHnrFBvbvsI7mJjEq0sm05O0Gz5+3r/8/37bGlkarJMg9VnX2ckZwBp05c0bzmIbhzZu3NB+RdwLoMjM3p/jM8wnfvwEJiakQ1hzXKxPk/IYXukpl6+/r0R6G5xtrjXjl3NlzNj0zI0lAxdewlBS3+T1rnYXGJAVQvjif9+zeI0k/XgcLF+kj9hfGCIaNJJYTtZarrw9ZtkO3JP2EnyCF8OAdKUljZD2lWODPpFFymF7MJQ+Wn10AqQiU8YhqQDTBdck3Z14IZU7uThEvAYvAlQ2qFZDosFQpqlYtl05YorppTz55Xr40N28M2Y4dvRpr6hw04js7Oq1/R7+9/94VGzx9WrHD4nLePvz8BWtuqrfvvvw9e+LJAevrbbOVuWk1xnu6u8V8HB4ds/NPPCZppdaeXqupSdrm+oaNDQ8bnlrDN29I9o34D0/G5uZWNeqPnDlrQ9evWyKBB1rFytRaNspmNNRhrQIQW1qyBjyONotBwipt+aVFq92sqGi+XijZvckZm5pbtGWKv5msGnCUXWlgqakQ8kjyOeYRTUzJ0wEAQw40NKKZ7zD5iGvl1xfyFHlzbbmsKuPPOU++Rq3IDdEBvMHCT9rqat4a6tKWrgUQh/QTptg+j12ejEJ7UsCR/Fpe+0oVhS6a2nU5NUNXlvO2o6dD71/aLFqBhkMua41NzWp4AzQhvgFw4zkd7DzOXgcuEa9Qu+LZE3tR/AX0Af2FNeVS4c5idPljPz9pOOMrhXwgOd7U5JTWBY20uly9Xbly1UaGR92wvr9foC6AG/enkTHOqAG1sLxsG4VNMW0AYAGKEAqf8xQvo7DOVJOR2oU3MmCYsPZinQN5cQE+kGOC8RC82niGPAfyB4C6PF9582VzgSFDnUEGHIq35W9mpn1nR/8OySsix8Uex/4gwENNxerqnR0QYwX3PfX6kBQ6Asgq+iIiaS62ZfCPYt1ROwAM2dYGeHlVjdGLF9/S9Z45fUZn1MjwiNYgu9rQ0JD2IckwUowP+beeSc59dNzUGqUF1sJqkH6qtdUA8hADPzbBxGpyyWnyP2JdYk++XFLOAXu8nue9jAx5YDy44onXCrkHJqwacJIhdnCYsyaQi87pe5w/vD85npodIR4kX/Xandc2vJnm/mTxy4HGAFu3lDcCsmQOS0Y7/B5zxFUuAgM9SEWx53MffA41SzE0qC3+5HtUeNG+92uP24kXt8fqr/jHCfvSxT+wj9z7onV+4st/zS/QdHjepn5oowIz68/YWy//gg2Mf9X+0TO/ZX+ud/ubNSr2/M9fsju/ZPYfnv1F+0z0xvjkF2z8C4ft3W1pqx/3nn/Ibf6UNyr21bmUk8sLOcKNTZgNmECDgMrZEUlthtETAYo3XxwsJG0EuEqmwgJlc3G92jYlMaCuCY56unv0PX4f+pz04rQ3OAMgFiq0sCOSmiheCF/MY50K5oFVWt8DEQMCMVLsWfgy0hJSPjQpHioXhaTLZYYi/dEDWTSInTlBEsrGJe8JmbxRiHWNdIJiL+77mKlTngi0u2AmFWWtHm5L3KN3bBljaeYFeRtPKB3Nrt8LiH4FbCFY4zXxXhxh/lAuKzYuvFnhW6EMmcJ0juhsGdmp+OsST0pc0f8LWv/8diymR7ko0A7xS+8cPuNRCq4jxf2Tq5tofyel6V8u5q1XPgrLVpdrsGK5arMYZ6dTto6Jbng0kj4ICHDX7POmDQGNd7u9WaAGicwLg3EUCN0g/USnn0NCLIBAqZPRL2g12CPyWknL1JVEyfWjHSWo8RdS+eG9+jUFwyxpNwbtyPB8/Hl4kixjrPB8YlFcTabwudHYNxYRhMQKHXChWMJ1x8NOGpsxmNcccC1MVx2lWeBMABI/GhUcTtwbLIj5xQWxgnh/9LhJEAlWMQ7lCzNxErWYHAjZKNYHTROQ7z4GFEUoAtMMooCsOaumyua2IbeehcwXm4L5E+gOZ/9w/yQ2zDdHgW1arQzvXPbB0TqV7aYCrAquWciBUFBxhoevMT0bGlah8AHaOLKjxOYIr3Hjc2coIHlBoEZg6v4FIA8czcXe4AWOpAxlYROwxwiRFRqEkU0S1xvJJIFElOxw9JY3HvV+4d74PoGtkDrlslAoakhIJzVKtUWNb5c4ki8BKDyZdIKocZYLLBnGkGsmOVQAl80qeeGLeSyKLkEsTKFQtKbp8tB3ZVPzhf2YRhG/UyrDZllTcsZ4MTYUZShYqVAQmASSDAlm46CdlZhCu6ZApqabN0i8UQSln8YNlHR0X92UUhrQopL758AEAtlI4Ly0uiKkJ0URCr1KOMUYIPAmMCT4JaCm4OkyQN1dXWraSOomsD7ErlOzOi12glgQQdudoHNwcNBef+01SVoQnEdD9shE4TO5ZjHlxPLzBjZBO8Un7XfcA0jqYlGsnshQifJP0cSuhD4uDRAa3+xhgVnD6+Pe7sGr7/dIQsCYStRA2q8q+Dx/5pwVC5v2+ptv63mtFzz4rqlFxqBOGtSwT0gMxJDCb4OksrFR1GrGMjJiaHCUMQTnLEeOJLCoKIofPzOohGJyetpGh0clo7SyuCjkT5G1Vt9gHV1t1tPXq4RrfWVNiF8KbrFpw3rlvoTUDGwTN4xnnTlQwQ2HvQBCAqb1T9GCgqY8n1KKJVinFKtIAt1sfk26tEgpUZCFrbd7505pz7qkF3r462IVsP/xzF26w8+PjXxR85d5T7FTsmWgmIOZHlrNILCl01vdspXFeUkzHR44aO9dfkfSTMiSkHynkhlbUeGnVvrvFFhzjXV25epVjTvjS1Oe50eCO3j6lHTyc7mMTU5OKLkmnmIP52zw9V5rQ0PD9tGPfkRnkxJb+QVUtKcwz2gEzM7NaZ+i+QVzhYQflDpoUNhC7LFrKyuWrcupaITUHu+tBllgJZH8oMmbSTmimEY0c5LnR8G5Sc3tJpuenJKfAGPO7x44dEisW/buzq4u6eGy2yH5yXp969I7th/kdalgU1PTduDgfiWRrHc+g+eKLAnoPvYYDD/vDo/Y3eFRj3cqFRs4dNiOHx2wr/3pVzW+AFwOHTkqjwea12vrG7Ywv6Rn2tHWruIHHsw1VdZiwj707AWrrWwK/T2zuGabiZwlc41qSpCYY2D/nZe/q/2NZrOK5oW8pTEZzaXt2NHDVi4jK5C0C88+K2mIq+/ftK9/41vS+8dLizmaFzPRE2DWNwUbIeRDc0I+ZqHp4OhIL6JF0AJrUsAckKKZjNYqTVXtETq3XQJAMZtQn+zZ+In4fkucqfMoSLM4wtLXWozdtO8ExLFLYDgiLzYfIto0ek4IPbiNIPf33i5GsLaDjxtN+/U1Z5CpiVb1uIJGBY0q5E66uzulK728tCBzbCXx6YwASchn4BdDI4Ezm+uFKdREETcUN9nPiK9Tta5XLiabAgqXneVzYcUVS1sqWMnMOsxzmhYOKMCfbUvrhf2EYlhtIi3NeIAyFHBgVDCZkHai8QVbBfYAHhgUz5H/QH6M62cPIZ6h4RJjvsYm5Ow4Lzds//69ai7VZtM2M/tAeRD3QPzE4EjOIwBhlpdWNKf5fnN9k3wrOHdUMMtkBIZgfeMTtLa8YCdPHrLdOzpsfXXe6tNpu3n1hp08ddqSjU12+Z3LVihs2uTkA+vq7JZU4PDwiG2RG6mgv2U7+3dJIpESyaHDB+z1197U3xPj41bYKNmRgb3ygXIAiO/fMJiECkeKJ1FrLZ1d9trrbzmylcKmmT0+eNSm741a2jbsycePimkydm/GqrV1dv/Bsq1v1thWMq1ia11jo5rK66urrpMOyjWXtcmpCbHfunvw2FEPwWprneWLQTnNxXS6Vnr6aNbfvHVzG1Wqs0eyHyXJJdE4ZX9VXhUK4yoEEXvIbyv46bGJbcEYbrTV1XXFJZwNIK8jsMGBHI/EnSEB2s6zFOcFduUWfkoeyx07tNvaG5rs2pWrYnVk6hrs5OlB+/Z3X7X+nb0ybYXtLWmmbE6NlSNHj0pKb9fOnQIayAto3VmAsCrcs8sBWpwXe3bvVqNieHRkmynPOcHZy/XBROxoa9N5dG/0nuQgWSf79++z8fEJWw7rV4zMwMoQO19IbD+rIxqYtXNg/37PT2TKTJzioB0xINY3NNbuYUaegMysF+3cuJyGO3/72PrZ78Cz7ZxRsbYjyWXYG0ByLmPyUDYnNnUVY4c8LcZoykuVH7GPUVh0kBvndXWzYlkakyL2btlTTz0uH5mbN4esv7fbTg2eElDz7tCQmq8wBodu37bBwdN28+ZN1SiefOJxa6rP2OuvvmHPPTdobe0NtjY/I9mvrt5em5t+oPvce/SIXb/iwJL+nXu0b28CuGqot3s3bgoIxXl+d+iudff0Ks4eGDxttyXhRnPZ5ek2KFbXJC1fQnWiJCAYDditctG6O9tkps2CaVS9pWyr+aItrq7bxMyc7d6/XxJQ+CUgbwiwhxjX9xgHxkm60Ey+VKnalNDtnGE8B8YWNQJiQp4hjVYM1Zlzql0AOgmNLuJoYvgI4BTYT4wK5HaSlkmmVFMR6IuibZDwdt9SABI1ll8tirlGs5AzngYGzC6Q+rAwuF48alraWxTbEHcCnEAe0K+pRs0mgEvE9LByeAP8rjhfOU+FoA/sNiaYvB2C0bq8B+T74GsAhUlnbzsTUYx580aAfCxSacVcIyOjqmGRtyJ7WpOqtaG7o7YQZJjXmMswyQLQrR4pS0A85QgmcK1A5PlUcAaMkHMvvijDBlgngtjYdKkD8H/WWZQOkoJDkBfyBh4FGnxg/Mzk+UTp4jq8SRobNC48j6gY4PKVK8GXIXi5heZlZNMoRwzqAcTQQvWXyzpjiO/cg6JuG0grFoaAhM5UH747LIkzNgzkQwEpUHeUibt879Y9P0VhohawUINNTE8JjMHnejPBZSOd5eNqH2qubm1qj/d6C5/pjFGuS/KLYq44cDTm6DGmgKXhNcjQSOCcCJJXUUZODRrOhFD/ipKZapwKnO3y12puBG+5GKNJwvqR93R2RQC/hvof0sc0qXj7OAZcpxj4qnW5tHME8jJfiIljnEdc4mojrgrxE86o+IR989p/Z0cu/f/NqPBTfs+v/o699T+eM3v1i3b+E1+20b9Ro+Kcfem137Gfn33EF0Of8sHv//j3HGKSh3/9lDcqBlrbZWpLNzPK1dDFZvGykZCQQd2mM0rwA8qIIBbkbSzkEXiJtlrPZlwNSDyXfBCifbMs4yYWNf4Ak1PTweTL6UosUIJ5GXjJzImijWNkY4fS63tuvOmSSK6dzgKmyEXHVUiyLdelk2lm0OJ/WH/+gM+CEAcJIUJiPV6ouI0N6+7pVvCdlkYiSBDfYOJmR7L0sIgeitaxM1D163LjR/9M7506K8LlplzjXuhoIWvp5ju9zyV3HBGi4qzM5Zy+zFdsXvxAEyHO2oCii4Fe7LhLZz5o8bl2vntX+CYbDgnpg3qgrs05mETHt5b/huRdvLDP+Mm0KhQcuJea6qYMtRfnZ4Ug4MCdm12yru4+W1hetRWKzKBpMYkCSR6owQTl3sDxz46SVY6YcAM4oebCc5d+pkzMnR1CoCTAdtDYBH1FM4L75/BnPvM+SJVxD258/tAPJQZibmIUAvco/aTiycPkRV4GwS9EGvs00oI2cSwSUCDnS9JPoXkQn4notUKieIHUpZIomniRNQbqvEYSR6yHBOBnOA3+N2hK7j+a0fEaroVrV7MK9HsmIwYEGsSsJTr3vCfJEEU1l9epuvSUaP95yZBQjCVZEtoz6JRidkfxkP+LphqeHagoL1h7Y1BskkDLV+EdgzPmd9CS5LWac0hciU3jY8T3Qfyy+MXmETqRxoJLCsnHQQbPXrBWMhnWmBdFvcgv8yqeea5Ogfb2VzDTisZZYqgEPUs+n3uNRqeSyAjFzPjMvFDkaFzQRPyfwoIafDSXRM9EcmRLczrOYZ4pCE2o1tITFlPDZe4IRPgs9hMlcQG9QoITESw8G14T9xI1LMWIqNdzFJqWYm+guDrq1VkcfHlginmqm466pqXZwuKc7dq5O4znlozMCfBgOTnizeUEvMHghX9vpqVU7OceuF/RlJUrsgY8KKSITmOUxpKM/WpoFMrBRihkkpiIqj94+LBNzfDZJBXBfC40BL31ijSgG6pxRkHPx8CXoio/jGwTDwDdsJY1xL4TdVUJmO8G00peF4u4Yvwg9UQCEExuVVgPjWCeQV1DvRp83CsIN81DmIIy9Cyr/xyLCfkCRUg3dON54UPE62R6LoM9n5tuPM+cyzqKELoDchhVEPgpmTIvzi/b7NyCAvRkJimEEZrboD9BsjNfhHTytG+bfQQCWEF2aPyBSKZ5QqJSxFS3xLncbPMLC2pIEfSy7hI1mNE7Khk2VlNrq2Xr62169oEtLq9I1q2wvuFykMjGsefR0JL0VEmINQXMNHiD10xkOkoKJaC9XQOb60/qXknQWBvS9U4nRdd2o2UK5SbtW+Yv+8+hA3vlf0KsANsBmTWSbIqGFJx4rhTpaSqSjLLHsUYoaqlZncmoMMx87uzokJwd+yfvkWEfLhZs545u6+vvsTffeN0+9DM/o/dZX6eRyHwq6n4Zp0xdxgqbJVtdW1WRVskbhRHMIgMqdODIYUula1UI8SIaMiicFzCoSnb2icftnYsXFRdhKksBz5ufZRUQGEcS4vn5OSWCyDnxXqBxAX1Q7GJtQK/H5Jo11drRpmIMez8ynqOjI2rQwRwbHh1V0Y89JLIMJT+1uqqCLXObseUZAFThzDx8eMBuwWDZ2rRjx4/bxYtviFq/e/cuJe+rK8vaB9m7SDwp1LAGOLdANcOGaW5pUIGuVK7Yer5oD2bnJFujvaNqanR8/Oc+al//2p/pex1d3WJE6PxIJyWzcE/msEl5kTTX11s6SVEd1kfJzh4/bMW1ZavAukjmLJFttkxjm5W2vFnAPd0bHdPfSFAtLi6IPcN6oNi8e2e/DQwcspGRu3bi5Clra+9Q0+PrX/uGjYyNqyjPXsh+4NKJvv6ifrDO+KAPHX/OaxWzyUyaomt6G72sIgjsBl2bFyKRgmJecU7SIGMOc63xM2MDLjKTOfqIl1WsEOPUTXB1/ockOhpeRw1xPs9j6YfsXO7Bz1v8Qtyvx4uX5uuoXBJ7hrl16e23xSCQzIR84lx+jmfNfEZqDJ+IMghYAAdC5FIUdmlY981xpqjYryBhif+Qp0MvO++/h2QN8yXGBBjGI52DnAWIyYWlVc0F9m0vsFXULJF0IKCN+jo3bXULC+3P8wvLii0oivFhMh4tFNXI2sCnCMY3MTKVZ4GUnD2tgmyQrVHMIamFkhoiU1P3JUu1e+8e20pUlYs4S9URjrAo2Cv5HnuaGC1VfFcWLFObCtIoSFU6o5dCPs1I6k2rSwt24clBO3xwh9lWwUr5dbv+7vt28NBha+3psxs3b9vaGihi9OY5bxn/TltAsi0wRpHRun17SDkcDcQ333hTDZm7d+9aLpOyXTv7xajgeXFOMdeiETxnMmAXS2fs3XevuuRdNmfspGeODdj48C2rT1XsmQvHbWJi0haXNsyS9XZ7ZNJWylUrW8oSoHKJdSieWY0V8xuWrqtz6Y0EXmoFeTmwvoQqlz8HBW3GC0QqHndN1tXZZTdu3tSZI/8uncGeD1G8p0lBHitUdxoJ4ozOJhpOFESJk1lvTXUNOr/Yt1TQk/TkpjU3wpRadO/FUJD9IHjp0UYFMTON+62tkiUTzgg8dfSgdTQ129V33vWYur7RTpw8bt/53pt26NghW1haVkMYYJ+aCqEITOGalIXmCY0BGgt4LUXPEwrcPD/iJvZxENL80RkfGMnEdoF6oYY5zWvOpWSNNzZ578nJKeU8xGWwSVibEYDF9YjpHdjt5KN85sGDB8R0Yl9gL8b/iIIc4DMkGiPyV+8TvAPxqCAuYrwJNGlUxPyd17P+JR0T4nrFHDWAARx4ol5S9KjQ6x42LSLAT9/T62hFu1cbcjehTyWWK+w7xWAwUVM1lq6t2tmzgwJajCBlmE4LwELciyRab0+vtXe02a2bN+3YsePyB2Lsz545rSbH229dthdeOGdNzVnLL8xCRBXbcv7BrJr97T3dNnTnthoUA8cGJenUu6PfGtvbbKtQsPXVNUkFDQ8NS6qN5ilm3nduD5HRyQh4aPiezS4s2Xpx0/KlrSAnh4RSyTrbG6yjtUkSmD0d7daUyynOXFhas7Vi2WYWluzk6TN2e3hUzXhMzImhaN4AlqI9IIYXfm01+IxMqakapYDdG8AUs5IbyT+KGKulRYADvpT/BNN7fk6cItY1De0KjCk3tG9pbhAgRnUMNc3dA0zxhQhPDgorFTCgdo+VVXl4uLeFBMDD7/NMYWU3t7VYS0uT4gWYFfxNjYa9nbwW5ji+WfhlwbD1ON0lbDU3azxnJp6WAojOTz/LkfmMe76ObMmRAvzKa0/JZl1GWHkOjPN0SiCasdF7ak7D/O7s7pa05eTMrEsKVT0XiUxirodcUKxjnbUF5Rx8T6x8ag2SBXLgl2Tskinr6++zTD1ybc5iZ/yI6cU0CGBKByw4K9l9oVwCTbUmNlTqDKE+oX2tUlF+BJNGgApqG0EVwsfNzzn2jsj44k1kgK28uFZnFHu4syjcb4qclPkk2eKkM7fcF4SmfknxIY1B8iCkF2EwSUZrekYsC17D9a2swhLn9wHUOuCL2LuxoUk1Cu49smEKhbyey0OpJu7nYV0nAnMVF2nuegzEHsNzEmgseNaqviAGUvANozkTmKHcl5oy62sBWJLwPEiNWlfh4N9e8Hso8y6vF1ivIdaT8kuoGXhNk0KYg4AFMFSo6d4r0UeR3IAv1peawsWCGvhiBLKegmcF9YSf8EaF2W/+6Sv2P7S9/Ig00sMazg/719/cowLpp4dfH/nCf7b/85Pt9rr8Kj5lV6c+bvaVH8Hw+PTv2OxvHLZ3I0vj0QsUc+KC9fyoy9+8tc20+HHv+Qfe8qe8UXG4udUezM5qgQlRWihYn6iLNdJ4I7nli+CVA45CAguSRNkPrRoFXmIWBG01inixiOJor4QtoP2KX0BBR+aFAAAgAElEQVRDgxIIAkIFa+oOu97uNnKaZCs8iOhFIDrntvyQB6sqCFC0oZBV8STgISPAkw3vjrrO46MNCxXh4oZC11/mNg/Nbwj8SFw4oGPCRVDI/znAlEytue/BNg01IO9p1kRGRfgQR5kHRkVElFNg1OGiKI69LegWhgKmKMqhSOyocWdRMM7c96PmVI/OWz+YvXAYx4wxB1kLWkv6u0GuhcKKy/HQJHF9cT6TL/cdiIbdXgqLhf3Y4Y3BSxxLisp1ubRlU0lpP98bG7W+nn5bW9uw+cUVq29ssRqetVWFEqZ4KfQztDc0ktHBTT/sEDPvYuLPZ4AuBTvj3Ww3zgNdrCIxKEkCJzUNaj0JQsaork6BGwcUCCOCaAKQbd1TguPQWFIgHFCKEcXjzAFnJEgGKciTONrfPVIU6CPlFJDYdNmFnN0su6ZjkFLQuOr1fv0RTaTnFR4iBzvzIUojxORMFL+gsQhii5+rQSNvDJeSiSippoYGMS9AmDDXu7pAzntyHrUOCZIYB+aA7jnhhlZ8HtR8rk/GXUHPkvULQwNKLWtNGupCYTl9mEIu00W9AwWvyIFAs0XLuqCCL88GRAiNQZLNIiba8hnzdSo2QdWR194gcUM03kNybtA2g5ycsxi8kC62R0CCsublNaCmp783BQOCKF6HuW0OVHpTo9ObSyUVDgjcaMRwX5LfCogumAzR60G091WCYKeWSiJrA1mj6KXx0ORY0mKBEh1/n2sBTadGJcEWWrIg5iTzEczUKOjy/qEho71mlcKMo/l5X/ZRkJkkEUIM1tYqCZXkT0Bg+NyiSQetHAkkN9NV0r4JtbUiJCZJkNAtsJ1qadT6nuyMJvZvR/77lonsFLI8fiYwTiQskt/SuvQgMTaDEgS1FG0oOIb9DugkyQhFCcaid0efjY2PqxALypNzgGfitFe5yCvYlfwgPkmYRk9O6vMoQjD/SMQiiwHJK/eJ2bSFxSV77tlndH8k6jwzN9UuuVFsCIw9yGd/8zOD9+Jcw5R4cWnJqdRxngXvFjVGkHDSGPgeIEQYBqCS3jDNsVhIVAG6VJb+PkV2GaEzyKLns2bQW3bEGsW4crlq2UydEh4aRKvrKyqegSJmfggVFczXYjOXe+IzxCpUEIv/TUZ0dvYMSfuhV19XJwQ/48qYiCVCAalc1jzavWe/zS2t2LtXrtoGJu6SP0t7oQpYpdhNmypER7NsL3ZC7XemDXslc1d7e5CAY5y5rt6eLlH0+R3OABK/2BjkPdiXYEmil06RhYFGEgBkPN4SXCeshf179wrlfnf0nh0/elANxKG743b06H41KaL5NSAAId/D+BJPoCPOcwW9xw1ulgpW2liXFNDBQ/ts6M4tFfVBAGPknM02iJVB4Zw19YBiRSYj1CXX2FjfYLdu3dGazmFcHgxQGZ/ZuQcqQjJXWTPsKSRtXT091hyKSDx3GuvdPV3b5y/759TMlJIS1j/xB4VMnhush+HhYfei6Oiw+/fGNed6+vvszt0hXQ+yKO+++66SdxgYd+4MCdnO9cN+AEHK+966dduOHB5QEQspDAxEMUUnMUJGa+jusNYEBdlr166J0dDX26u5CuKTwjBraiO/rmIaMcbo2JiQvmtry7Z3L3IySFLQmK3Y1WvXFWuqCbRatIHDu+25Z56x/MqK4WfW07/L8JMAGAOLlnEBDci6yKazdn9s1JYWZmyrvGGNDRl78uwJs1LeEtk6yXVU0vXW3NFnNWlQfjRsEzY1NSlPGZJzTH3ZC72wkrfl5UU7eeKEik+379yxn/3Yx1UohO3y0h9/VWdbETSkzkez9nZkiAq6f5oQ2juIk9VAd2CFSyo9BLSoGR+YEzxgniFMsYh4pEgu9Ge1qmYsrCE8hNhDxOTTOexsyeiPhqQGzzLGLxEdHZlmjoT0GMpZFQFxKc1yR+vRPADcI1ZrIiEdfeaWCppIS1Yxsgz3QfwRGKRIGkYJRuYGZ0xzS7P2dvYpSbACIAixDv+m6IkptXwbckiILVhza5OVKm5UuZEvaC26XncsgpQl+RObypz7FD8pbILSdakEB3CwlzDPYPCwv2LEWpf1HIa9hLhms1qxTC5jxTySaKamb0dbh5qZiZQ3jGgWMe6xyRWZaxcvXlRDD/nRhvqcnhHFGIBNmzUeo1DcU0ylnAOkp8twCQwk8ABxXFL72MjwsMaW8UK6rrG+0W7fum0pahdVs7/7d8/ZqeMHrK6u1pZmZmzo2i3r6e23jt5+u357yErlqk1OPbCezj6he6/fvGWpLA1tzsaE7dsHi+KitYPy7uuR9NPA4cPaN2go7d+/R2AimonME+YnsqGMIcUj0MvL6wW7PTQsVhnPtrkuK+mnkdvXLVu7ac8/d9pmpmZsZHTKdu49ZBOzK3b5xpBVU1mr1BLrewaGLCzNkEyu3se6tsbmFuetro6CCzFGQo1M5iOsTOS1QGOTjxJv4dEjuZMgS6QGF+d0e7vmEfs7TWmaM4oTKUjVuoSRFypr1BzK0PhPJW1xcdmNkIlLN4kBHTUePcIicj/mVh9sVMBMw+Q2geRltWpnTx6xM8eP28id23bj+k2rSWTt1JmT9p1XXrcTp0/Y7OKKmsY9Pd3ebEnUSKoPKRmyBeYRcR33owL04pLuiRhhZz+yYB7bEZ8qniTmr8vpLMnV17nO/WbJGnIuK0w+xL0QbxPLwGKbeTAj2TPYDo7WdvlOxpH75X35TMaPfaW3u0feIGq8S2++T5+LXr8AVmV88zwHEVCxuiXGFI0v9tYN+U3x/q79r30Jzy7OAjV9/XdZ2zxP4iZXM/CYXo2QIJcbxz9KVcVcK5VwDx5AHDS4ojeR4uvylmWS+JIkrLkxa+fODNr7168FadisHTt2THKoN2/csr7efuvsatP5hzzapUvviG35+OPnLJWs2juX3rMXPnzO6nM1trowK6ZGR2ePzU5Pa6/bdXC/jY0Ma+wHjp+xK2+/Kxm5nXt2WX2QHcZInELtyuKK1VqtHTs1aEPXb1mlSi7RZFev3bT70w9srVCygvIql8dlHA/u67WmuowYqDlipkSNvJPAPWCmvWkJa2nvkvwh7AQ1yHVGuRSgGEjlTTVYXd7WgT//L3vvGSNrlt73PRW7qmN1zuHmnCbe2dk0u8slTZjJpkSsCMsiYNOBsICFYQOyPximIRgmDBgQYNnQB9GCYJoryaBEUaK43OWm4XLSnZtz6r6dc6zuSl1l/P7POX17d2kb628cTy8Wc2/f7qq33vec5zzhH+JzIQ/wOBXWQ1j46nGkUzp7YcmRm0cmtcrlUD/zrIiHxZ1dG+jrsko4F4kvHluQH8TXzuti5c/0OACpIpOMR0w9JU8pZLWasy61I1ZgLmu7paLiPLEJySvyUfkYMXgMDHu8Xi5cOG/nz5/T2kJSUCCWdFZrZHe7qNxMoDmpYODHsRdAbkhBMXhxYGBE0QuMJYCS+3eyn6IsoxgZ9brNzc/bg4eP5MWXzSOpW/FBIwO3YEzOfSVLIM+WLFAK+cZWMZ3IpRkawSamZmffAgDk/fj5MxdO2/DwkPaDywq7oTXrm/fndd2Xxmtl7rUkiumf4NER2O+RyRQ9syR5h8w0frHKwYkJXuex/yS7W60e3F9ySK9p/azg+XAt8gOt1gQC4t8ZWggwBsg2DJTJh8WWDUAm1eIbGzYxcUSxi9yUvP/M2TNiHcG2QxVhCoCK/CBcEtrNtfGZ4DP6Ik2nAHi4THoE1mlYEvIB1XTy4Yx9QpcnptYhXrgpN7WLA3cjKFHPSYMZB5vEnqdAUUFSDbak18EOZo6DIHnOCkQNo4h6P63zzwcWNEAcAKhYTq4TcjT1cAJQl3vI2tY1BWlPcnnuWwQ7sr95fb/WzF/9QYXF5v9PGFsfanP+5v9s0/+52d8/9Vv233/ht+3x7/+slX7/t+zC190H4ie/XF7prQeH2A0/4lFx+DeG7He+9Q37+vE5+93fvGVv/aP/b4OKv/MvfmC/PfGR/ealr9vv/sQF/W37cPrXrfAvg3fFT/uZf/z1PuGDijOd3ZpKS4qBYEbS3tujpFrmfWkQjzk1rzhkKBZJBmka8TNsjosXL9r09AsNMtisbjSdUUBHP5lALQZGmChzaEUEhiPhXWZHOr57e4Gy501fUZ+CYTabmyaZU3O9aS5JHH4O6rqCQUZNR4KnGBY0vdCo04TTzWwVhqEEh4YUMiRKjKIpdpAwkdmw2B77Qt1wfWoeYzKKGVAwzAVBEc16vIHjpsocUjRko3SKBhFBIsn1cw/RW+Vp8XI6LT3pLaS3mMg7i4F7TRIIEjLSL/2A43DbU4PIkVzo66Mn63Q3R7WGoC1zqO1geu7+CVH+5OVQI6f35nmLYi2Uiw9IYnIoJHHorMdnod9HAgTWX2Pf+no6VUBzz1pbOmx5dVOFyB76eiqm8POAFeHFd2zeRjojr8u9ZA0KJS5qn1MaI7uEJqH0oJlaC9kd5KkkmQRdEEkP91ShEARJKRROMDriNdW4F1rENZV9rBU5yGGdRQmucOjGwZyuMbIYlIT7OpbeZcmptC5F9lJaSgOk4GvhEyynLvtgyZvDLa3NWr9IFzmdz6m7oFK4P7xPZLFoyBCkQlQQaPBj0npuyqZtbW1VTRFolPI0kLEyDCQ3HmdYAFI80uClcxgQTzK1C2gN1pmeUQokdFa+E9BgMf6E1kmzrLyHAVaQLpKJWUNFEX4INDWjD8rW1o7Qj1rZSUcmiMbp1KOAXGE9u9lZpEvy3Om/KtGVjAaG6Y4EYmAF8j3qSQrNDjpja1vJFkwx7gXNFf6NJr+juBK2sbGlxkM0EFehF+QweH2Pg4HZADsAvUoQY6GZIoOswD7wAUQ0aHRDsIhOEesg+McQQyVPFhAe8ijZLQb/huaAlMdErKjGDskRCSDXrhgWPFXQtuSBs6bVeAeNk3JTM1F3w+AyUloLnQXb3UUruU0NOJ732sqahr1i2dT21Wjk5xV7JKnhyDzXYS9bc87R5TLTDfuSZ+WDxSDXEcx0EZxmTbhET93SDLT3MQdsk+wDzLDp2TmthWwmp/tO/OP5UlDRzBP1N8UQM6uGDOcNDWAMd1mXXAP30weDLiXAZ+PZ/42vfc1u3rpljx4+1FnmiKbQvAvyIi6t4F4grHcKe/Sj7929J3SWziv0b2myBBM8ebsElg0a52xq5EKgm0sWZm9XiWlkUfA8eB3Q6KwpJazhHlFMMXdDk5YGOp4h5TKoRtcTbseAuc656cU+9ySi4SKjhPMPqrcYBKmkhorEcRoxkenAotor7llvrzMpASJQbHCeaQ2lkra0smonTp21P/nWd2wbzxghozmjU96UUMMWnVY/H2GL8HdnITEeTUiuiuGQzo6ANOI92HM0ytEeRzB4bmZGKEbJnTTnFZ/YVKzDQleXmnignjjzKrveiHrl8kXb2dyyyRfTduncWSH6l5aX7OjRCd0rzGNpqHMPhXhcc5Nv/o1rPfCVkaTFvgavDI4099yvWqG9xa68clFU+6WFRevrHbB0GlBEVsUQzzDfkrc//pN/Y5dfe0366iAjMQokHrIuiGdoe0cmH2sCJDPsNvIscqsnT58qtnGms9YZQoAe1vmWSunZT89MKecC0UpRSx7lOVBVmvOYihObGH5Nv5gx9nZ3b4/dvnNHQ0sMu9999wc2MjwqKZr7D+6ryc7+unPnnp09c0Yx6Mb1G/JkKe3uSjaMZib3bWF+wa6+ddXuP3ioNUsR+d577ymWDg0N6NmihX7qxElbX19VES3vigaeQ64bTw5Y6GwVUKKtHaTvrj19+sImp7h2j09jI8N2/uxZO3Zk3D547z3r7R+yhaUVmVczGDpx8rjOU+49bI/15SWrlHetsx2kY8lGB7otUQVtlrFyPWm7pAL5NuvsG7JiCckLP7MwT16am/PGWmubhi744njDO21Hxsftz3/45/b6m2/aqdNnLJ1vtj/79rftgw+vC7iiZm2TG1JypgjdBjOQYjaROGC4kQPHeKImIMP6INHoppEuH0URyvN0liAN8ooaSuwjHywXJc9HA8BZdS6fwvmkRgCSb7VaQC36QFGyA/Jdc7PHaFrNmaEmhtgM7l8WvSlYh2Ki6suHifwugwqYRnzGGFcpwFl/zvaMuYKbTfJZaODy2cX2C0ARSTy1twcJqB4352Y4SCyGXZXDpwOmpqPHiQcyKK3VNThoL3Qoj9fAem/PtnY2/Z4H6QvOHpounFOcj6DKQcty3QwtGFQNDg3KjNlR3ru2i88QLMFM1jLJtPxhiNXcf2R65OWmBrezAThm79y9Z1OTz3W+MABGukmNVjTIaVqpYcRwyHPuKIvD2mUwy6CSzxVBEUg1CVBhDYM1Al5jc2PdCu2ttjDzwr7ypbespwsvkk1rz+Xszsc37bU3rloqm7dHz6dsa6dkS0tr1lXoFsDn4+s3FZfbOju0ls6cPW83b3osAOl+/foNO3f+rE0+n7RKec9Onzoh3xX8KuLQnUZjZ1engzda2mx5Y8seP3nm5uj4zTXn7fLp4zY/9dQKLSn7/GcuKPZsbJWsnsjbVqluz+YWba+esH0NtrwhkwnIUs4Szu7mVmTq8ja/uGSpFM8/YU3ZZvf/SgNccgkZzig0z2GBSA4SxnOQNiMPJ5YxgFTuozrCQUKcTciNNjVz5nut0dVesM6ODkmQCVyRSFgnDOK9ogytY64ZwTleBrxk4ofqUWvCtwrt4brQ3+dPjdmls2dtEImzhQWxUMaOjtufvfuhvfr6ZZtdWJGEHg1HakOx1U6fsUePHuulNEzcryqfhrGAn4TAQiF+IMEjH6E6hs0+yKPRFkFxrGlQ9DTXWfvkjAz8iHtHjx6zqekXfiYLqOK1cqxJiSdimQapKRYD8QdZLRh87FF+ZmR0WDklZtrRsFtgkgBAYO/BhNrcxPzdJWWlTBoYXlG+WPmUUM0AEN2YlrNeQIeA3I/3Pg4tYkkmZHmQ/BQtPyDdy9Wyy71I5gdwDPK4dcUv/CmymYaMsdHFn5qZttbmVnvzzTf0TKamXkjiCLYNNcL4xITdvnVL+/fShfNmVrWnj+7ab/ytX7O5F0+ssrdjifq+dcLKXFrVPekeGLDHDx/qnDhx6pw9fvRYceb1z33WHt2/Z739A8pp5J+yvWvb61tiRT5/MinpM3SHnk5N29PJadtPMDBF0sZZ/NmUWV9PQbJPbS3NlgVIVEMmsG71ZNrWN3Zten7R0rm8lWvIifoZQDyFbaAhb8YZBQxVuaex7yJmtEB+5KAuNy3wVxg+R9WEWGe5RHf8cmUADb31/boVd8hjODcyYu9SDzAMdjAXzG9qDvdxKyIPS3M3Qe7LgIr9nhfTDU8e1TQMGxr7YrAKICkgZcI6O7uVO3HGiCFhAJZabGkJH759O3v2jA0NDwqQJaAbLJtKTY1/AQ4C+EogwkpZtQRnED48L/1RXIqJaxMIUvEl+kLAaHDmgozb02l7onjeJHlrGUVThyifNw3+1UzWIN9lWzk35JNZrdqNGze0B/jiZ/Dp4/dYQykk8NpaxQAaHRnVfQQYwPqM8Sn2Z7S3pHjBaeRnuQCp9ICCf5UPWlyuTT02mVXvBvlJvIp2tUYAFkT/D2pTSZEGT1lv5tOXcpY57Dt5xkh5xNnt3B9nXCLfhJ9os+4DDG2uIaoITM/M2ZEjEy/zgTAsePuzn7WpySn73vd/EOK7S8xyTTr/AarRP0zD4nc5usjAimtYQI4whHXJbffoZM0CgHHvCu//uCoG1+ogK3kwMgCueI0kFYwgwc065kt9gNC2QOkiylIJsCK52oDelMuasznpSem5hX6VvheknvheCW+/Q+wPZ7bgU7ovf1t5rLG+GibAIu+rzwhbIz3wxo+fWIc27F+FPw7Zb//RN+zvnJ+z/+PrX7e/+QdzP3rRl37Dvvl7/7G9tfSH9ovv/F37DgbVv/8t+52r2/YH/81v2V//Rz/28/YZ+50/+m37+vlV+91//9fsN78XXu7/dlCBX8Wv2zf/6G/bO7ZtG11ttvBTMyp+bBDxl9z2Hx1k/PSf+Ude8hM+qED6aWlx8UBKiYOqu6v7gDXB5gf9QNJDEiL/hlJJ8gpK4JNJIY/4inIHh6VNQEmBFKNhIskYmlpMgEFLBJqVuAZ1NwEUKoNErPxSh89ZBY6O5osEiOaUDtuAQKugsV4u6SB2BLzLKrlvAZhjbzxLL7ZBA9vlnmTCE2UzRKtDvqFm0rANBjpiUeSyrv8epuuxgc7BQrFHg8Unqi5LJSRbpMNKokaOSd6Qlk+FI0s8CfPmuhvy8j5uwCqTMB3qJF7ehIwN22h4dCDP1OAgLAeDX0fBx0m7kt2AaibARUaLGh5VD9wyHQrNJkmyiKKLjEnQRA6G255cBs+AsFEOkEZ+ky2XTcn0i4JrfHTIVpfXhDzZ2Nyxja2iEG11NcUc7RcHJC6JxXUHmS+pxLwMuXwemhZCVIna58wRUf1pHJTLWptuUutyWbwe3weRynWCYmXNQhPlZyN6iteJeoCSSYi+Ezrqg3zXISaE7m1A/agxEH7KGT1u2Kd1F9fcIY8Lv0uBdXOoCIpMG61x0dsdXc2gh+Isou5h7Dhq2aUeNAgLe0pJl/w1TPurOe8m3ej9cm3sVWiEPqChmG9Scw30Hcht3leof5ooxR1/wkHzlw8lVO/erntkNBq2ubkVzF5pXDrlXmgLJH+kYenPlwaxDDeVZKBbTZKCXjt0Rqe/kgxy+ENbR0tde4nnV/VGkDSSzZRcRSYJ+08JQbWqNcDzpCHA+8c1zb+9pPIW1Sz1xNaLQ9JMJXABscD3lQQERGREdUV0BauBmCAzuvAarCXWoxqzjbp/FgrBILMBmkaMk4bTZ6NsCL8nfWhkbzJooBcPKL2RqSB5syC/dPg6PSGEqeD/riZXyuUq3FTa5ciEpP2Rdcw17NqRI+MHBqYLC0uiUzMIUeKpdRQl4BwlHE3eSODQ9lRyJ98YN02m6egFMOiwZivtlrTOK3WKVR84ijnE88+49vTZc2cli4VxpGSQwt7X8LLmlG7uPz/Ls43xgkY4iENiCOgoUaiDp4XrqnrixnUfmTiioRrDdm9auVkaPwPqSA3FJM044m5OA15HdzXcvJ4mZtNLeQ4fVgcJupoXdRo6y9PCPz8FD/eSNcn1g4JXEgmSmsLxAJXlDQ+KbMke2r6QXsRlkOctzd4QzTbRcESzGKkvTNuc/s3AQsihjOuLs65oyFN4xgNTSH1M6Ri8MbxNpWwH1HShUybMrK/FxXkVtol00rZ3d2104rj96z/5U9sE8a376uwEEm3WEpJsPFso+UqQg9zJgam9PGi8iQmTgPuATBPnO9cGapvPowISOUINtCvW1d3tyCakIHaQpHKJMQqKFDIOra02MT5q25ubuodIzVDUlip7GsRyg2mKMrwG3YbMJANUGr6sCy8+Kj7EDuw0DX62d1QgI/GQz2Wtvb3Furt9kJlK8Py2LZ3BNBemVsa2i9uKl5iFCjxtCclb4tejeMIAMuXySsRiTNCj5ix7BYYUMTg2s3kGPEcOP2K0+1gRk2tChXNfZUqcz9mDB4+0106dOiUJND4T59n0zKwGISdOnbCPrl3X66DdfPPmDRseHtG1PXr0yI4cOaJ1eOPGbbtw4ZzuNzIyn7n6hhpZ6Am/9uqrGj6T5129+qZd+/hjxeZjx47Zhx99qIEY954ikcEQg4rVlRXJIUxMjKpohEUbkcNgAQpdsBn3hWjc2iraD9+7Jk8r4sixI6M2MTZq46Mj9vD+PSt09lpre4difyJttri8oMKc+FEtIytStXwWE+Q9a2lO2WuXzlhr1j1RKgxYs3lb39mzwbFjkqABsZrONFlpp6hhDLE519pqt2/f1mCkv6/X6jVYwwWbnZnRcO+L77xjmHqXazX7xj/5p7aysmmNhiPmNNgM8R85DfZ9RL2xj/j8OusCy1dI8CD9Qzz2WBVynyD1JUACZrB6rSYVxH52eyHsYAaXhfBhKeslxNZQTJMn03UgdotNGCQMYjODfbobWMHKciSR6kCUmCf6+3kzEPBRF+cxZqo1R0yyn4kxaj7IC8iBPtwXzlYQ62i205SI7x/PRjX4czntC96TfIGGsiSkMj4IJV9zedEgP8jf1KwVQUwoYRiBkcVIrswzQAaK9S+mJJIRmKCmM9LfJlZMHDuqpjR60OxBsWfJ9aout8dz26CuATgQ0N4AIeI1c000jbiHOtsbdfvhD//8oGnNAIUBrO/rnO0WaQI5SzI2ZPgA7HMGAUhTIk3kQCFqEwdEIImJDOB+ZdfefuuKDQ922eb6guWSCXt4+56du3DZ8p1dduPmHUukmmxvr2a1CshV91YCVS/5TD5/U97u3XuoYSzsiJu37tj5c6fVHGcwe/bMCff4yODR5wxBhiog0x8+fiLD2q29sky6WZxNMOCSSTt/8qg1Kru2ubxkP/szr9rC3IKtrmOG3GK3H01auqXVrKnFNkHVlyueKwU0KSm9AFY0M5Fk3d6xcpV8kea4y9lwrjMozqSTWlNc/+NgvOp5idcOrD38HTAMFxM242hYAX44U+r4KjgymNbZ8OCQ5TJNGnr0Dw5aOUhiApp5MT0VhmuOnHZGZxhI/EhTwHNifobrs3rVMomGnT0xgdiVNSoV+RMB5rj/+JH98INbdunVC7awsmnPnk/axYvnlIsgtwdQ4/79+8oN+MKzZnx8wmZnZ212bl55M88HqU3AE0gGIR80Oz8fUvPgaUjOkwZEUpKBOmfU08dPdO6Sx2DojBwgbGDWtiRDAjiLuBOlljQ8rDkyl30+MTGuM4NYRR5y9NgR3ZfZmbnAxEJG1JuRnPcw67hml0VOKictwpJSnuzych4zvOr2vN5BaORLnNHyXItill4auxxOqMOEYwq/r/y67qwZPCp0vtNjEJ7Nm+ewD9ryWck/Xbx4VuRGUUkAACAASURBVACByalpDQwZXDx7/lwSPuTD7O3lpSU7fuKk3bl9R54beFTs7W7ak4f37W987ZdsZfGFVXa3NSxobWmzzVUYla1iTSwuzNvG5pZdvPKqPC6o0199g/Pzms7Pvv4BNdgTaYajGSvv7EkKCumnWj1hq+ub8pvAowLlAT4njFE8VFqbmyyTqFs2nbTmpoyrEdQbtr1XsfmFNVta25I/Da/DMJaGOfda51Ua2VH2lfd3qMXIwyJKm/js9UZKe3V9fUP3m35HZIlFwKNkoQLLPjKdNaRQozRlpWLJ2tryqj+jgTS5MQeTD27d9FdKDqWqQHhSWIDhlkgpD6tzRuKphoxutSw5PsCifOWaqNXo0zDQRDGhxVrb8WxzFjzXC3gFo+Te3i7r7CrY0NCQ9eDHJ+asDwu4Zq/hYfB5w97lOb2+pj9CXRH7RxEsqgGHADges8nVOOdhhnE+IwMGQAo5KDWYw17wGorzuqEeCCs0qiGwJzkz8OCYejGlQSr3lpqH2p88m/2nflxTk124cEHs/+ZmTOx9iC4JZfongKMCgEEAomrFAFKx58VWl9k8AAHv/VQrZTFtZP4dAG7Ut9RcGhoGlQl6ctzrCFRwkALACTy0ajobGQqQl9A7EuAtC8DHgWnUaTwA7xc5yFjDL3I6sTMc7Ec9gJRqobND+SKvExVFOD9VywfvUc4IMXXli5gRUFIMliD7Tl7t0k3EI2f28/58fp4D53tEL0ffTm6kKx+4RyKX68AQZLNdbSA+Uz4f91uqH2LTul8Rf4jstOizpX5j9DYNDP6IRlSHKQwr2BfwdnmuvC/Pn3MtSh1S26xvbrh8V969qHyY4ozcT8CggrvxGfsH3/kf7DeOl+3B+9+x3/v9j2zS2uzMz/+i/caXTtnA5kf2X/7yb9n/FA2q7TP297712/afnGuyyQ/+jf3Df8zPmxVOvGP/6d96x043zf3kEOP/aVDBJXz1v7bb/+AX7XST2YOfclDxl5po/3gSIWmo12zydz5nn5P21E/7mQ+94Cd8UHGq0CV9T8nWBG1OkMkEWBqYfBEUCGBsQg5khg407fkdNGUvXTovKpKQ/CERYeN4bQWtKil0HlNQNdGUTDrbwJM90jvPSNSsZnpOE1MBzRu60igPzdHYdOT1mY7DqCBxi2gyrjUa3HJNasCEiEAA4hBSwIxBmIYe8k8gWijSgjEoB5S0ADFS2ttVkydqtWvi2pRXIKFAUWMofF5vkIOu8s8nMx2vGmOGqwaYI9+CfqtkXwi6TlknkaBZFem5BGoCX0SEanABAiKgseOK5fpjg06HdkgiPdfzxEMHR6DveYPOqYw+Ifd/IwDTkNa9C1PfOIiK6Jv4nnFQocYosi+ppA30ddvG+oqkTISAXNuynv5BW1pZExW4tE+zzyfukWLoSUaQ6xFVz9G5ET1DoBYjgEYwRqCZjJBwWldB09+9ETwhEyoBRDGHq5rZNa3DUydPKAHQIUXigzSO0M6u8ehF9+HhhNMqJcF0yDzYE5aUimcl34H2591YL9wl/UAxfMism99T2hbkgsLCOTiMI9pRMlPItLQwQU9KS56/M5iRtIoOdr/el88Cr0CXSSE55GcwF6aYZ32RgJDoyMh4fdNlzGCkcO2gNEJTRIg6UMyVsmSS2PPRD4TXUeKrgsbXJDRVhoT8vnxYAgJftETJZTn6ggOe4on3xhQ1olBZZ5hf8p7sNxVSOvQZOCXUpHO2QCOgMtx8Omp8ujyTGz3L0E+aqZ5Q8nwd2duqQs69IVy+jeeMVEOkdPLeND00wAyoOdZKRIBJBg7zr61tDW6VyAZZAVA8cQARkSVedPlQyenuPgTxRMnpuyomNSTyQZES+bI3s2iYs1ji3nR9bG9C8Q8adATpLbTDachG9oHLeLmoKshRklGKG5pP2VzakeSlkprAmPJJBmzfqbExDqDzzHvyDNwvyGWnkE2Q+mzQOve14P42fBbQpqXdsrNAKhXr7O4UO4jnnRGaq25DA30qFlvb20T/ju/J54oybj6Ybdj25pbWrFOKoWJTpKSEtHJTWLBnLiUoY8ngo8P1C4WcQU6pqD2MHi17APS6WA9Bm5kflIQJKJosZwEG1e4tgYme1g5sGBgiops74qmz0KXGM8k4hcRehfMA1JQb3PLs+d3YjGZQqDiNhJOGWVFWC/3+HW9oJ9k3xCOagAzAGGZgTBzWRDCllhxbGDzyPqy/uZlZSUqADCSRZQ8To2CueOM4abs7OzYxMmLtQaIIPwKQpxU8nqpVSe/88Te/rSYSVHbWGC8ibyMt6X3LNKUlF6eig/eW1ATGtY4ywwsIdgiNQ8XKhKnhoiG9hmwuM4DUheTUggwF/wZzhfUKgh2ksmImCXs2Y73d3XqdEgjS4OlDsUVhw9pFexnPBrbe0tKK9p3QzvKzchmM6el56+hoUVMXxCXsEg2x6iaJiJOnj9r01KSjCvcASlA0JzWo8EYPQ6OybWxjco5xI6jFsgbhvT19bnKeDZ5LYl1xrjl6XLIC+/uSruru7RJins/C+l5ZWrbe7i5rb+8IFPaqbe1suHSBikxAHwynknrGsDrFEhLAYl/PmZjLOReH8zTjBwaH5Mnx4UfXJGtBnnXv3n07d+6sfueja7ftM1dflVb/5PPndvXqVSGMNzc27My5c2q6cC9OnT5lH177yE3bYQKA+mI/0OwMUnWSVJMkgDfRiQld3W0a0NHs3CnSAEzb/fsPbXVlXRIaI8ODdvzIEQ3ANlbXxNa6ePGSZXKssX177/2/UKHumv/egE7YvtUF3ti30aF+u3j6hIZh/Bza89V6wiqJjHUNjFoj0WTJNBJfsA9B4KWFPGYI8eF779ni3Jw+a2cBvf6qhkPHT56w19+6Knk5vCK++SffsUbDpYUiE1OgGjXGYgHuOS/fo9GnPQmyPwyu4zntAJPDjNqXspIwL5ChIjY9ffJMz9f15Bn2wtbjv6Ciq2JU0BziPRge8BzY3/J8C5rxL/Xc95UTxXPKZZuCPGookg+lEjpjWEujw8MHmuUCs1SrNjo2Zi+mprTexeCjwV6tak0gzeWNQm8oEM+4Nhh0DhpwzzCaGcRkSc7JfwL5qJLOKm+uefOT2CtvCDVWvfFQNxoIIFFrAjbwf75Ay1Mr0OTZ2th0QEKioWY3jdr+oUHJ5AilSpzCCDzbZB34aOzsCMkIm4KY6nmX1yc6r3mWsEAb7knF/f3jf/WvxWbijIHtxDVpCJryeoBzEc8nyXmGegA5C62bmjd3PMdGTszPyEvnz9vczAubmZq1X/7FL9ipE6O2X9m27bVVe3z3oR05dsI6+gbszv3HYlSsr29bob1LiOHoQ4VeP58llc7Zo0fPdOYz3GdAceHCWXv4ALmZmh09Mm7dnZ22sDBnLfm8zc0s2cmTyObV7NbtO3bh0iXbrVTt+o27ntclk1Zoydu5E8dseXbKmpJVe+dzV2xmetZW1nYsneuwuZVNW9rctQYSTLm8bWxtOUmWPDh4/dGYPHn6lC0szts87IYMA2QkNFrE7CS+oS9PLocHBbkRjMj2QiHo4nuTke/TmF+Yn9eZoH3AOR9ybCTFXIqxSYMK2BnEDgG0yDGDtxnrnHODRlTMtdTQ+gk2he9ghjpCumd8IN+UbNibr1yw/XLZntx9bD1dbXbpyhVLNTXZ3fsPrVipWqWRsMkXc3bs6LgarIB8Ll+5bN/8028pNrJvya0Y1sMMnp6d13mnvV6u6BnCVoPxNjs/54NtMRqRd3G0NANCENfE4ukX06q9BNY4csReTM/YxiY+PtF/z2vhg1wvsEmFwN7HjL4gRsWjRw9dInW/asePHxO4hSG2Gncl92SJsiqME8ZGRzSEARyFBA45h7M3fDDq/osO6GN/OPimfgAa85zZ42n0mVT97IXSQV4uJolqd88Rq/uhHlbTFy8A19MFcgS5G0+jN15/VRJij59OW6GTQcXrYljACMIniTMO4ObxY8ft9p27GnB+8YuftfLett27fc9+9d/9stVKW7a7tW7ZVMLa2wq2vLikHAawCNJa5Lsnz5+3B3fvakh28ZVX7db16/I1AzTBtWFY39vbL1sygAHpDAO6fdveK1sqkxejgoE7YA0Af6lk3boKbWa1spX3ivIHaFZvImfVhtnU9IKtbRVtr7JvKeKvQJfuN+NDVfeTpHYZHBgQOEho+hCLGfLBNCZ/7O7pFuiA5jFxi3xXYDZJTSH7WxXzO9amYvrp0Xg9s8egogWJKpdmxoMMbxpiY6yVyMfEzi4iOZRVD4czAkZFe2uzzrUEhtcpNwiuJ9ivDC2QTKKfwoDdWTOVclV/x3dtaGgw1N1l9W54TwHHSvgrdtvRI0dtcHhYcpX8EsMbrk+N/X0HxO5XYCn6GUtOx97k3uh6kbMKPp8uRQu4xXsm1EPsRdWvSHxK+qjmfSMBMF0GCYkluA7Eq2iK7IBDV8Pg/l+79rFYbwICFwqWb2vRkDPu1wjumxgf033gzKHWj4oQYsYEtqJYKAAog+oC+5Y8a5faNbAJOI8BBykWBK8KHik9EslrMSwFnFCtCazMF/kmOQixXexy1VaALzy/lboIjEj5RPqzpH7wfhy339eD2iXqPbo/DV/q4aGaINkwj/Vx4E8OwRAJUAm+QlwP8p3+uUKtQK4v2TMfdkWAn2KK8lTuFZ6cyH75YDrW+C57zBnkvQsHzwJuBjSCsgw+cqGnJ2lHvx5+R4O54Pkacz+/F/HcCL2a0F+KvTVJ4gZQo6TsVeu4fLXn9niQuZyxA3Ed2KUeB+xbBkRIYn1yBhXcsCH72n/7X9h/9auv2ekuT6hKW6v24Jv/0P7D/+yf2Y2Dtlf8w0/+vJW37cFH37G//9/9Xftfbv7YL/y/DSrM7J3/8Rv2h78+YZM/1aDCzbK/tvu/W+Yrf+8nrvLlN4Kp9trvWtu//b+Gb/+0nzn82id8UHGmq0dNvMiCoJHEYcSix7ALIzwSIuhFJFEEbQLF9IwnQWzO4aEhNRgpUjRaADlGA393V9rIHGS8Fpq2OgwxMxKqi0LemQTZNJNipoZMpGEV7BwUOhQKHEJswsikiAMDdOxA7EAfjsUimzYMrAPyxZHOPnUm+cWkygczMtGWMVraUW4cwsFgCFNIGuJMyIvl3QMUB0FO09JgnCd9+K0doYhd+5NmhgddocqDKTUSU45ic4MnT9w8aZQevXQbXcqEQldJVpA9Uh6gZM0bmjTjKKY16SVZCVImcVCkJmtI7iIqCCYJz5PJdtRBJ+hxf0EcExi9oeKIY9HgZBQdgixDH5quwXQvJvFK6PkRgqbuKUluiw0N9Nj83Kx0TkHGJkF/lau2T+OmKS3ddJI7Rz+/NE7nz9GTxBkKnjhTdLI+IrJCg6RMVusuDr84kBiaUWRKgosDBf34BtTGHWmS4q+iiX9AVPjk3FHjfkC5H4XYBQE14SbOjq5SE1SNrzDMQB4MFkVAKHrx73ROzacCQsNzuSDxFJ6nUIHh3vFzHEzSLA4FlEyWM2lR5dWkDghUtGAZgHhzNbBegp8I76HBYkgeY0NUSKf6vpDuIBTlNRDYGdJORzMec06YGM3Nar6SmKnRugdiuVXPmPERRYsGa83IQdWV9HLgs4Z0YO/vq/HN53HUlGv3c2+IByAnQWFgwvraa69Kegn9Z2TnFpaWJE8Sm6rEDTWsD5pB0MRLYoaw9jGRpXGGCTiGu2vrq/o7a5zYJnNeikrtGU+quT4xDSQ7RWLp6yuiXGMzip911li7D2XKZe2fQqEz+G80QiPWGTnch4g88mbMnlCV0j0NEgjEVuIpe1gm46WyGry+skLDKhR0oLX7ertsY2NbWqtCJMVGDlTeoOFbqdVtoL9Xa5v33caMLOvrmIJDhusNk8Yscc6RnsjGNUv6D9mI5dUVSycdlSddzeAdwyoDccm6Il4osQwG6DKYPjBQ9qEQRb/u9Z4XC1XufS6rpmpne7tQmRQuxe1taei3FdptZW1VyaTLa5VdVjAkgPK8CINgkl6GDJjgMvBEMoT7qXsffDiESKmSRNPoRmKsSbGaOCGJLvZp8AbiuUviBMPxWk2oTDWJoTQHmR8xiQKrRb5FQXuX74Gm0ftLzxV5qx0Vp6xzDUwkd+FyQfyfZ53DjDaYz3Ke8lx57jQbOANpplYqsNaS1tbWITnE5uYm29jCWJuzLKXBDvsumsVzrb7vahpO8DloTMVmpDRVkTSplPRMWrgn2zvW1+mMBL4Y6lRgbUh+4oj96Z9919YAK6ho2IfcrmvLMFxOu740cYC9KO+boCHLOqRJy14Gvc61SdKlJciZaUDng2Qk4Wh28u8MEJjIlDEDJ2bImL5h6xubyh92tjf0DBk0w1BB9ujc6dNqTFHs4yvBunk2OW3jY8MaZK5vbAlIwLMQxVsmjo74ornJtfHseY7E2ZQYNrAVjtvTJ4/dVC+BhxPxoi5tZNYSn1+IwzyMGXR9YaW4ySlDC+In8YkmLGvCG5UYRmJmWlZDkYaPmvjIQQTgRKrhPlEwRuSRsrQoA1OBKIIc3eTkpD4DMgA3bt5UTgZjAq1thvZQ6JeWFnWuw3pgINHT26cGxZ//8Ic2Pjahz/r46VObGJ8Q+vrR44d2+tQZoTennk/blSuXbHZ23ja3Nuztz7xlT5490748ceq03bh1Q0VhZL9yHuDzQeHE/cf8kbMKFD75EHthZNQd5SjeYQrRiwKV+/zZlJDdSEmdO3VCwALyJYp40Maj40PWVmixD699YHfuPrO+/nY1NNeXi3q95pwsFKy3O2dHRobslSsX6T1KyiGVbbKZ5TXr7BuxSj1jyVQu+OCUBFygActeeP+99+zurdtC4zPcb2tvcTCHmX3hS5+3rp4uDU7+4A/+2B48eKZmOB/KUcHhfA8eV+xxPetgaI1mNzEzMvj4L2vjcBGr84Ice7eo+I7sI3Er+rZwHdzvqB3Pno5GmSqgNTh1wEmUcFVMCuxe7n80rpbOcvBYi95Z3EcVxLAgA7tPEqyhuQ5KmnszNTWlZgUxauLIEQ3VVpBVCwbjLo+QtwJMmEr5QLNZBqKhWcl7iZmca/ImCX/fcfkk1jHXiu8MGtouSYepe1H7F8kgzhXiLhJ7DMM4N7kfyIZxRq+vrupaY27amm/WgAImyObOlr362ms6j4g9SD/VAbUEM3LuzcjoiMyoOUPFpJY+dVKIVEdxwpTDF6Vd6Pd/+o1/on1K/MMDhZjDMyE1g8nHfcIPgkEf+4VGspDxQ0O2tbMlxhKfg4E4MiWgq0+dOG6Jes1ePJ+2v/arX7H2lrRlUzVLNxq2PLtggyNjZpmcPX0xa7fvPLIX06v25uuvqPnp9VlFBq/ounf3Dtq9uw+so1BQnvLoyRM7f+6sPX/2XB4VQ0P91tfTY3PzM2qGry6t2KlTp90XBimQZNq2dkv29PkLxTkaXIXWdnvrlXN2/f2/sM7WjH326gWbnZ6zRDpvq5t7trZTsa1y3XIdnbYFyINdorzRATv42LC/xo+MG95BzydfmCUzatCmU00621gHgGJr1ZJRh3F/l1fws2gOyFxnwzJYpf6cm5uVpKGAboGBzmvvVd1MGx8ghusDvYMatmxtbquZy890Mvje3VHsjvm/pMkOSRD9eLMhnaBeQyrHa55s0uznvvxZ625vtTvXr9uL58vWWmizixdPW0tHu+2UavaD9z7S88cvjppyc2PLXr/6pn33u9/RnmTvk8MysF5cWlJOpNwrDCo4J0ZHRuQttLKy7JIqNKwCwyT6DTKoIN/jTMykfGA+PDys3+P88cFBkw+CAjveh5rR29DR3gBZWKcwPljTnJ+w9YjrS4tLvh4knxj8ueRBVtcwQzKAu0UzcoXgfSNGLD48YWAh1YDQJOT75G8HtWpgxTjpKSScwQfIfepcUpKFwmcQGw1LktjETnEtJgk48uBGrWyJetWuXDlvzyYn5afS29Nur776qjyJ5mcZIB1VjQ+jAhko9i1n7ltXr1qlvGP379yyX/mlnzHb37Wd9WVroZGYTItJCTgh09FmLx490po69+oVe3j3vmLw2QsX7db1j5Xz9PcPqplNPl/o7JbfzI0bN62trcuqtYQ9eT5lxVLFqgDdLCFWADFufGzIPv/2m9bZ0WYzU89tZvq5zoP2joJl86326OmUbRfLlsgSt2qGwgQSqVw/9c/K6kqkpmgQBjBFktoMpAoFgVUFqhRLxMGobFueD8+J2K66DQAODLqgr3/AjMHfdLeooUGjtm9dXW2Se1JeSWNfksquVCC5VEBlDPAZVDRltc53lFenraO12Yqb2xqgUudSh6Jokcx4Tu65EAbY1Pdu7q1h+F7FsumEpK2o/8h/kY/b3SvKcwkZS9Yesl7IuiJzDjNPoEcpTiDduGO5rNc47K/oA8nrSAo9k1H9Qf5Gjc19Yo0qh6RJLpZQRgDeYOqn+EOdJH/XBuBFamcARpiWu3Qjubz32Nr0npw9H1/7WGAdYtHA2Kg+E35o8uQMDXRqLPa3mLmJKKHtPYXIfOG5RjBjlGt0IJWz7ZWPwh5Bmgo/paSzJHi25PaShySpgq285SoLnO+8ZjR7pj6QMblMnWFHAsaDbUx9BAPR5Z+Qez1gV6oH5pFVyhfyenBfEj6A+214f8wHR+Rw3oMhHyoWtwQWJEeHEcf3yLeoZbl27qcGMGHooNeVeoLnOnwfYB9ndexZHI7z8uBR/8mvwVl27vlyAJ4NSgd8dleLccAl90F9RDmzOz6Z/5N3qocUQInx2YR/duBfALxGz0o+XxxaUHu8jHvUgA7K9PqmphzwE8Ko+PEj99O////5DjCoIEE70OwTNbBLAXlmekYNBx9UFFWE0KxkQ6yu+sHGzxFAIxuATYROsSRrai7HEqUOVGDp4HKpGhl4h0Yb25ffkcRToHG5gbE3fGW8WKuFZjXNH590EhBBgOITwbVoI6uh6YMA0VJFqffGvZreKirdt0IUXhrE0LnZ7GU35Ob3CIKgrDJNWWttb7UtzIODrp1MawJLg/cleYva9AQx+VMkXfMzfoEmkpGyvhG0BQOrJA5SuNaIHiEwRwNBhhcRleuIOS9KZKwGajhMuGVKTvPbo++BlE9kxIj6FjwBKJwwzItBmM/kGq0UvXtuGBykn2IDN/6s06vj/Ns/IX9HhxYUfKE9b8056LZuXNvU1CzN6SRamDQL0YOs815Zq5S9eSiZmkDbFeKGhJamOw2kpNODxWpovJyQ0yRRoE5501ZoShC7afcvkMmuJYWuI4FZkenervX19inZAoGtZJgmLA1QCuyQvEfDZCHTA/LIP2c8RH1oI1Rx8NNwSqzgy25MzUDDqT4H90iT+/Cekc4suqkog/Fe+n81aKGr02ioOAe1TrNdzxMjsMAEiabnQpdLTsWTANYoer/h3dWk5ppkWqlDdl/JgaP2A7U2l1Nhy2tgJMy6gw3EZdMobBb9NKsE7IUo4G54B6KP4SN7UIyoIP8CksIRB/45eA2aCazpE8eO2507bm6HX4ZM/FrcbIxEz4dxbrTp6Bl0bJ2iTNNXdE+hJoNvBxrmrS1aR9wrmpQaRgSUQ/QQkS+JtghFlqNQI9VfgyuGi2FNkwS6tJMPslybnPVpQtSAfov+D/wMcYO1p2a7rhU2jzeUuE49jYSpQYlZKnFSsj8heeFnpOuKdmmtYT3dBdHJI/md5UWSHptlJLk8DwoOmqVowotGH5I6dGwpqEiUhYKG3p1vOvDZoWgSA01IeGdeSA6AJFOMBpJ2Yq7LhanQxEw7eAL5nkC6wXWTubHE8WTDJZRAL1Mggw6kQ4kZaUtT1ppzOesfHFCzhmfuvwcrzyUdJAeSZL2X1UwiSY3mcOw7kjOh01nDQU+UoWfcHzxDzh8hx4IeKxR6GZ+JAZVWgstwV+ge/Ao6OtTE5nxyhApx3BN3nrvOFiWtScNEzZ+n/0/mhMSOoCuNF5BL96Gpq92sdc33OFM5F/mzfGcSDTdrw1gb6nQRf6eCGio8byRw0Ot2bwvidGDrBcM7eTIhAYe5d86bVR5zKCZ86ISRNEhbfdXr1pFvtpZ01rIqBBggN2w/UbeNnW0bHT9if/bddyX91JARJu+HDnxGg0oNzaTJzr3PWlMmZ50d7coFkGdC2klGfBimU0Swh5BNCf4sGtrRZAm6vww1nIrvyGkK7cWlFcVraVdLM9aNt8+eOSuU4eTTZ3bx4gWxQ6amJqVJjK46aEFQzuxrminyOQn+FLwPZzVnH+uC50yRwd6E/o9RJUO5n/3ZL9vDB/dF4QcdXSyWLNvULLScQALlPUe0wzLBvyOZUmOfzwXy1YdnLskW1xufQRIfiYQKJMWSSlnrjZjRjvcMORHotW2kJTKSiKFIdhaGS8M8fvxYg1z0mZGtYI3iEwYKr6ur04aHBu3hw/vW0VGw4aFhu3X7tuQeQHIja0TRzrUx7MHTglUife98XjEP1sL4GChmEJ1e7InWH5h3Dx8/lsG42DBd3TY/NyfD2831de3F4eFBxfc5NW7d6Lm13SVB5GuTbxXikOL27u07trm5Y8MDvXZsYtyqpZJtrK8JgMAawoy2pT0njeZHTx6rkdHX32+JRlKoS6RX0ApH0x8YRUcrrJiSmEeSTLSUPZtbteUN/IBarbOrV7EQZHwjjalr3r79p39qG2vrdnRiwlYY8GQy8k3Z2d22sSNjdvb8WQ04nj2bs//zn/3L4D/k8ph8Ea9YY8p1w9CW8w5Wi7Ov3J+Hhj3PnPwy+lbw+84idcSrCubgIeHrxqUYJbkIKjUMIA7ALkEnOko/RNNHxW2MODUYAtXPfc/7gJbcSmhLP5OiwaUjY10+Lho4SgZUMpsun6BhGWbw2zRoPDeJrF72Kc+dVJsziHw9emUAWmBIznrq6uy01VWk/hhykzf4eQYDi0a4I9XxeXHZK+4PAwvALjR6+VxRo5/PdhcCEQAAIABJREFUxKADFDcG8HjNiIVB7hrYJU+fPbVBBgM0TpMJm5mb1X0mJwQ8hEQJjV0+y9iRCcWfrp7uIJ/hQ2bloUiKbG+7yTReOz099r3vfl/NJe43zVnpjpdKdvbsOb0GDAnkPKbn5qy9tU0xH5AD57DuYSphe7s7yk15bdZ+W3OL9XR12Nb6sn31Zz5v2XTNrFa09nzeNpbWxHYr7Zvde/zMpmcXbXVt106fPKnYjDQqcoDL6ys6pwYGR+3m7btibTEofvjoiZ0/f8Y+vnbLck1JyUBxtsNW04BNzUuPSwABiJ+Mcm7fua91BCPhtcsX7cTYsL3/7ndtd3PHvvLFCzY/tyCPikSmxV4srNlePWn5zm5rUFPAMNp1Y+y0Bto+0MefYmltVajwRoK6hRzDfUt8P9D2qytesfbkIYEROjElyKjRAD1z5owtzM1pf4j1qVqhbJkmDLWTXk+mU7a1vqF8E/FC6leYcDxrJFowV2cALOnYwJhSDnIIqHW4T4ARMr5DyWTD0tIcb9iX3r5iE8ND1pLL2dTTZzY/v2i51hZ7+OipnbxwwW7df6p6g0FurFOQI7t27bpys82tHckXjoyOCnCyjN+a9nBe7IuBvl7FZUCC5HlO/3bFA5fldF9IDK8Vr54+s2YkkpNJO3rkiM3NLUj2TfsYsBklcfh8kVHMHnDwhjNu+/v7Ze4e65vRsRH3Hlrb0Pkq9i+5Y1AkyOeaBFahES429X79gOFC/i6/AxrLIa+MsZC4Q52h+KQ82z+eKpjQ3ItNbg03hDp2RhjNPzFq046KriMPo7zM3wtz5lSiLn+HixfO2J2797VvBgZ67Py58/JtWphfsmNHJ5SzAHRDSpFhHrHtypXLVtrdtsmnD+3f+eWftb2dNdtZX7GeDkA3WT1n6p2egQF78fy55MZOnT9jDx8+1Fo8e+WK3fnwmuILXiE85+3injXlm230yFG7e/ueZbMtZskmu3bjlq2sb1mpWrdkkHSFlZJJmr31xiW7fPmCdbTlBSycn34hiSZYFC9mF60oGSUYvciGIvNb0D0VCEcSOw0xKlDFkNQWErop+hztel5ivQTJYZftRKLJvfr4M3tK2X0A6MnMN0jpqPcCqK1WtWq5bJ2dHbZP7A6+oAmdU76DeG9AMcrny1VJlkn6iVrcgvQT0lACZAVwSZODJjkPcvms2CIM5njKMI+VGwVpVdaW+5DhP1MITO99H3KWygJMEUMAdJBLkO/ByGXwCPAtm8rqtb3PAuoe1qyf4RpCh8EYtQKvqWZ9aFLDeOTM1jAiACzpVxBXGARQz/KzfG6XLArsvFD7sc8jo4s1pX5EvWGD+NZsbQnUMzgwqHutegTWUBjgiZGPVBLnOkwCqWZwBnN++fCRfcb7k5dHqWvyUq/3/Gc4gyWbp4EvgAzvvaivEfaj6qJQD8cBp/etQlfs0B6Wb6aGFMSokONQwET5NsV6z4G8HncwFv0IB+V5r4yzlT3UUejQOiIHd/aDe3qyTleXVyRxyvOXCoSUQiLb1a8vDgCoechHDytoxOEIr3/4z/4+XudyD136nf6Ym2pzP92Y3YetAlQE/zKAa+T18qsNm0DswhjjDitiSAYeoBom8oBj3VeXn9UAHslR1R8vZfL0fnkHW9J7/XRQcfik/vTPn4g7cLa71+Yw7Qq67ASgTqb0bPrVVZfgkHyNS0yQ7FKsQHGkaGbDjI+PeeALZlyRJkiQYBMREJnYs/lIuji8tfmiySbfC4Y7tD6EIAGxXXMUslPCXhqkca0EYCbJFEBoaoOsjY1LIeWDRp0frI5+FwrtQLPOD27FCMy+RDdLafJ/gEAmWIWGHU0cJEpohHS0F6S/zL2J033RI9HGbkZqo6JmVUSLKKgH9oTTyzzwioYW0CYy8gnXrOZ1GLY4o8EHQi5r4+iVODjgeVDgSP6jWnH5EZlLO8XNke00RRxtEilukmqQka8nGFyrGAshaEbqfWyGxsGQB/CXptqHN4GKOSWOJkZFtbxnvT2dQiIwqGjK50VnBkJZ5dkrAHMwhgNODX4fePh3fIAQ308IeBrEogU70iiimbXWQuOdhojkuEJDcm9nV8Ux94LGFxIfFG4kpCrW0dYPaFUNGkBBB4Nm7jmJhk/4w/cPSRuJMaPmpaOo1VhQMhNlonRGvRxUBDS3PCoO6H9hZhbkSRxVxJonEfOD+IBJI8kiGrQvTbyl7y6DMepwH2IpYVAT03X4JWlD8ZbxgZxYM/J38MEGXzR9aNq63I/rTaugRit+c936e/vU+KKpRkOqUivrPmF2JRkc1m/DG3O8JglwV3dByAYvOdxHhWSFC6BgBxFCMkhjHdRjlPQhcdHnYDGFMYs35N1PwKXqfKrjQxKX2XHtcCRoXBrMKZJ+b4QAESvCdXUdLe2IHH7Xzdz8/dwg7FCzvFxRE5B1JS3qbMYp9xSJQYufWEHTsqtAQ4Y9x2BGu12JH79zwJopVa1QaFOTLpFw/X99DrEvvGklVA8sg5wzAjTMC5+dz0H8ldm1gqlTZ9X4CibNSoxCYzj6zsjPYW9PdFlixosX004J5nVD84o4qmaWGmQMLijIDxzA3BR1bV0xQ5IdosrEoY8Pc5CxWFtd9wSZfVNH+7/JCu3tdvmC0+KRMZBXUNhXrPeIYuH7NB78DEGOqSSkCoMzzhBpv4OkkTxWWbHAY1tAQoUhCuuK7zNoEMKFYC9Dc/95rfcUTBCnDTOBEWMhSBJI3xX/jSb3GKC5rsFCGLa7n0fwExBF2FFjIIYpcIjF0Mxp4FM0xkF0HNC7NnxADWEQR3HK/agG2SdGNJLKIhHGt4aRDaMC37dcK58FxC/3wjVnfQAixgyNPAyxM2lpghdZu/kmaQC3ZvOWZo0lkloTIEBLtYpt4VExNm7f/t73Jf2Uwhx+31liFEacZaDk2jrwrGq1lrZWDS8pkihmOQdgenAWuuZvXcMLkIF8/lLIFbiHraDYhULz/QswAITiyvqmYorOvUzW9f/rPgg7d/as7unzp8/t4oXztrG+qmb50WNHXUtfUmWwoDCNd415zgKZ9jY1CTHJHokFFLtGXiLJhC0vLluh0GL/1s991d599/t+3oIFRjM64VIAkoMRW4nC32XYaECh7c79zjU1e4MJ6RhiDrEiINPoyvK5iYNRM5jGIlGHwR1odBWH8tnyWMaz0cAvMKmQmKHp297RYQsL81pzoEGRJ+ootIudgFwHbFaM2+cW5oWSFIiBU4X8KPhoSCogaVbcK0oShdyFfGJkaEhsNNY3TRs8g4iX6NyjFd9WKAiRKGQ86E0kxvhMGig1aZDCsxB7te7MOcnhkU/WHHlIM+3J46eSwGprabFjE2O2T8OAIRuoPIZ2abO+gV5LN6Uk23P71h3FKp5LpcQwri4N653Nopo5X/3y29bZTmMKUEjD0k0tNrO0YQ+eTlsy3Wqd3f1ikXHG4cfCOgC5yD0eGxmRPwBrmD2Tb3Hm2Zlzp214ZAR3bvvH/9vvCe3Ms4gxNbIOaabzu7xmLCZjs0LSpcgjBLPJmGdxxkl6EtRiMCSlGSuPIFCKOku9sejAHQcvELe0Zxh8woQVe4J74Ya0nK2gC4mt/LtYDHg5yITS2TlChubyei8GUexZUhVJLHCuAYbJg9bL6AwFmSuph9C04nOzlz2+ev7FZ8HjhRQmnkfkC5JtBETQ0uJsSLS15ZfWIkqMxvfUGLAqkp6PRzQ1CEkNHTFDfzFtC6C5kWILoB/uBfndZ66+pRjPPRHoKJzL5HkYCcOUOHr8mOE/R8OrJZdX3EyKXedeR7wmw1lnc7qkjDcNHBVMvt3d1SOpUZ7zzRs3PDcMDESeHTFiYKDf+vsHhJp9+OCB7q8DXBiO5cRuQmoslQH5uSNqt5qsALCQtshlbHeraL/0C5+3of6CZbIN211fs521LevqGbB0S7t9+PEtyzW32+4uzwTwVyPkvBXLt7Y4WtQydufOPRsaHtbnvnv3kV26dNZufHzLOjrydvzYUZeQyaZtbXVVOWG+qVnXwxB0bHzcqg0fVPBU+N+rl89bV0vO5qee28byqn3pC0j/btnDB9M2PDFhz+dXbHFjx1q7+6wkfXH3lIMlo0YV6NlK2QaHB8VuYSBNfMVMG2CGJF+VTzCNbwjdThynSRf9uqIcB39ncP3s6VPFI+0nzj5p4HOWko/sS4pye2NLOSz1J7nFNoC6XJNG94BbqIMZpEnCOPhzee79Ulr1oN4Ra5lcu2oZ6spEw968ctb2y1VrzqTt4rkzVtzds0dPn9q9+0+srbvL1otIBRZtfGzUdnQv0nbi5En74Xvv+d6vNwQQ6u/vk5H22uaGYgBMmI21TQ2AB/r7ZfxMg1q5YqyV1ERkKzWUV3G2IR0D040YgJTR0+fPXDqY4T25iMAwjspVLRqGBxE0hYpBb2+fPXn8WOsfYMqJk8dsdX1dZvfcGmfgU7uyY52tyEBlfX1N1+O+d17rvmQVO6I8Iqs5M4kJPON4H2JzLoLhHHnstZBAgkGqRaA0DVGrMov2yjFITCVcYhWPCryM+ns77NLFc3b95m1bXlm30dEh93m6e0/DBvoY3EbuB2fefRgRDCouX7LS3rY8Kr72a79g5eKGbawsWHszYLy8rSyuWGdXtzU1N9uzx480gBuZGLN7D+4rjl15+2178vEN5U8TR48JAFrZb1h7oct6+gbs0eOnlsk0y2/m3b/4wHbL+1aBPS82PiwCGugpGx3sseNHx+zo0XFr72iVvxMI97nFZbv/6Kmtbe6aAfyrIQcDQDIhpQqeiWR9K16vSX0BaUrJADqiP0ob8Xd+LzZpiffKMQ/YeQERLl86B2ypFyPZ131dK4OK7s6CpBUBEAL+kMQXHhCp5AH4UnUR4NVgpo0yhjwqiM97ZQ38OBPw3GHoSNZA3KaO4Bpp4LO2AToymOHR5/OcPXGICCgzIelj6h0/E7jGqvIi8gwGpgBLjp84ZmlYwihYGIMw77FwjyQJWPI8kt+R/6K8V4p6z33znhF5FYwEV2Fw6aFYfzEwlbeBwLYwkL3xDZOL3JO/UyNwfeSSXKtUISS1WLNsnvWRssHBIV0HQ1V8Y3muDFUUD8OQ0WUlqV1/VBXCKxNn7HvN5tA31TtBktF7EsGDQ30OYqGfz7HBr38PgKI4yMVXT12KUIsLsBX6EbHXJekv9bPCcCVIKzubgRregT2KG5I+YmDk69EHJN5F8MGZ9+tghZFLqw5pbtY9ac636HMBMiIv4Xdi3nU4nrD2eLYa9Bz4xQYZrzAciP0FlzSG9R4krwGgyHOnai052ChuKC/Z5eATqr5jAKBoUBHuR8Dy+akS5QXD1IL1yvc0bApAGAe/+nXFPgZ/Jn/TswyeWjwnztVPBxWfiNb8px/i8B0439MvynJs3FF0ChEog80FFbggm5hOknRTCFOgwMLwYi0jeihJNzIHBBcm1lHDlwYPG4iiiWBPIU4DTehaIYbd9I4GHNvQkeBxAuxNXp/eegGlhCmg7gkeagjKeM2bOIeb+XFTUyTIdCYmR6FR6s37QHcVNdGbbRSrHe0d4UBPC4VatX01VaQJnWtWAOLQFOWwWLTOzi4V9l5cEVjQ/s+FQ8fZF1EXNxZwnjBQfFKkebM7oiw1UAlGT+iVE9wx7lJzA6mdoKOfznhjkwKVQhLEGZ9DpqSwQ/AlCPI9NJdohvAchGjR50+p+FpdQVbEGRTcXxgHC4uLapTo2ci8OUzcg7a+N9S9MSkEFNeLPn0uY309XWogYXxFobq2smbtnd2GaS/dhzKaNmEgICRhmJpzP1gHQsgcOjzUSKdpJbqz6wAyKKIoldwTibuaT8GctoxvAlr660Ljy8B1e1tFIdIhNME4XNS0CWwbNbuDtqLToutKtL1BHIsn16L09rMnxCrupXf5EoHA60giLAyLIkvDp/KOHHB0Or4QrvN4UCjo1V/q4wo9yRo/0P/PHzRChEgODXENKqT/GhIPGf6yR91jBsQI+4BEiYOZz6/hGAikFD4cSTWVuGbWDD8Lo4rGNM00mjkwl8bGR2WICoKQYRcDOjwLKP54PhQ47J9Lly7a5OQzezH9QpJMrlftlF/2Pc+ctUbzRBqdgSVCDKIpwdAyepSoARqGe3E4yOel+en3041D457neXR1Fmx1bd0RYqEQdMkJR/87orOiJAckAk2GOPxwJKtmakq2S+Wq9ffRfNvWfVQSJsaIN5UOmC+WtN6eLsnVRGkp4gGNAJJYyXnIN6GhBJXYwX/Z12riqIDEJM8RPTw7El5ir8w2pdeNdqgbP3MNYmJguBb8GxzV6UMpL0R9cKbETo1uR/F29fTahx98IIkaya1J6sgZbJ7sO9JfaA7YUsgOBckw1gc076jnebCHg7Ywa4cmlu8Ths9JFQGDgwPW19OpGEuxwH6MA2/uIYhChj0+RHDt2VgE82xBJVGoxEGiig9RuGlOubeJvDJohoolwZnhpuyuS+oo4qgbqpilAbBLf+lz1/YVE2m8ymKONRDOtbhHuSegd0GtCwUUBgro3LKO2ZNRK92vwRsBkTLMfmAQyPrdlYk368IbgmIi1U17T7InknXZC+vGh56sSZ4Vv8Na3ENmKwv9OScKfmwagNJfWl4S4ohCT0PKMGwutBf8/oRVDwqsXOP/NRW612/cVPEBApCzg+sHFSx5yLZWGxjsV+IOarjC5yjuSOZP7BQAD52Y8G6r2KRo4HwiJoNikvwNhaWkSmhWLdnc/LytrW95biCjQfZcnwpsDVyKO/rsSJOwfh48eGgXz591891EQuwAmpLsazXW9+vKUy5euqRzgNhEMQgjAeQajQkYTawHkKJ4Kz158MC6Ch32lS9/MfgiIFvWbBCY8i2tNjM7J4ZIs1B9fg5TSLIWMD5HaoL13D8wqPVEw6EcZDBpHsLAQHtaaxmAQCJpi4uLirHUKMPDQ+F+bereCMUoWQC0/HOSleJLvgVBxo4ci8L53r0H8lgYHBqUnvvAwKD2J4MHGsM8e2TyBgeGtD6J1+x99vji0ryMWvGCEVOip1c5HfttYmLC7t67p5yChufde3f1e5zP7BO07WOTIivvhJo0u0GSe0A2fT6a2JIpCew1GtAcXbdu3lZjEZN0GrTVatk21zfEcJhfmLOxiXE7enRCIJGPPrqudTAyNqz3xIcFZGhzS872imU7Ot5vX3nns5LwqjIYyzRZsVSz2/ef2OpWyXoHxy2ZhqHhkiAqvqW1XPNh9d6era4sK9ZqiJrwQeLbb3/Ounv77Z//8z/UuuN8IsaApo9eVwoUypMC0leDBR+OI4NC7IzFLftWqG+hjgNDlOGBpCs3FQdhfYCAJc6zZ3kNDb5CDOabq8trNjQwZOSBK6tcd1Vxrr3dQQA0SzlX/JyBlYtsGfmANzlZy86E88YMe6g5nwvgAi+MkXckvrgXBeyprBq7fK6+nl6hcTVML+1JNo8En9grBqhQhiVrac07K47BOggVgYYyYozJa0tMS0yl9yXb1ah7LsV7sF1gTSeSGWvv6LQPPvzINneQkalZb2e3AFU0ZJHEOHnihAYBfJ4SQy/QoaDx5+eUz3LftzXMALGb0WCgTpMrnFQysQwN7uZci+49Z130ASIWd3V2yVeF+PLs8WPtW3KC6r5LssK85roZ1vH+MI04myTPtbtnx48f1393S0XtCaRPiCHEJAFS8HtK7AuR/Cu/+CUbGeyS9NPa4qLNLyxYZ1eftXX02d0Hz2xlbcvmF5bszJlzzihHQjI0XsgrW9va7dbd+9Y70GeNZNImn7+wV169bB+996G1teTs+NGj1t7eateuX1OD+9GDJ/bOO1+wYnHbHjx8oMHOdrFk9x48EnKZYWZrU5P1FtotUavYzsaGvfPFi7a+tGwz04vW3tVtm1Wzxe1dS+faNeDmeROvM1l09x0FTNwE+AWbgdwxJeNffI+4Tz7QY70T57q6erSOifPkb9pTyYT8FtgLQ4ODOuPYx5LXYtBEo0z+Zj7M4/wnHo8OjWid02RUM08+hDlb3ViRRr1LzroUGrlEbA79+LDCh2SwePFAqMu36a3XLmoYsjA9ZYN9PfbG1Td17nz/e39hAxMj9nRmyVLZtPZ2X++AzqaRsVH74IMPXUbZyAFbNeBiaIKxO34dMN3Yv/19/dLgR5KIGCEGJwE0IKrFqsykxYLga2ZmVlK/7OLjx45pyAdoyGVsXUo1fkY313VWrVjg9brAXKCXOTPYazSbMdMmt3TgoYN5BOhhSIbk5v6+jY4Oa1DhoImqwBECLIZn4Swzl6tBVo4ckNd0WVtnm0eQndheAaokqaIAXFMDMQyRNICXnJuz9GHrRaAfH77Q2qI8HkbFuTOn7MatO3ouAI8uXrhoDx890ufBTFua9SDxOzvFqOCeXLl80cqlTZufmbJf+aWf0xm1ODtpnYUO7e3NjW0bGhxQLFlaXNBaO3LyhEzIYSSduXjRbnz4obU2N0u6C2AX8pYjE0ettb1bBvdtbZ1WLJXt2fNpW17ftpb2gmSzyB3I9axRtc6OvDU3peWXcebUCRsfG7N0W7uVdvbsg49vGsIEG1sMK2ASZQ7OJ9Y1z4UGOHVDZH8rHknuB0WKjDMuZGruDOToocS+YU8AxCCm0Qvi97jvPHNeEwAQwAPuAcChbqTWqHtgtsGA0/7nulJay0yyJeGKOXGoU4p7Ze1XGDC8p+SJqK0CapHPIPPkPOeEe05SDzHcpA9Ew7YN+W3yX/Y10mJpQJFEdcyRm5XjKNbX3T+IIT45BFLkgPD4YgATB+vEfmI0a11DA9ggQswjo+zfkxxW2AcwMhgoUH8eeJOaCWBFvk+M497x1cZZCZNI8oXugUHPxr0IXOaZxa8meqhZuB71C5SXUH86IOOwuIV6APLQQX3CGWYRGOH+qQyPfZ9p0HiodxGlyQHa+leUXgKQBTDUaykfcoSfOPTm3rOK7AMHB7oZtzNP1SeK4LrDbKlQ2+tRBwCrvB0D28P9PYhNDZ0J7hXqbDLOBdQJWIvkiNHXlX4P54HUIg5qex8WsTbIAQBHco1ScomMkABWjDE/1tDU6cRP5XEM3UKfxeWuHaDA61AD0Fvh2pX+RlBykI9ygLYzRyIAm/sThxERpnuIaHHQl1APJPJWYmDUcMNBieypTwcVYWF++p9Pzh04191n86Dygv49mw/0Gw0PkiUSQZoEjmZPCd1BU5zGMM0pAiXIPUcwO8KdABBpmhglsQGR9yCBJFhD6XN6tjeFlCwJeOuJo8AhoYlOY83pnAwGShoOULxFtBPXpLonaPrHg4NATSFI8OJ3hMAgaIfiUSE4BNho7M310Dig6OBw5GcVPKAO513SBkOmp0+nraurXQ1eN7d23UZvmiqF0vVwz6LGbUR36T3C5+QnNR0m8MjEtaJhD/IfHAMU0RxcJAIckPKiqO1bGwOLICPFtXZ2dQm9SMFOUamJrJI+/8xisuRzQjiQ4PPvUfqGGy2pEKHPfF3T9Ig6eW5+FZDakttx3WCK0pf6gS+RTGjtJhMN6+3utK6ugs3OTKlpQRGGLmquuc02NjD9AmGIDiIf3guCeMjx3zj8IFmKjcV40MWEVhqXeyU1P2m6sE5I3mVo2turZIfHwRqgWcN9J9FnraIB6ZRll5Th4PMmoh/+JCE8TJkqh2RZiXLwgYgRQM3Qg4k/NFRPXriZburuzV9niXgCrUFMaFbFQzl+/nj6HyJheMOVwt1VeNxAKZXypiO698G7g8/HZ9KYIwwplFg06kII8XhhAlH4sE5pfsXnq+tLeENfa5J/3y6qkcGeV3GRSgvZq/scDmPtq/2GmmqYaEYtbu7rKKZ6mxu2tb0ZENEuYUFMkDxcLucan5E6GWQyYGRJfieYbSlZVQLkSZBQ6lvbgZHitH4leYE54SgfNFpb9JwdvR4a8GEoxnr3wqpuhY4229recXmv6EMSqKuRqUBcQEZDSGgQoGJAUUB4bFKCEBATjsIOJtk8i3DdPmhwlpmSblDD6G23gjJ1JCwxi+RKGqxBi5y1xDAXhKSa3cF0nn1NzFXDUoOEID2kotH1g13SKUpfuQ8L1yu5ETNbWl6WpB/FYmzuu2RZaGpHH50g0eef1dkFDAd8IOFrIhqzR/quBpHVinV00MzbsWqlZGdOn9I9oyEIChZmhrxtkN8Ksd6ZCM2OVA3GyySjNO5A2DD4iQmvzgaSbtDTQSqEs8wNx3y/yach0IzdS8WL5qas64mLxRMYOTSmXLLLDVn3E/ui8hN7iQsUY3xpeKDXSjkVHNNrxWtHrcm0NiB7/blW1OTnzxTBNIGFxmnDP4VBi6MaNczjDFV85Nn6M+OL4l4xpVIS6jgijfwvLq/G/WZvsWd3trecKQgiGkYGEirhvtAqn3w+JSSsFOdoVAY9Vpm3gZKUvwxndFXsKNY/xePAQJ834RkyYjyLoSDyWDR2hXRzfWSGBrpn0OMx3FSjluYgyPq0GnpLyyu2uLRseyUYmQ58cGM4Z11Byee/rDkNRXd2ZDS8trxq0zOzdubkMb0mz4cGNrkJEkfIyPFs5mZn7dz583q9qO9KXsN+5Qt2FI0dDWF5fsWiteRz9vbbV+39997XoKaeSFu6qVnIW0eX1dUIV1GOlAZ7TG3YhvWAkuzp1foENZtj+AirEeo/hVqCBpgjyDgDaArDkOC5M+hh0VNoHzt2VIjg27duaeiL1MaJE8ddUi3p5snkGxHtzh6IzJmhgQE1GRnKcFavr60rPtMMm53ls8PIS2oNHpUut9nz55PW19utODM7syCPD4ZknIPcH4alpUpJElIU3VFrnL2KRjwMF5psxDJkS5BF4PW1VyQP2mF7sDaQ4cBUEUmCOv+Ws7nZefkd8P2JiWFDng1961cuX5a2P/Hl8uVLjjCs79v9+3ftydMX1tLiOsp4SmxvwRhIWGtzk506dsSOjo3AlfdyqosuAAAgAElEQVQc09L28MmkvZhftXxHryUzzRpUeK7irE3WPvuR58mgnMEv2w6jdcxLjx0/ZseOg35+3z7+GKkWhgfkUe5vRS4YQTK8ZjSLjvILNPZj3qKYZQ0N8qLWNywiGXMGTW/Oh63itgY8PkjGq8W95LQPg1RRqVhRs6XeABmLjwIx11HHeKvonCZO4bkDMpV8nPins8LvD69dKLRrvx49esTe+dI79u1vfesgB1tZXwtm92k1ejwWgir1hgtSY65jXtbZRJODmAKyNpnwwXGlUtIeo3kMnoD9zrpi+EX8ZThR3yfOZiybTipPlXRD1tcOTfbdUsWHhrV9e/fP39eAuaOlVecEAxPyVgyANbDc2lKMWVpdlhkp9w6UOjJRJWIqnCXkPTizaUwDGCIP4foSdTWIaTjwjHmWvAd1DRJSkDzJpdtbWuzRwwdaK8pVGMqQf4V4LclM2HXIxUlWlc9Z1TAFiSziPmhc4h+/B7hB8qOlonV1tFijums//9XPW2tT0rJJ7veehrmjY8cs39JlH318x2ZmlmxqftW+8PmrGhjduX3fxsdGbHV9y8ZHx2x4ZNi+++5fWP9gv4YCz6cm7cK583br4+tiN544fkznJ4bP4xNDuj80UwGmwFRSbZVpso+u3bCW1jYr7VWsCwZdJm1tuawtL87bF98+Z9WdolD/m7t1W0Z+K5+ztq4B29ksGTJJ3IdSbU8splo5SC1y3yWN6Axgx+C6xIXXRs78Ydiys7Pr/n8AWIIkJQN59sGxo8cU7/g9DUCUTzHscuAKuRuSVeQ4x44e188trSyH4VHK2jrabKe4ZXPzC8EjzpnbBzn+wZ8CmjzkUCTJrB1w/PiHfPbq61bd29OwBymt4aFeGxsbFYu7WK3as/kF29nFQ2hMAzBi5NzsnLw3WBuwqojd5Oqzc7O2vLKm5pPq4v19mezib0KsJu5S09Fklnl7aNYTb0ZGRnQnMdMmXyHHZDh2+9ZtZ8kGSeUInjpAzIeaRIoCQUqUYfe9u3cPmMAjo0OqpQC2OQjYm5Ji8Squ7YvRR3OcZ47iQZRW5f1i3RnBNjwLwJBcl2SMiRVBcsaZGJ7nOPLbQYVep/maEvOcYAMLS/8MCxupFf9n5NByeKalk9bbXZCR+bVrN9SPoEZEMvHunTuS0gK4IHa0JcRWvHnzjnW0t9grr1y01ZV5m5+etL/57/01a8omrVF17zmMzTm/kYHraG+zxdkZSVH1DAy690RHh527/Ird+OADsdSOnzhhk48f6/xobeuyfHun3Xvgf8ftpIzkkwbpzbZbqqppvry8aNXSrmVSdTt+ZMQW5qZtqL9X+7ZvcMi6Bobs+vXbtrS25b4rNQfOcUOI09xX1UQywXaWMnmbpChTgDcAs6zoLOCMZRCwtLSse0+uStwDAMle7Ors1qBBXkv5nM4sci7kKeU/yrlUq2lgwKC1iZxQsrBVr7XJJ1k3yvWRRGL4iDcpgE8HUOLHFnsjFTFVXZaSNcZQnbzIpYmQf21SrRc/F9fk8oum62BIkWt2ViJyopxd5ESAa/G0idLcqo3XVv2sNZOcL/dCMqtBxYIzAikz1bjURwyZ5VXjQCnVitTbgUHvYBtqZWfFuq+o91aILwJ7yVvOB3BSrQiDB11EOEe8NvfYE+WXDsChoWaiHnMmfRjmUY/Qywh9DdaKswocJBeN6GNz3GVXfSJEzFcPJrAK1CcL0tdiYgSVAN+XoScR+jfOTIhgTJdgF5guSFurLxF/J1Qw3ut4yRaIlY2G9oCWQ42t+w+IUcwcB6VSf8bhCzkxoJ+eXoztvTfE68Y62wdbrrLgQ128RHYDe85lLFmHkU0U+1A6k2B4UGOEM4ffVSxjsFV2ryyGZmKnhZyXvzOgIx7E5xXulv4T5en9uXqPQ8C+g8HPSxbJwT07PKg4OJcId95zVO8mPfBGfC6HfuTTP356B/7q3oHThS4hktRgDWhTUFGgM2n4cpBFOQ42Ac0QgjKTS74I2hMT444+h/aVwJBo19kNyNQEtB1NEyGTxLpgclwOmm2keS59QwChYSdEcaBa8R6uU+jBE5SUptfBCEi0qIBUjX4KPvF21K2aghRCvJ6ogoEiG2V3iLtIWoTmIv/Ka+o1hJpDQzFl9aRrRKNpDKrMGQAuQcV1RQ1ikmuMqyIjgmk8QQ06GoetkspA4SfQ0t7g3vvAxeUQttXYDSgRNYr2pYvLkID3jLrrBCdOZNcRpHHoiQfPkf9TYDmSYk+NDSWmgVIW5WEUIEXBd407niOJCkZvUIMd/eINd56/WCTBe4NkOX5OUQcVcCnooNVnraMDuYmUjG9J/JaWVpzanckTVkVrpelIwabmbqDzehB3+ps3JIO0TNBxjMMCaf6D+GvKHVx/pNuxfmlCgUqm2UKyBmKCKTvyALBjIhI3eoJw/bqOQGOWXqfuTxiWBYmkcJwENkU4EkJj2wd0jlSKe+LgNA9hIrJFVNgHWi0H8GHUlubmh5AK3KMwLzowr4vUQGeRuF9FRBOQPPI9H6J5sQ39XUOavT0vDEXL92RCe4ymQmhcdLR1qDiSCS7a5Uk3eedeQY/XGhO93hk3an4EPxjWjBr6tZqQsCSWaEfyuWEVqEkimaNUGHg6ZdIPfhoUm1pnh2moavaHA59kkoLaD3SYLH7dkmcQOsSbIxQOrFFPGIPWaYhnfGZp6LJnkP5SE5ommieerAP2v6NTPIlB+kF0y7obWJHsS0kooE64XyS33F8SOiVLJCoZ1/+M/hhKvGS8hkRQLjRwkG1gAOAyTmIvhefPfZIEWTB/579CzkMRFmPNkyMZumvg60wa7k+MByw9NeT5vlCyzUrq+Blen5hN4543j3qr0fRVA9es69fyuz4UcnO9SP1XYy/EVt7HtdFdysiZGlVra0Uj+Kytr62p4MZomfvghUXK7yveRvh5EK9oJMl02Ye+KrBo0gtx554iij8h9ZXGquSuPBkXXZgGNR4V0GMly+TxP8qG0LyGIcda4FmBbHJpNF9bbqrkQ+vIesIoz9cacl7eLJVWO/swkdAwj/ilQZIQSxSfaVGC4/AkGoRzR0HBgkz358jnBYFNzHazSRo0zqpwT5ZGw++10OBCGLqMUTTTxeOABn8cagkdBgq/uVkxUbI/mawkN+bn0br20iCiFVWoqAjIqxjv7xvQwFLoLujqxW3dd66FtYisEw1dBgVqJDUaAi8QD2BKsLaIQbHIo2hDb35rZ1voR2kKy0QcZLJTnmkyCTkleQEanVW9OUzFVy5ftJkX02rMjQ4PK7YTDzCjZe3Ozi1YobNdgyb3y/GhHbkI8Qy/CvYBe1lowCQyUe1WwkclmRSjYmR40O7fu6+znzEEkgqMKJDvKZd2JSVBAc65z9may6RtdGjQ2lvaDkAfzTAw90q2WdyzHWIF5z4objVxq9pLAjAIhFG2zU2Q1/hhbAu5ymN58uSxPF0o4pGT4XsbG+sy8uX5zM7OquGFJ8f0NP4TXdbX0223bt8UyzM2z5EQisNFnj/PGuNWGKLsCs4G9xNpsvbWVj//Q0FIY6qto11nJxIKfGbWrA+lGS5MSIKKZw8QhWfDdUhKLkio8expDnUUnBXqA7+ElfacgfTsyRMBPNrbmjU43tvZsatvvGEPHz4QchpjzFdeuaLmM8UiA5wC/h3SXGd17+uaiG6dbXl79fJFod5dWjNr0/NL9vDZjNUSWUtmW1zKK7Ai2fNCU8vLgSFlxQeiSF21tUn2kJjzmc9+Ts3DH7z7rhok7LtE0velCt8UOVtNqHMQfpzB/IwkIkKlyfW6Bn7Z15yQqZ5fSSZPABPPUzljGTAp5xJ4xRuCQgSqYQtaMpy9GMmm3biU20EOT1MZBg65sBpV8hjKKkeX+WIA/PAeS4uLGgoQt0DWv//+h3b58kUxxmj2PH/+XJ4moyNj2k/k/5xzsKneePN1e/7sqYajayur2n8x3gEgyTYlLc+gMfi18THxpuju7baRkVGXXeOMS4O83bMGAxX8pYKhMX5vaG6DMN4TmjRl27vuWVer1LSnMTjHWJlYf+HiBcsyAMRHL5XUfuf/rKO1jQ2Xg2OlwDIk95F/VFKN8irDA0lUMLwpKF/RcCb4i+hcQway0CE/k+fPnmlQoUY8QwoBm/z48drEWd4OKnVmwamTp7R3N7c35KFA6gdTy/NOmHhl62jJWXW3aL/w81+wjpasZZPkYru2vLxiRyZOmmVb7NpHt6xUqauhWegqKJ7xnHjmPDcMfnnNP/veuzY0Oix0Ns/m3NlTdv3aLevrLtj46KgYFVwH+zMLswE502pVXgQwAGBA3773wBuMlrJBmCJ7O9YAPJWs2euXj1oSg+C1Lcu1ddrt51O2h4lzS8Gacx22vQkTrm7JprQk5nTfg/FqtikvkAg3SEM9ckrJCTlilmeMDCEgDQauYtio4Z1RPkbsunr1qn3wwftai6wxYoUkMIKkIINHMTSKu97Eb7gfFF9qyudzWrszs7M6S8g/xBSN+kOB4RwBA8ofYibBHlSK0LDPf+ZNKxWLNj05qbOMZ4y81fz8vA1NTNj712/azl7VThyfEKIfhvzo2Kj+HXlcWBIg1ll3AEgwUuZL5yyxqNCp63/+HEbFxsF+8mZcYKHu16W9T+xA1pNGHp/lxIkTdvfefQcSBlAaOXD0kfEhgEuySE4klRLjgDxNDLIgzUg+v7m5IekppBBDx033mngEQ4J4Ql2H5xP+CrFpFq9R9VEYWiD5x5nNWUJfIQK2qHUOcqrQEBVzODD31SQNzdGD4Jp0GUNv8CYUG1xq2p/PQG+XnTp53G7cvC3AFoNSZCTxcEKmdGxsRDkD64X4+OjxEw1OX3v1sgYVzx4/s//oP/jr8o5pzmestbtgNc73jU3P91NJm5mc1D3oHRgUg4WT6dSFS/bg5k01zyeOHbNHt27L42lk/LjtN1L24NFTyze32u5e2ZZXN62eyEgaqlRxEM3y8pLlcxlrzaWsu7NVssq0w3nPje0dyb9NzczbZrFkjWTa1mHAphlIu6efzg5JZHlznPXlzVVnuvB3wAX0KjiLqf+JM9RtDFQBrHmfA3ki9pbn/pwj7EOvNX1PU2tXyxXrQM4IP5mQy8V8FIS/aqtgciwwHHVXOi0ZXHLBfN7NsukVadhQqaqeECsK8CkyUCG+Zhia75OT7mqdo54gf0KY48GTg2mi2j0g8CXr6r6MDCxgdUf2jsBjFFApYiFy1V7bcjZHtjX1Fn/3OtbrEgc2uneFmtrUGeENObsk4yjvJcylHUypszt4UwnYGPocznCirfOSmSAmo+RXfYAbJgEHzCjlDqHWAzZJLhLVQuIeibV0jGHehA+MhwP/VpgS/voCUwZQprM4nXVO/h/lpSWYGGq+cGGHfB1eypvH/ekvHeqvIIEef8+Hji8HwV6R+KBC7xu83vissb6TskKNPe79H/6P9xX5hPcSHagaXCED+MnrMvflcICqeh8KUkE5I3ijKD5Gz1GkWZubvXYI/caDexsAh/4iHtt4VzGW1HujHvXekoNIfRjivU2Pjj6oiCV/jJhxUOGfQVf4lw0q4jMDlMc58OmgInTaPv3PJ+YOnCp0uVa/pFgc8cxGJzBQjBAE2JgcBBwCMtOu14QkiIUNyFiSf4pcGnX8njdU3AiZYEOSSIEvSqbvuGDQ640KSdAEky0m364NSrD0Tcs1UNSxyaM2G9+n8OKg5L2guXJN7m3hgVboNdHEPJFSM7cJbwY/ZKTJ2Aj0NGEaXC8bBBTIbhIdNA6rAUVNUYpu5+qKS8pwsMukqYwppntB0FijQQ6iMaIf+czSBZW2fJB7IrBwCMqkCpymNw0x1Ovq7tRnU0GzsSl6d3FnW4gxpvwUvyTSHKYET1CXHGQc/J3dXWIYcHgKUbm+poDIz5JE8Gw02Q7MCoZCL1ktmAG3OUMGqqbQj84KUHMNymPNadTQgrm3PG+eUwcoMdFMa0KlggAb6OderQi1nUxnbXl5XTTvUgkvBJIpN2aNbArpZR6iXMdJsxBrQcYmTp65ZjdcLIuOz896A6BDzW5p2de4J1tCUJAI03QBfURhEguf2KxlzQh9zYnhKg4HeUH0cpC8UENHaEAJOCSP5+5Nb1DInty4kbMjFuNXRBY4ytAbGUI7MuhJBMpE2B6HgwxIoTggiXJIOhDl1eHPk88f5axogvAMuSY0bzkghSAo7bpcCXRfXaczmqQ5Kf1X1zqmCOQ11HClEYMkVNobUTQvKS4pHg8+V2g40rh1Kizaqq67XejsED3/xYtJb77km93QLAdl0pQUR3QC94PGLPcmoid47uyz2OhgHdOkJ9GIhqMuKxUk4GBdMHirI2+CUW3bgYGo+904a8gTBG/4klDQlBTlOTbHy67fStOEXxKzh4Qd5LeYWk5PjgaAzgbzoiDqwCOpFdHqXoB7MhGHbP8Xe+/5HGeWnXmeBBJIg0TCexAECIKe5VpVXaZVqnaSZnZCGmlC82FGERu7od3983Y+bcTIt6q7WZ4segOABAjvbXqz8XvOvQlwtnv2sxQFRYssEMh88773Pfec5zznebjvUYJKewfZrVJJI9P+FfZ9DaA1pWKAIkN7NhhtsW9gOwNG8uVeM/guBLZv2NcUIA7EufY5PkOsmydkaKx6g421kayQtG09RsnWsgnAmBFjkWeHNfBpDh875XOqCMZQuL9PjUkkr9x8zmxwoN8uTU8JXARMIOkVkNXRofMBEJIv4gvPKPuL5gn3GwBBZrTBDJp1hm0WfRm4p+xT1kcN1RJSJd7k1Gg7SS1+EmoAe8MFgB1wIBbpnEM8F2rqtu6l65L68+l7Rc2E0NBT3MbETJrTHdaJtjggtsy//XlmPTkjVMzRSJakla8vzy7nBmvKcyl5sHRK7wXwRnNB4+cp/CUKLrPTrFqp4mwwEm3WCWBKo+lhejDLXgkJN6BqpdbQNcBSRrYNcGBzY8vWN7fDaLZr/vrnaqgYnJqesr7eXhWLFPaAdc5qqin5BkDlfOI6YKN1dXWrOMTHgD18/eo1u/PFHZlMnxZgNznZUT4VwSyO+0xxyJ4kU/fY4cAe1682oM6DuggO3LeZ6Rk73NvXGPbY6IgAqvX1Dbt6/ar2ydLSqs1duaR7BiDE9QBmalIHWZi2NjEFWVcKceIo+5iJkPLpqQ329dhAf69rSdfq9mp13TJdeemLz1y6ZKzty4UFazaq2sNMykyODVtvV1agFTrJPD/lWt0OCiXr6u23LYym0WFXvPWRe75g0gP8ci2A3DCZMWiF5UgjlM9OXoOxqYwUx8b0OWITHoNZDMJ5PeIq/kVMsdHs8PjdLpNiJhqJmbBXZepYLutM5Dwkn5ufX7CpqYsiMogRpjMFSbGi9iDG0MSta9ev2bfffmv9vZhwIx10xn4kpgMuSFYnjNLzLEqKo73NNjY3tO40FQCdJZFWd0YsOQIa+d25Trty9bK9frlkf/LLn9sXd+5Itmx7Z0drf/HiBTV379y5Y6+WdiyboRGBLADM6aZVSzXLpNrtkw/ftcszMwK7U5mcraxt2zf3H9veUdEsmRGoHBvSEVgQmCDNbJ5xZ9ujC39ydKQJvs8++yNNvv7DP/6jGlZuJkvzlHhLI9SlMfXbGEHKDNWLc9aS++MNHmQw3LyZ65ZOdyJhw8ODkh+Tz0cGhq03sol77F9ikwzXjT2XD95xnAtMTiDpgEQHJBXy+KTt7x9bvYZUAibpTXnKMNXMRBOgFPGJBp9LCLaJ0Q0IwITtr3/za5ucmLT33//Atna2FAMhGzx6+Mg++PGP1RDguQFEY9KH6dkX888FBqyvbdvBASb0bWIUXrs+JxCQs5iYwd6VdZFin8tfcX5pv9crkicF0CeHIB9Q3Eml7fDoVHELGSDGSzWtlUpZsVCymemLaoDT8AY8+8M/+tQ2t7f0uuSbxEhiElKQTDAIXKrUJasiVjw3ggZ/BxOfSM+ZTJyJIeS5krxiohl/vvV1NfMAJr+/ey8QuJvWQE4zMGaJY0z/cHZxViPDxbnCWYH8Lb4LTLKfFE+V51D78BzPv5i3nlzWctkOO9o7tL/8i5/Z+EifdSYatrr8yl69emmX525YT9+IPXj43Cp1YmbKmkxzVMquc16pa/Kbe8T0yDff3bWJqQu2f3hk23sHdv3KnD24d1+sbBj8NP+5x/hRIOdIvKFmoPH5zrtv2fLamq2ub1oJqjZrlUhYf67LGpAGykX78O0LNtrTay8Xlmzi0iV7srJuC+s71pkfsKNDzveMywBZ3SqNqnIbgWRtyPUN2v4h04XOlKW+IpaxVrQDOM+uXL2qM3Vrc8t9otRga5NEFufBxx9/bK9evlQdODQwIKIAMnmcnz6hirQnDYiq7e3v6/nM5twjRdNQCWqeHp0BTCsIxAugGue0591vgmhONvKzvyNI3v7kow9sc23dDvZ2dX3IlF2+PGO/+tVv7L0P3rN7j5+JecukMU0I1gRWv/LaZsK2d7YVC4nLNJzYEzrzuzw3oMahUby8tOyyrQFo41ppUCrPrNdt7vJlPSc0KgTidaYUOx8+eNiS1NVErZpBAHfVIF/qUqN88awwGcGep5HCNWK6jpwbuZU3M5Ah9bqDWM76ZbP4ZFEDeu6MpBnYAfe0pakOoUlSrC6B4t5dLnVMM9WnFn3N+VwCToPJs6bJxXoOkxQtj7mqWRvsdW8cy8eCszidsRzxoz0hE+pL0xft4aOHtrW9q0bFjeuYaz/SuTsxMeE5Qa5bcRsSANf07rtv2f7Ohq0sLdrf/M1/tdVX89aolWx0fNhSSDFCsGrgIbOvCSMmsXrk5bRouXzeLl29Zve++loTCDMzM7ayuMiwn01enJUvxd37j6w736eJy4ePn9vxaVlm2jQhaXqmOnguqnbt8oQmOZCdHOwHB2B/VKxQqdrK2q6VifudaTs6LYAkuApF8ArD85MGIXuGXJF8jXyY+MQEKo0y9oPn990+vQd+wISBJpNdPSLZ5r54AozD2Ub+EO8TfhLImnJ9TEUq32OP4SPXSe7o0xVMVnJSEudFrmtvt53dY51jNGViLc1BQS4tvwIRMKmXIMO4KTfnAMoRTuLB18GJX+SOqsNFeHV5NAgIki+STylYgatOTF6YkFcJUzUQawrVsmIiUySey1DnMOFOHepxQDlNqM+cLR+xgjM56Dj9yvv71JgD027+7tJQ/BrxSCA1eUIwgg8v7SoMQcovEmi5dgfQfbIoSkI70O+SQnzJV4RkM2A9apaHRgE/4xOeMbJJqkGNtTjZzvmlfAZPtuBr5f50odkpoobHndDjDH8PChJvNBJ9ut2vMaxRawojogj8eT7OBgWL8OLRt0syZfgKEReRNW80VKdwHTTXiTPce+qCOEnvtZuTuUS8k0eLxyw1isKXE3idHK0JCdYoTDk4waSqmjkSRoRL0fjCZwxsTYQLf93WFEmoQyM5zqfBwu45N0kSGxVn0yW+HlGJytf5nPRTfBGmhwLGSa7+Q6Pi/H764e//JlaARkU0uuYDqcPe06MDiwQl6l5HoyuKBg6KyMbl4YHpJ/BMiUHaGX8YCwY2ZGe6U4kAhQoHmsxIKYaV3MBCcsayZC5kluzBSgCSOtSeUPHf8QDzzqqDqmIYZzwhIxjIXDAEC7E0gjktf8pUkFFDz388wPImoUPPN2Ciwa6mGCQxfL3yWoxPimwHc/y6+TeSNpkmAY6qqHQjYV2fpK0AdRyI4JqQ1ZI8T/Ap8EDqprkcExSOBSQSOjsEXrEuy8tL1imQuE9A0/DIqIoQxjNJyjXOD7BVIkHPSncbIF7jlmEN9RGDJwABWCEwMFRJGluHqJJfZ7dToJFYM9aJ/u/R8ZHAezc+chMtHRjSAG3XtVHA9ff12MHejrSmKSRJXmHWcJ1okKPl29YBc7TkiTECr14ZBOPzqM/vzS7d/1A4aB8AFCODEgy8ojEYhxAvJB+RbFaMXPY2a8m9gzEFI4niAvkKkl/AHDVAdM98D1OU8oaxORLlkeJIo9ZS525oVrRIDm+O7fFzJDpqmIUDyZOaCL55d13MMYEWIXlvHehnIYbEX8yYwO4//3zEUUbALe63/CUAzaSNjT8LzGiX+5KkUqPhmp4As2WXdGMNuRDWkJ8HUAOMdCDKOQlozbLHKYb5WXSBHUSlmenFpxvqOouHIkEj3sVTMZeGhge1l9UYbG8TiEgR4yBrVZ4GgwODAnjY375Hz5hTvBZ7WgC15Cc8ieC9SR6i5BxFLsU/gBzX71qSFV2zj8jGcXVn6wNE+URI8JqgUSNTeKWQ3tQkCZFXhU8xyMBZ64MnAGOfHVobgFKtH81WjGR5VjB9J1Z5zulNhpDksVcB9cXSiVNLsDAY5Zd/SrjnAUTms7Mmblqb9skAdy6VLA7f41rkYaGxaE+sxPhN0qgiVrUL2OB5FRMosDriBJDLAPpUlpiuMpT3ZBsNdcWY/X2tLfeMWjKunTeczRtIMl7Fj6jTdnYP7Ufv3RQIhbfJH//iFzIZ1bg/64rJcxqWExqzjOPSzHEjbRUoMojz+EARwWd034JTPb/eqPXr5qyRebL0pl0GjevRiHjZG1LsAxJdN/z18wXNakB0aafDHmcaCzmS0OCJGsvilUrywM8eaaJL/gC16obABWmqBkkm2GRMcEWJKuIvsUMTJ6H5xTmliSQxRj3+8fPS4A2JNbGYs6thNetIeYMJYAJgkYbOgwcPrVz2KbKJMfcnqFRIzGlMYZDqBR1r0dvbb69eLdmrpdeuVx0YkWocaIqwaRPjoypUfVwaZli7miouB+AG9cQLAMZcd48NDg6H2Ov7n2BKM2x1Za3VPJMOeRL5Iomy+hSQ6mCfNuEzt0wEaYYrpjkhgc+PjMP0xWl5XgEq3bh2RcaekC0mJsfFWEPaCdCNveJ6ymXlI+5DUtEkwcbGtg0N9et1VJA06tbJmiPZ7zMAACAASURBVFcrNjU5bteuXrH7398Ty/HlyraNjY/Y7uGJDY+MCITe3tyQ/AvyKRhqvn1jzrbXVuzy9EUrF09cC5rnpq3DTqpN29w/tEoDVhZAM01hZ1iJHJJMaiJBn1UM7BjzAKRzzrYPUmzLS0uaVlEcMLPl1ys2Mjyk517To3xGCCFBw5gYzDOmkXBkCnTfkMFDJsXJBjzAS0tLNjkxIYkpcpBrV+dsZXVdzy/SitKDlwxPTuxL4pPLDpYE6LIf2M8AbzQdeDYBCIklnKkHRye2+GrZJieRNhm0Eya4AhuSySmajHu721apFOQFhNn7L376mf3DP/yjS4+ih39asLffectmLk0LaMY3g3XTRJikHesy1C6e1G3qwqB99ulPtEdTqay9Wlm3X9/51lY3jqw91WFlWNM0+hQfOIPdsyHw1gTCAErMzszY0dGBmigffvSR4srf/d3fB18bXhutam+kc46Q46BFznOBL8NJ4dTlp9Q0L8qLhokn7iexVNfHFFmtqukgq1cllUe8oHHCfSZvU+F9cqKYBBDGehMrAYZq9bJyqFqdCYrYVOWZNVtdWRdxQ0QR+W652aOzYpGh65cEG/GD5kuhUFIz5osvvtVz8c7bN2328iXt563NbRFkICkNDw57I0z9mbrNzs7Y5taGbaxv2MH+sW1v7cmXCK+v/+U//DuZAH/9zVf2ennF167pzwDPF2tI3CS2jI+N2OBAn21trCu28hlp5o2OjWuaAlIDZ7PMUZlYlE9Qj8AxfDIWF15ZOpvWVMWt27ft2fNnAoAIR5zZnFeA90w4qzmB8SwkBM4tjlEa953k92V9j2eERqdPnjIBVFLj9sGD+2pMCRRTPkH3kaYVbE00332yTAa21ArdOd0z1UVMIkhWqml7h0fW25MP9U5Cz8/J0b4lGvg/HNpf/MdfWF8+Y/lsyl4tztvy0iu7cuWG5XuH7f7DF7b0ek3rgjRZsVK2pVevtV9OTwp2YfKCTOC/f/DAxqcu2NHpqZjCM1PT9ujBAxseHLSZqSmx3+8/vG8Xp4mZTJT1aSJvY3Ndk9DHxaItLr22BOdxe7vlyOuoqzCSrpTtR3NDdmtu1jbXNi3bN2DbpbL9P5/ft75RfPISVsUcmDXJpqwOqUf1RUogNnuOM4Eaif0IGY6GKhMd0aCXpgJgHLGbRh3nHaCvCCzJduVgSEvSYCEGEqtYb+IcPouScAwymtxzfFpYeydpMCnPZBzeBO22urriedxp0dnCMWmLI1GelfrvJxNWrxJzSOAb9smHH9jrpWU7PjpsEf7GJyftm2/v2js/esdeLC6oYQZATrzxidQOsYAnxidFAnKlgoQ/Z1vbauLx7JOvY8INA5wmhiaFA/Aogowm6n1qGIUD6nHyc2/cddrY6JitM5UvH64zY19yDdaW+BWJT5HdTV4+PDyk61FtJF89B5Ed8PTcLOYrxLwOGXRD3DgVmcslTV1a0ycjXVbT82r03PHMcga6wD3WtdMJPapflRdQnznI7o0K9wv0STqzTuKHSFt1S2VSyr+YbuN3S8Wy5dIpxcXR4QFJPz169Ng2NrdF4Lp27Zp9//33it2XZmdte3vXLkyO63xEdhAs5J13btvO9rptrr2y//Wv/8r2ttasUj6xgcF+7VmmkzO5HBvJTo4OJHmXzvfY0wePlC9MTF7Qe3Cm3bx50148fmrdubwNDY9bsrPLns2/tCZS1bWm3X/wWJ5KdcyJmzQ+kRmq04Ox69dmrCeXsoPdHevsYGI8L6C+UKnZ0ut1K1bq1g3x9KRgJxCAQv4vcg0kEE0tHGgaM+a/TMeT92sSAblZEZZ8qphcIoK4TLJ63eIgrerQIHkEgQr8geaGZE/bEzLTZiqSc5RpXBFozoHa5Dncb4B5l/Fpt529E8tmO0RI4b01XS4TYvdlIt9wL7oOxXRvMpLzOEueWkXy2FXOQeSLm2qK0yDhjJFEreR92hWn+Z68506Lhj8G64TkX4PPJqkx33M0JVym0pvjahDws5LVBaz3XE7fD00IB7sDHhDCiOfZgMousRzxk6huEfezjLaDAbTwjiCvRjzjeY5TDDL8VtPW/Z60XEG+SAohbV4vi92PRG1LXttrSp+88HMt4lGqp8PEh3CXMJnPNTI56ERejxWyuXhjEsDrW+0NfXavq2Jz4ryyRATjIz4VicmOeITxU5H0Qg3sYIDeF7I0v89+lt9ZwL2oU1Aj4Rzg++Shlarvo+jjyeegLkbiU8SpQELU2oUzXjhDkKYX2TrINmpaAnJsmNDWa6Uc79PUHuoOQe49IjdqFEly3j1DJC8dGk1xP8TJFv+dN/1GvK90JpcVV+f8d2LzSaRrfvqHiYoz4OyHv/3bWIEb/UNKlEgWI6uaw5mHkWYE2tvxYSRAUvAQqGDyEU94ENH952EhKYFRB0svyoNQUHDo0N0keaEYEwseMCcESVfUcTa0g02wLIrOXo6Hm/TfPUGMRtcUcQSr2Ln2QOaMXv6uEebAjKVgUOIC0BgOwmh0zGuSKAOYOZMHQKFL4RI2Lv+O8Rua/gB9ANkUrPy8JijETK+oKIEx55Mn3TpkYwDjNaNcRotVG8b/OEzoBJ8UTtTI4IBhBBhTx42NDWdGw3KuJ+zmrRsqeF++WlLC7TIlfkC4BJYnEWIYVxz8lL6nNCqZmnFGa+gLOOOf6wDoFbiE7IA3XQA7Tk7wEHBGg8tnhaMkavgHuSQB8WggauKlQ0UqsgkHB3vyqCDhAWgAMCtisstIZTB/k8KewFI/JOM+FPtcWtae6PKl8eEogRD2LMVHPDz5N/YfYFr0SwBo5HsAqxSCmNiJRStDZZdh4PBypgJJuzN3W4d4+Iznn/hWwyE0HhwY8sMuTl1ESaVWwnLuBWCh8CZn0xYOTkXQ+M3o4gzN1rMQJKiU9AjMDMUDciYYCgcJIp4LjeYqiWsTqMH+Zh9LDobioAyrBpk0T1oEuiB7loTx6VJiEYSnOJIWZwB+BYppyomCxZMSSb+okUXy6PuTa+dejIwMSQeWuEKDg3tF4sUeZe8B+JI4uLwbCXHSE8OoFyxmghdH0r0MXh/esOQ93azYGVlnBlmA2c7S9gQoTlN585U44cbaDoZ7EqqUQWOhZ/qq0jruyrlMjZ4p1w6OCQYJDTGH99YkRphciuw81pzvqagMI6w+jeFmzSRckqeh4UbDFZZGCf8HPECynqhXaVB4A0Is8ACICHALABj3UYwzAW8uCQfIzLpFyQ+AeJJ1n2RpBlab7xXf974GUdJLoknSF3UfhVhE6r2QsAvgF89u9IAQK0UFBlq0Jfvoox8reQSIm7t0ye7f/16/R0Ms7h+Zo8lrRBQjsZC5Jq49NiZh++t7GtF343AAWRXKFFhMZakB7VN0PvbujVwaNDTDJbMSJvZk5qo82AFLkklNC2BmXC4FCTEKP28ayL8oSB8hxyeZlvAaAt6D/IAmDySZ5ZMKcY2ipBZ65TqLam62Hb2AxG5G3zfI8XEPAdDiNVt7QxIlrqdK86Cg8wqw2VnabXbl8qz2jryOYEMpkabYckm8nnyvLSwu2tr6puvqynCO5J/n14ufa9dmgvSfS7kBsgkgaNQddGUiCi136cR2aKKCzww7D8YoIDL30qeSvJAizui+ILSiB8Plsny/eQ7Ac0whpwJMo/ouxQMehKwCABxTckxRXJ5xGQ0kea7MzYpBR24yMjrqTOYglxWnGUVgUAPf97IDTs4i5YRpVMs2PNBvoyND9nJhXqy6NJ5QiaRt7uzbQDAPppQkbjRrNZ1zH7//rj26961NXxi3Zs1NIclETqtNa3Rk9CcSUCC7NIdpzMTmA88VMlY8L5yz1vSYDACqaS6a7yfHduHClO5xnNhjP9KkYRmR+KApw/Qn7PaV1RW9BiAuGtrsD9Y15mY0FwBrJifxbCrJuJUin31Ko4sGMsU+73EsRmy74nOr8Vmp2s7OtkBAxc5qTQUkRBURXFIpNbQBcjWxZW0yZfWpMOSQIK3wbPhz7uAZz1FRQFGlcGKf/uQT++1v72iaggks4gr7EL+K3r5+5SPffP21JvDIvxpVcrOEdWW6LdOZsvd/dFtgFMM665s7dufLu/ZqZds6iJ9OHVRjS899KB49ZriUHmDQ1bk529/d0Zn1R599qrzvv//3v2sBrOx99pMaywBqgBeS9KQIbrMkDUXiawG2e5cktXLZtJuLRk1hNStSlkl3WrqTXKbNGz3duUDS8fNCjeFCSVO1TA/AIkRWsFhGjoDnF28cB1C0m5uAOD61RkzjdTVBGIAAPF4IgxBgWE8MXpkp5vMsLb223b0D7YU//uOfqbnB9BnkmOXlZZueuSTjd6YCIISQV9+6dUMTAeTMfn4j5VSwd9/DXySraYBf/epz6bBzniH7xXPguQfEgrIN9PbY1IVJAUR46OS7ke5s2NjYuMxHaVSUVZA3tNdo9KsBHySFlpdXbWi4X9InTP/ceuuWLSwsaD7m4PBYoCZkWMBTYnuj4nIWLATa+JqkbeOsQEYssIjVwEGmMEgGKdWt63dYF2obGsinFdbfJ854LZf38PhGHUWcZV+wh5T74AcW/C+IYUhV9vbkrFYuWa1yKmPm//QXv7RmtWT9vd22uvLadre27O33/sDq9Xa7d/+JLa9uah/PXJpR0/ruvcfW240fSkNNKPLgh4+f2MTFC4plO3t7MtB+DIg60G9DgwPaE8Vy0XokCYO+fLf8R6hH+Awwtl8ur1giThGxX9vbrHByZMPZpH1yc8omB/ptc33Ljso1O6jXbX5z19I9Q1apMFnbsN6Bfjsunlqis11rJlKRADknrHA/WJPRsVE9Q6rpQs2nRkaauoz80nNCZ3VXfHIy1AfsMZ+O8+Ze5O/GXJrXZ2/rjA7mpZwX5IcQZAC1IS5EIF77gR/05CD84YxgnRc0Kio0/pwE9ulHP7aFhUU73D9QzoWE2uj4uH373V3tw6fPn6tRQQ4MCY2zm+eYaXniDk1jmsVO1MAzxyemffI6SCmnkftbUcxW7kR+EUhTnPPkwr29PaFuIhfgOfRcDgIbpJq4Lu6P4/K6rLd8skIexPeQr0MtgeaWN7e9yc/EHrUn9aSa7oHswp/EAmT/qGf5Hc468szIAOcMak1PVCtOeBCIzv11YNclZ4K2fAdxzGXwPCl3Qog3Khws5fMIU6iWLJVKKqbzEiIs0SREVrNStAsTYyI2fH//vq2tb9vo6KDdvHHTHj1+pMk7ZOioWWgiIGO5vPRa03xI4K2vLNvm2rL9zd/8F1t9+VyNitm5GXmMAIbiEzmAoTaT3p0dtr++aZvb4CoNu/3BB/b9l1/qHLh6/YY9+PobTadfunzdEolOe/DwqWVyeclL3n/4xE5LFStWqcNpnnpDIJNO2shgn/V2ZzX5mU11qiFGNnVaqtr27oHtHxesziRFAOLZD1p3TZo7cYSFGxke1h5jfThXiK8RE2jVJqH5yvOiukasc2f8RwN2TTtwfZLm8el0zk4WH6k/NJmY8NR5FHAYNhj72gkZ7WpW8ssQNXf3TiyX88ZczDfJeWtBBYI6COKQ6r04cRNUAWh48yzQwASDiUbcnEU+Ielr4PmeN2HIxdxPLmX7R660wDPQJg+MuscZ1fReB/FsxDolyh8pd5UHQwTlzxSbI0ivqQnJK/nPRqlANSgCgdQHJ/xZCh3Ic3I/LivJBcTmgprsQe6Xz9bCR9Qw8UYEPxLrtCiT5PJr/l7RSzA2KrhvENLk+RC8/+TPGQhiwomQmQ2ESpqHbzYqPC7G2tOxjdh08L/F6OkySGdkZCeLxUitgOtqAjLBDv6lYYLMSbhnclnsHcXH9nZNCpHzgh+SUx0cHmkdfX2coBMn0WPjk3sd10NksUB6jP5hnjs7SVqE7EA2ZJ+qAava12uKSEaLKgP8PBM0Xrs6xhLr2Oiz8z82KmLD5OzY+Z83KuLPtUidPzQqzm+kH/7+b2EFruT7NHIqcDH4IcDsoGCGOUcAoACl2OFBJFHhYaRYcSmOpkZSY0eZYopimMRN5pjortPd3N0W+MLoZWTKEBQEzuDxUCjIvJGikyQDQDSyVAXQBj1nNBJ5Ty/cMBXscMMkeWF4kyLqz8FAc2kdl3ZxDVghkBrL9mDvoBwJGQeVgxsVgTAUJgAIBAACHwe/2J4aU3ZGK+/Hvzkoy8FfURJKkFSwCka2gDx0PPmcfGbejwTCNVGrGgFHJ1ZdYjM7LZxoXBJQknUjOUNKAwCBkVSKDhis0rUPkyYY08KqZu34LARRCkJJ/MjIzwMtLFkAVpm2akw3GNKGBJxAyeuWSgUx5nQgBiasNNGjhmF4Dd5HAB4BWaaNVTFf0f/tyiLvA+iakRdKSrIjNY39UyRoFDLsu8iQiiOJsZEUzZA4yKL5lAMKJMawib2rzT3R4dh0YBfghukfmfMlEmoCra2v6aDSYRUkrJASYM19fM+lo/h9CphYILQYAIEVpKJT0gbIPrjZksYLYSOgpRkkWKJkVPx9b4C4tm5sVMSGSBwf/R8P+Jih+++cTWHI9BbfgWhiG3xd+G9JmgRWCpqxgF5MxDg7GgaZF0OAGfJL0Ci+AzaSrdGEkQOMfElahIRfTTVfF2SNaDigtevL7swoTT0pMfAmiuufl53t3d0lSQm+/3JhUa/DPaSwVlKMNI8Kpw55YaQ7MVFzgCoa4LLX2Dc0oIhLam4UXVaNZ5AkHDYv9wddbb7U0AtJoYxgA5MVtg0eKtx7jRIrkWbM19lckmugGYRERPCQARxSchcmgBRS8CsQa7/akgWKY+qOxzqY7/fP/UTEqg1eDsTbFttN0xfe8NJ1lZnwwkD8SPFAz0xo3FFgssfKQXKJa4lJIDHDPRfcWExSRJKeagiE4It7xXURd2muys8nFCWeSDo7Rk3KcO00MXk2vFnnu1PscIFhSJ91OBh5jDSYs+Txp7h+9aoKQJivQNViwqAPDXsYCayMS3RQ2CBPRGzs7emXrCA/B2veJ82cURO9G2DcArLwelyPGo9iVpGUuvkmBbmmFgBAwsgvybjiQJCBQQqKpoeKD8WDtNXVzPEJC58EcK1fB+PabXtryzXgk+02ODAkZjAGqTL9i/KHQQoOXXmdW+Ge85lJqmGTRy8N9oZLPRBXQqMl4ZMWzhzKWLFSsmaCvZPR6yHZAnPv3t27uj6e2empCypkNd1DQS+pOkx+MzqfYSjfufOlAIdYUOm5Czr7YBvXb8yK0czn4H7z0HAdvIeeRRoPYaQd8+3jk4LWg3sIM5ufp5EUY4KYRPKxahfLjecJUCFq9/KCmu7CUBtJxyB9BMOOYqVer2jvDA+PiEnN5AzTBIAMsEXxdeCzMe2D3BGfFSAfsgR7CeCFazo4PNAeInbzeSiGiCMU10N9PZJe6evN28nRob1eWbELF2ds76ggcLu9A/buqRf/eBnACmzUpE/++N63NtTfLfkeSAuprm7bOSpYvSNjxVrTChWKQJ/2AkDivGetnEnXtMLpsUAEGiBMZjKxgXQazzjr75KcbdqXkswoFmVGT+OZ++xNQxi07unE3oDUwb/7pIXLPSEDJRZYmCQiXzounBq+RMQaGLmLC4tiJccpLIo3JMm4dvYVTwgxHVAs+gARK7mOg/0DGUVH6T7ACCYY1jc3XM6ligwETS6zcgmpmR7XaE7wmWAOT1jx5NB+/tPP7KuvvhKAzeeHicyf7Nd333tPRszr62uSjYMVjrRHqjMpwBdwB6lMmlpt7Z32emXdvvnugYDdhnx6klYPU1TKHUI+wBnrU7DI8LXZ5Usz8g7ZXN+0n/zhJ3p2/+4f/sHZwVU3ime6VnG5VtMzSswE4NfnTDmLGMCO5iFNPMAUYgHTxbD/IKQwxdKWaEr7PJ3xiVeabYB83APWkufi5OhYEh4QLpAmlUSUEAByChixPCMAtjRHU2KKY2rO/aPxqunV0LDEWJ1709c3YPmeXsmzAeJAKEFO6eXyspj5N6/P2UcffuggTVubffnFFzpDeJ4++sNP7OnDh7a+uW4XLkzo3FQzu42JtYwdHO7alSuXNVXLOtx/+NC+/e576+lBeq0i1rDHn6Y8i6q1hP34/bf0/KvRWa4IPD45KdsAmvCBYOINAJ/KdilJJ6IcH5+IBU7Tnnjz4ccfyv8BY1wmawowlNGTT6V0PmU7M2Le+oQYk74O0nAG0AxVnpDKyOgaBrPO7lJZeT1NrGdPnyjWizHZjmxl8EMKZ2skKfDvysPVAM/qc+GxwsQNe0Ua8AhvNGqW7gSIpAFyaD//2Sc22Jc3q1ckObWxsmpvv/sja+/osi++vqd8mqkMfBbwBSmcej5WPPXzh/34annZRibGrFAu2/bOgV27Mmvzz17IZ2ME2Thk/JhShC1fbVhPd6+YqTSWZufmbGN7216vbcoEhfwAPyI86E4ODyzbbNrHN8ft0tioHe4dWLq7x757sWgv1g8t299jXV39VjgtWx+eVPWKpLU4T/Ey8Ul5Z/rSrCd3JoYIANIZ7HUeewpijybwMfhuNFXDcD5AlIlT9uRPNP9qdeoXprhLIs6wL5Buo6YReSmR0GQlZ+8h/hiSE5zWM8gERnzWdG4Glq1yvTgNrXPQQUX2TrCxsh+//wc2v7CgeEQMwcSds+rJ8+d25coVW1l9LQCfZgSkCSaShodG1MAlt8MAfnJiXHkY5xV72Y2yk3rWmOxhn7u0J1OieIo5Q5tclwZYvEbWTT5qECkCMIkUlK+ne1AEIrUTIIJsp8hiQY9+fHxC780+UIMh2a6zAVyAcwsZoAhaa6+V/bxCYeH45Eg1t3LQMPkQ8xnl2SFv5BCIjSHHGrpUF7pMj5NriFHcQ2q/OPUmeVb5Znij2X3ZmtaWRP7KZUyVs1ubGhWJZt0G+3vs+tU5e/Dgga2sbYo49fbbb9uXX36pxiPSh8RK1pr8bvHlS5lkk1dsrC3b9saq/V//x1/b68Untrezbu+8+7bktYiXkxcu6JzlrGZ6hTWtlCp2UijY4MSkffH555KKu/X2W/bs3n35e4xNTFsq3WUPHjy1dC5vxVLdCsjsJph4ZmrAp2SQcayUCjbQ223ZVFKTTBmR0JAIbbfl9Q1bWdvSZIUlO60iLIemFXkbkqlplzBCM79SUfOSfcRZreZUkDBj4kyejpIyPXVfwgw+Xk42IEYN9g8J71A9Ro2PfGDhRPUB6wy5i4Y75yf5E4oK3GOB4uGea5KKPBWz4TA1zr0/PEKa06fPiTOcbdSh5GaS8tV0pssTu3QTNQPnL2vkKhQQZbl2rks1ejRzDqRTJv1VqwoEJ99MWrOt3Xb2D72eC5LhakTIg45mj8tuCOMKEz6q9QHsoyRHq3/pNZFIXUzvM31Aw0Ov6/UUxBuuQ3VjWBO/TieViUIjXCxU/kyyQFYKsqyaLopYVlRjCCi/6jnOPp55NSIB0D2nVl3XmhALbx67A7qQoPwQYl38bK1GhibJw4RHvPZzzYUz/MJzDF+DqAjgIH304/Lmva9xBNj9d/wzx0YFBAYnMnlNpr0KvhMk6YnxeTyJAt4iFYUgncs5C7GB+xTVXdgzTEBD1gJXoFalXhSeEeShHMdzGW/2LbWY6r5AMGRdY23HZ4qNCu3LMHGiCbQgU0ds8amYIA2qxpZ/lrNAGO91/Pzx38OaBHxF0x1BKSX6P+oamFCqVnzv/NCoOFvEH/72b2MFbg+P2urKiorNyEiGXQIbbnFxUQGBB4pDAgAXAIpiDaa/s3rLYjvpZ8QgdS3B+ACLuNaGbnpF3U4OK5grqZQHXpdGca3taPgUAR1neziYBGOWAMSXAHgFG9fb7+ru1rgnTRSSOwIyADW/T1IU2dIEDw53mg/O4m8oMeL1aSSg5+uMDmdZwhgB+OBzIrVB8uOHSV0Hp4NgzpYlgeYAp4gfGBwQ2w3WKkw7RiLRdKdoiKZLJNBirPT36/1hcGEuin47a0oSDEOIv7M27779jhIhTMxIhDlWBgaHVcSpUVGtqRvO52O0k+tmLQieFLtah05nHYtZJKNbJh+YHvDPy7o6+7xdB77ATMkywbT3QpmcVnIltVqLXcDP+/h2h0Z5uf89+ZytrixLQ5zPPTQ0oiQdBm8HRsCwx5HjkGyXgyw+cuxND/l2cLBJssJPL35WMl9BjohrcMClLqNskif+p+8F9rjAxO1NgeN88Jcvkbhwc8SFxVcyJQMYdBPTUxVtXdmcJTudTcpaK0nhvZXQO9Ne+z00RwDd4nU468OnJQCjIiAdD24vJLxRcd5IKVIN4vhnTORb+XxI9ryh8GaH3Q/QwIaSLqWPp+pz0XDCxL4rGAYjFRaYNMdH6CPDonSWUhk2aDDOogBTgyeA+6xFNPcEJEFGi7VqFSPBBFcSUGI0+TVwgFK8aCqrWROwRuL81s1bii2wn2WKWROUKimO49NTFWpIipUK5SDxhsY+AC6sZB9l1dh1AM/8GffJDJ5pGGd8Zmliy/Tdx4u5prhH3HjcJypy3TkliYB/zur2MXOSEDHO686gpjna09/n9zg0OWGZsBYspIxYMd3uxAcnGbxe/JlwCSOkmABevfBVwRjSFWfBkNy2h9Fjn/DxJk1an5UGEz8Xx08p1BU7xf7kmfGmImAKn0cjyIqt/LvLfmDgSHHhOsdcOxrJnmBvIa0RN13QOY1687xujL08y3F6Ik4tKE4EGQf2HgUDmrJoogMeiO2GB0PSTc/TqaRNTo6rOAIsFrCQ6rBMCnDdpQAB3WgSsK/c/8MLF0BS9kc8D0hQeU3YwTxbnDFqfLKvyzDt0pqkqEnCypsMNH9o7HLexGdIzQnuE/q9mmhBE5hmmTeP1AwBsMbHqL3Dnjx5IomqK1fndF6UqiXL5DKKG+xJzkreP/o5SK4snC8R9OJ7EfyPWs+wDuP5yDkTGwM82wcnxwInKaZZENaHtdLEk3Tsu+29d9/RFAJ7FjY+tttNOgAAIABJREFUWu0UMNw3Xm9nB43mUXkOvV5+3WKWu4QQRL6agEbOWW8QMt2SEcjGmc7zx/lLI4A1XF3btJNTWLIOMAF6caayBwFpOY/9eXXPK28g+p7TFJ0m6WAQutQD1839xliZ9aHJCpDXlc3YrRs3beX1a0nCXJ6d0bQh+41nmfjBmQoLlNhEDnP79m0VMjQo+MzIa7DXYH6+eL5gw8PDav4DBFy9PGMTo0O2trIs2aUHDxfs2o1ZaySStrK+LYZ69GPhc9KQL54c2Ts3r9vuxprVyqfyt6BR+npt3awjbc2OrHXmemzh1WvDPBZZBtiS7EP8rgAr9RmPDnTvgNFlXq6GrZMp3PCvqRg4M3NJYCzTBjQFenr7JGHF2c/Zsre/I9Yu5z/36+7de5p65WylaUMuAqj16uUru379ukBYpFnY84CxAFEjQ8NqDJInXL1+zZ49e6ZzAumKp0+f6DrZizDa0dsHaAOs6OvBmHNL60zcJF9RnO3otBfz89Kg9slA93rJyny8aTW08bszikv4fezubNpPP/3UvvjiC2db7uyqScdkqwNbbTY7O6t7PTw0bKeFI3v29JGtr60KbKoGpjNyTbduvWXP51/anS+/kUwOjH7uI42KpEwqHQxUkZ9oE6APUAvIQiNsjelha8qbgWnRX/3L5zrbAXa4H7F5EnWxyxV0+clbnAFaLtcs15W20eFh5YXyN+hIit1Mfri9uanzDgJPOkUTr93Pr1y39Q306WykuCb/Iy/jniPFKc3wZEpNy1wOMH1XUwzy6CkDBpEDN8RYJwZxHvb05vXzXDdnJfJXAD2SNE0iQeVM7mqtoclTmgVcy63rV9UcYaKIMxwprNgoWt9YddnTrDfQAOTIW6vVkiYqfvHLz+zatStqJh0cHNlv73xhC4vLdnrquYfIJIoNbriNnxXyKciU8FkENqcziu06g2giJQELvA4gl2Tf8nzsbG/b1PRFnwRPp+z5/At755137c5vv7atnV3rGxoSOA3TUmBdKmuD+K00moqN7LH9owPJwPA83Lt3X7WQNxyQDSoJgMRnADnLf/z7vw966O1WCdN7buLpjP44Qcm5wTQmzxP7ivfL9eTllYAXDk2qTCckpYYN9OasPVG30umR/fIXn1lvPqcz5fG9e7a6/NquXbtpXfl++/buI01tkbfl+3oV+4rFstWreJB0qWlBPr62uW7Z7i7rHxy25/PzmqjYWt+0RKOuxii52s7+jo2Oj2kShzO6Wava0cmRjU9M2Mrahr1e31bOTG4u2aVqySqFU2uv1OytmT67NTtrJSamu7rsq0fPbOXgyIr1pPX1DlhK5vVmpUZN04YQxTVFmGizguSCzs4Gzi/lL5rEclIUAAx5BPu0O4csqbPwOVfYB8QP9g57Xmd+W1KNap5lnk3yOfYJ5urURpI6QxIUIErgVLtiNk1ADMX5N840l0Ny0O1cStRiPkvTH2Nf/E7qDXvvrVs6lzhrkJCBpAeZYGNry2YvXbLVNW8UXJjEo+JIuSSTbZyrPKOQ/2gk01xeev1apDZyOgB3nku8YJBjYp+TB/OeYvkGM2rOiN39fTVdiGmvl5f1TJO/jI6N2fPnz1teg1H+VxP3gYASyVSaOqx4U5trVK4vD6S0pvWIVZzHbQmftmYCXQQdEYUc3MPTjlyXCR3yzIgJ8B6xfiMmcV9ivRTNgqlZyHXJLyCh8TvI88CkllRVDdlCz2ck41IsOes7+AZqEAFsoeoMcPZrdzYtM+3R0SHlO3v7BwKq33rrlt2/f98ODwp269YVTc7RnOA9F+YXNeXy7rtv28vFF7a7vWr/5//+X2xl8amdHu/Zrds3lV9A9mAa4+SkYFsbG4rvl2/fFjLNtRJPV1aWdS7dvHbdvvztHRsaHLLpuRvWbh328Mlz60x1W6GMrC2yT+2WTJH3nkhulxy0UuJZbpMPFiQKnl3yOxQKMt15+9XnX1q1aXZ4UpAMFXtb8jXCVjznJM8lR4SIuraxIdCZ3IuGmfsWVtS8Y08hjcw9QK5X2AUqCNZmvfle4RkyvdeUT5hKSLbpjKqVkXvutHw+p0YieRxEEiRfmSQgjkt+VNPJNavhRaap6JIdnlSsO9ehPad9T7MFiadgpk08Jg4AIjGJRhMOAmaiLUiI44/WwzQYTdqkiAMibwSZXfZ0rLd4PqU0AWGgvdM2d/f0Opr+ROJIYD3kM58ijeRBchFe35U0XP6S85T/xUDBv0m2KswQ8BxwhvHfInXWK1YPXnutRoUmqiPh0ye7zw0jGGOAIrqpQXD2d7Aq4remjMJkt+dX3hSJnpve1HP/zYinvIFgthoV3sQR3hI+kDcqHDCnYRIbC5Kn+p0waPyu+1vwpecfAmxoAqiuDlMGei9NksSveI3I0nney+95nem+VXyxhxyrC76SSZcfh8x0fIz8ru9/agO+7z6taU2C0sAQ1hXIU960DaoBkop0qduoJiOMQo0y/xmf8I9+fVElwfeNfPBEMvM6nOZ565OdGxt5c4Lkdy1kNNM+a9Lo3gf5b5QnkJAkLgt3iBLpPzQqfueu/OGb/4pXAI8KTBqlXRu055haINBj4hxlEUj6pFeO5EWqQwBjHJPi0CVx8iIvK9YYX9H0hsMQ4Obo+FCFPUBvNAIDAHdNPE8GxWKRJIYXLVyXxtcCU9QNqp2ZrC4n42Ak6Dy0krBxDWyFSoJ4AOXDfyp5IqEh8PEeMgfXuH4AMhMu50RA4H29MKHwcEaqrjUYQsGeohDlEIKRxGvyKQA9BRyWSkqieK3YAY6eFQCbUT4EcJRknPWSwQ+MynTKdnZ3rK+nR5rUgHMwGyjWkH/wbn6bWAdRmgczKLHdg2EwP8PBKAaOwG3pA6gh5IHfmywOVjtwDkAmwCdoHCIl4BrLPpIoqZo2N2CLX9z3yGqSIVMdVpYnKupuh3tAYYt8QKVet0MYcNlsyzjXGzjB9Dzo+EVWgq4njP7qWmiIUWiEpAIGEkV/NNbVz5KYwZrDkyTle4nmDfcc8zAKWo15RgNgvYebMnGPfdzawUm9f5AmIrl2JNc7+2JWKnGpC1BhfVw30o2X475zVlNgUcAUAxiKExChmx+1Xn1dz7rtGH6pwRHGJX3cMkpFhZHTwJSIDUMZOoeDHektHhm8RmDTUEiRLO7u7gdWAd4L7mWgd5aplz8/8h5oGW37ulDssaYUc0xJuHGda/xTRKpxFdgbDnLTbExKtgWw4vDwxFLJdrt144aK1C2koHjONFlUdHZOPq89iAll1EkVA6eMhAZAT6cMH/lSAyWd8YSo5Q3QFFgYJZLiXnVNSk82FNsSNFFh3qEZ3VBRRXMs+lyg1UwxpHUw2O4u9cECeeLoiW2U94GFK91U7VGSWuIbviHux6IR02CwHMdB2ZswPNQklWFcrZUkct0UaNyrOua9SHNUPGGSgV1gtjiom7f9A2T3kLjzvc3PADpRQEaG+0D/gNWbdcUKeSUE5jXPz+raml6TZ9HZap7wKvkOccPjXbnlAeGx0xknkh5q9ymZyPzTBEGpLFDTG0DOsOrKdNqlmWmxbdkXag4HTx9uDPurs71T7OsXL+a1t2AwT4yPuyFtyosw3lM+A6EZJKaZb+SgYQqgmHEJAoblw7PhHhtlPWvECk3nRAPsWk0FPq9PgeOjwe4tommedErnHKAd/0ZDlj3DlJGLLLlMCK/LOtCM0R4IE3M+AQbTyaW3XF80TOiJ7eNNY/YFLycPpyBRhmSea8ey9xldxwOq4Jrx8dyj8aPfRYs7IZ8YNa2rDevr6dbzDkPT/TJMLM4oN0WMHRzstY2NNYHfMSbw3As0OMGDoahiFjCRsXvwHJo8fD41ergXmhzwJF0NM2lNuxSB9ovMs33SifvAuvLzkCEo2iQhHxi1GFjDbmPf3bpx3dbXNrT+c7Mzvs5IqAS5CMCFrZ1traaaR/ILyAkMYn1g4/K7sNpopqjhWipbFqCwXrHxkQHrzXdZrVLWuqa7cpZIpm1je19mlX5WOmCSQO7QmjZ36aLls2l7+OCuDfb3+f2C2ZvtljRDqdaUQSY/XWMfieTgTFaMYrmwEixGMzX5iRKA2BhPEz/4H4zfixdnlA9owgYTzdcrtjC/4BM5FEXkaJ2+d/hSM04m110CbmGAXpya0v2B5CBJLsVrJwD4NByxwskJAOKHx0fuSxJkJPDsItYANrqsovvy+GSFCUwnXiJHBXlDYFTTvNnU1tQ0K9cFagnY5f1/5CW57iNrTyChVLaf/+yn9i//8i+K4YD2gEjcW8AOfBJ6+3ptdvayXb121e789je2tAxISFPep1kpEiHdvPfe+5rg/JfPfyuJB8pt1j8aH4sVHGKeZJsCSJHPMf03ZkcHB2pkffbZZ4Yp6Rdffh2m0IryHIlsPQAlmKRqNquY5SxkD1ZsdARAGCAlLz8F+Tyhd5xM2tHhoZ4rPFiYKiFWETe4PnImAZ6d7scjsDw0JMfGJmQsTTMom4VxXJQvBhMzNDAAbjuTKQHMnm/jPdPeArEcHEAbnXzbm+DFEmxP92bgftIQpjnjscRPUUmOSmqlqmeS3BZyQUeHF9RuHM2z7Xnhv/v3P7Vbt69bqYixeUZG23fvfq8zqq9vUICzM29hXHaIXDE40K9nX7l4YLYTe4mlkj4Mprvuw1NR7rezvWMbG5t25eoVPQecH7Fp2Tc4Yt9+e095ZyqbFeOe3B+PCsxeaTq7d11CjZAvvvrGpi5e0JqvrW9oegbAQ8ayxKtCMeQ4LpvC80is5vPJByzUHjrTBZS7rJomrDs65Uslr61sxna2t6wBy7ZZt6nJMasUMTzHPP3Ufvnzz6xRr9jAyLAtPX9h66urdvvWO9ZsT9uTp/P2fHHJ9o9O7UcfvKtpDs6CwgkStExudFk2nbLXqyvWlc9Jwo7zfXxkxNZXVhUfMSEH6No73LPunrwaHTyvxB8kfiRfmey0J8/m9QwTR/t6e6yKKXzp1BLlU5ubGLK5qUnbWd+0sclJ+/LBM9stndhJyWRSnUl1yTeimWyzEqa+kgoiT3CZR57tchmPMqYlnORBfqWcSsBUQlO5jQbNcppvNeVE1JTcZyejOdmA3+GaK6Wq+yslk7azw9TZiRqLNHW5R/nevmDKztlYEOv7+PBQe5vXYv/TvPOzKxrkngFZNFHUQOaMk59Zwj7+8Md2//v7ApYh32VzOckiIoU3Mj5q+3u7+txj4xOSwOT+OMDUFAufL2oUnn3qE5cPcw8q9tQ4BKsUMXw5sNzPpjx8bMIBUhq4u3t7al5TO9CQ58x4+vSZ13gBYIuTFREkdNDUPyN/59kh7lPbK9eoVbX+Lq/pEs2ed3me6JMNJhY/v0NOx7MNsS8SMZRDBak9GoUOpjqrX3Uk+QzEJoGQwQNQ5AAnfbVyvehPp9qjzbrzTBs21FwjntGkIImm3ksmTOD5zNS4DQ8P2KNHjxTn+Hyzs5fs8eMndnR4bDPTU2og0SjlPqyurCoWffDB+/b02TMrnmzb//bXf2XzT+5aMlG3y7PT9ugxE1U1uzQ7Z8eHx3awt2ejI6N61g+OT2zi8qzLusrjZ0ONwS9/81vJZF65ctMKxZq9mH9lXd19mqZ4Nr9o+4fH1taZVv5A44L16e/JWl8+ZwxLDg32W4bnsmmWzXXb9t6+ff/ohSXx6kD9oVqzrlzeZXoldwbTmlzKyXYjwyPaXzqHIUBlMsrNWW+aBOQ33EPuDc1nl5CuC+Qldkk9Qb4HPslCU0oKGID/8jFoqkbzhqw3C06PIVjhYdppBwc03J0QVMYDLpvRdR0dIQ0Nqc3Z/5rm59kjz4CQhgw0IpKcrYG4mJD8NpP9TAPSlKIRQs6Bb5xLGXO6uycEscc9BnS9TLWS6yQ7bGt7n6PAc5/oWRcIcdQk8qmU7C1NOSfQ+lQS5JgIYIeOpne1Pfdlwpu8nfoydCU0c43pSIgtoQvu8pNvTFScjSu4yXYciPC/t2SmWw3xUHeHgzpibE6A8+dMU8u/FyFnouJ/3qhQhUIu71XBm82UWGS/8WeQcFLN5/iSy09506YldRV+580mipOJRU4NJGVhadzjMFUmwl7ALmNt0j9w5vlIM8tjXvSI8BrDm1aOd7h8uuNWLKzL1J35bOiag5eepJLDbYkNLE1/hwl71f/U99GrQoll0EsP2Epcnt/fqPA38H8Pfw+/JBI2tUOQGuN5PS2e6rykaUFj8YeJit+5EX/45r/mFbja0yfAgQeLQ0FJYHePEkGmJlQ49/SoI8mDPTg0oGeHcVWx8ZtNBz9DsYDZ38bmpgIS7CQHuLxwRqqB0XxpWmpc1cesPWC47IxkiyRl5Mwayf6ECQoKOGnC85piRzsDmUyRRAYGCoU1n0GjgDAzUimB44DrBBk+B4xrGtZcI8msGxE5Q4cElcRDhmscRgFoASQk6DkA68GDolbGU9JMd+kZEq0YgNzw2aWAuE5nkzoIIDYtxmahAxsTNJjBfF6KVgLyNMzIo2MxK+TZoYL/WOuKISoBC/Yxr6N1l962a2+LtejNcO+Iyyjax9pIxmEq+MELG8YNVaOEE2tFkiLQKOjPa8yaZEddbmf2eyg9SzYlj6KxvoT19eSlY02Bx5eAcEy3YH+idx2ALF8jDkkfrYxeDNqT4SCJRr+AvYy+xcNOTJFgphbZAtxjWCPsSe4XUhB8j4QxAio6ZFrSNxyaSV2n2HBiq9QExLhkkDc9+B0HGJEnoiHmk0AC3yhCAQLLDqyfsSO8mDj/5SOVrr/oWrpRBsp/6s0f96ZILJa07wIrgu/JjyH+dzAFl1SRGJ3h0G13k3uNdaOLHMBB9pV0cMNd1JxtNDRnFB92ZrJTbGvWnOdJI7kwJ8NhDMNFmrMMwAczbkAMZ1DASAGI9amXKD9BckziygFOUdXT3S0d8p3dXYF4AGOYiZIgYlbo497RAMybVN7U8skgb2AwIdRuyPcAwFGEnE0xMOnFmHT4pIHtEhMBb8KhHY12qTd+AES1TsFYjgzOjZxdOsAThQDAhmshLgA+wOrZ33fwyWWaEio6HUT2aRreA2CZZgHPtBLn4AHhiW9MVhKSiUNfGAy9VKqJccvrVMmsQyrDcwNbbGtrx4v3avBHECsbdrYXkjw/gP1MOwC6ufQNjFzYnlWBXpJwUsPS5QE8efQEN7JOYrImcCBIIrSYNmrgOWCnhJL4gFm4GMA+cQMbjILk+rUr1o1ZpgoaYpkDpUwpaKqi7Bq6K69XQ3LZYRenp9wLxLdcyzxezxLrzZhzMKFl6iLGOYFtQUcU8E+MqzCqq8JIjXFvTPpzRcnlTRWe9TiFFhsOxGOAMZq+FKcyvq4jZ4IGe8YNWZFRkG+EryHXxR5lzXyCBEDRZQmJOdLJrVa1h2GyybNJhWdOYIXOFMbqT70JopjZxnRINvjJ+PoCysuvmn2qegmWdNADbuc1OjQhye8SPwH6mUKJBoxMuiwtvQrGn+yninTod3f2bB+N6gKNRaYe8M+AUeRnADGdT+pFnO8fL5CCib30pAGVTCBoa6JLklLOjPLnFka4T3F4Y8vN6WFRT09PSwecZgNeEpxJe3s7kr8i/jJdCdmCs5uJjzi1yOvGxiX3R0BJKFbIE5BVqBaObLi/x8ZHh2xjbcWuXr9uHR0ZW9vcsdXNXetIZ1tSFuwfAHXOxUvTUzY7fdG+v3dXzEFyIqSwLJFUc6OGV0C5aielil4DYFeLgIRHYI/CPkRfeUgSVQ3LinhRtvYOb0zTbPiDP3hf95oYzzPOmn31xZe2sPhSBToAOE0N1iHmO+xNQFSA+5mZGZFM+F1ASgzV2YODQ0P2avGliCbsK9aGvEV6+khzFt2jZWho0OYX5tWwRYKI/yP2Dg0M2tbWpnJFvsgDaH7JW0u6xx0yiEXWaP9gT3GGidCuTD4U9LBPiRWwAxnkrNu1a1dtcfGlmmFIuwGmEC+5t1wLoBLx9aOPP7bubiYNdm1xYUHPTmQ8sp9GR8dtbGLSHj56akvLK9rj0jH3wzTIj/r+ZD05v9hvNB3KhVMZ+NKo+OWf/LHe88uvvtZzSmwDiHTw3L2ujD0aJAgBbSTng+RaaH4jiRUPeHlU0KRGMqSzQ/kxvhicMcRo6UMnmYJhTX0CmQah5+PHOnNL6JmLMAMZxQk4gGxtbXiuAQodBUapn1/cr2I4M3lQ5QsXdJtFEgqxXDmOGqI8vz7dRDOLtROYookYJgaS3sxIu6cVJB0AKhr8NC7K5RP75JMP7PpbNwXAy6sn2Wkry6u2vb1n3d29konjdZx85GA+YDlgGc8w1yfpJBooIWeuYORMg5FJkUyX+291IqflsYr4SqOMa4N1m+3qsXQ2Z3e//97KnDHSKW9YTy4vYlRPd17xFUBcfnYdHTa/sGjDI6P6OUzm4/PGOaCmSalkB5AlGpAisiJMaXqZ/JRYHmQjiTk0qjkHIR5pkgYpmwDKDvbB5j+w44M9+6v/9Oe2uf7attZX7fhoz37yyUdWLhfECkdWb3Ntyz76yaeSSXn+4qXtH5/a0WnBpmYu2ql8/cih2Us0zdIyen749InNzs3alqbfijZzcdJePHthA/m8zV6a8YlhwweCHNfPPa6HzyCvCAyf944FqLMHYHBiHbC5umLNWsXGh/I2DJli49Dmrk7Zs6U1KzTrVqiYdXflGF1S/MFIG/13yTMBPmZpoNEgCrVAmHjlWeLzaho3TCZFoIo1YOohyh2RS/rZndTZyPozjUYTg9jDuYq0HBJ+nJkjo2OaQCEfS9KEx2Pk9MQqYuV7vcREGQAQ9zPmcKFnoWc55gTkdWpcNRqW7kzan/zyl3b/+3u6T8SWdKbLkOSi/qSpiiQhuebFqYuqrTmXiJ3EK9b80qVLHntPTnQGsrf5ol7jPGSagn1Gw0E1mzTuPQfUNAPPXa0qIJrcQmbupYpAY3LNJ0+eKvS4pyP5hgPXLhUafcn8MxPzmYqL0n7RFwTCC81n/rtQQBIlAnouf0oOjp8QMdvlSBwcjWQ6AX1M/dZqyvk58yTxJJ14Bz55f66L6UkRSALZj8+nBhKTYEFKjftNkCI+AXIj/eTeeT7JC6gHOZIp3smxERsa6lejB38mfCCR5Pryy280qcPEGPfl6twV/YkZOTnSjZvX7cX8C0tayf7qP/+ZPf3mN9aVTtrMzAVbnH+pBtiV6zdt5eWSFU+LkvZioecXXtrQ2KhNzTKRyfq4r9jS/LyatZdmr1mz2W4PHz23bFfeqvWmPXn2XB4VyDch5aSmG3lzwmx2ekJTV6XTE9VMuUzWsrm87R4c2pPni9YklyHmn5xIyo86AsnXCD03a035Qg7294eJIZcE4kukupCrxSYRt4NJXK8FXDWAmjjiPpLlCZWKngmZCpMT+WthYM4ZKuJG8DUjB+e+SDrHEnp9NSrqdTs6psGXtHQaUNmbuzQCo2yVJm1plmVdzlQThXiLJv2cI+9h0pOzR1Jh5XKLACpfQpQqonE4MmLU1eT4bUk7OKIe8vNHigeBlBQbAqql5eXBOpw1LFk7+a2Fms4L+FhRq2qVFBmkEz8zE1aulay9I6hEiIAYQGkZlLtqQ/zZyFeUdJCwgTOps4jDqK6PBud6ll0yNoLzZ42KgBW8gUa8gUz8nkaFE4OVLoULcl7k75uoOHvNWDty3cJ2RCb0mqrlpxoNvf8/1+X5Cp+TnCria5wJUrcI0sRRsp1rdDzAJcBVY0E8jN4jwsMcE3EvVMe7iPVRNonvu1yWN73dL+esYeT3xutgNfFpDII7MolUhRQFYTt6hODPSIPrDP8534g5a1Scb0zERXjze5LjDtJT3KSoXEO8HxwelDcdzx/nww+Nit+7wX/4h3+tK3Cttz9IIbjcEA9Sf/+AEhSM8WATtwBKGJOdjHq2KZkjIJBojY2OhlEnD0Yy2AXcxgSp0+UvADaQNlAx4oid2F3S/wv6fQAezob3xMnlWhzoJ2AQxDmkCHf8Fk0JAH2BzgmT3i9JLKOzJHkaswtgd5wWIcC4hwNGuIDMbh5Mgg6jDGa12KrhwPFCDgaBe3gAoAFISWqkNeJHgISBwwHdVGErYDT4Y0jXOwRF9wPwwkZ6h7AYOtO2s7ejYMkX4/muXzpkT54+cb1jseDRY/Xkg3ukiQSNPrbZy5cvZVoNY4jEl2ZG1N0DTG+xJUPjhSCrZFbgT2fL5yCyfGO3W5MOsK7DeLFG5cI9U0IZutlct34nyNvwcxRlNCz4fZJqQAbYajQpJMGiUU7kaFzr1LXkfZQ5JlD8jO6PZH1cmkEA3Dk/BdYnTk8QwEn0SVh4P4zhZbTZbDowLO3XY7EWAZMAuySVwAQFgAzMwGRShSmMQNhMc1fmbPriRXv69KkOPq4P8BMQXkxhwJowYcK+4BlS4yVqFJ4zyVbh06RAcBZRnN7xQ/dsRFDb71x/IzYqYlOCf1TDI3TpHbh1wz2Bf6qf/DB1mRY0RxM2OTkRfFeQC3MvDSV8oEPtDjCLXSCzKj+U+TcxdiV1kdE+lVyQphlqGq+OyZtAjOD9ouec61RKeMbIRx4E/5Kjg2PpUnMfYBULmNF1tEkORex2sW6DSVVgjkTAXQlPwyWhJJ9WZNzTD/H4vNOUxBtFhvSh0RTZ3W7U5U1P7UU+twzXHFxVs0oyIYyQO8jAWh2dOFs5ShMoicCPpz1pp3jH9PfpZ5AVk/+LRuFdxgUg3O9bwnp6AJ+Z0HFTaBWkNZclQRaJe84+Z99S7PJsZbuyoVh2Zol/dsAiZOXcJ8M3jjN6YmIrFkqx5M0f9O1hcbeZAEkSvX70svEtYcS16iwoL9J9H8eGRWSnsJaADfwM4JhYTg2AYAeVMILFUJn9g0GzZIw0Bk/RxX6hCGu3t9+6JZZxQVJUJcvlsnpdClJiLWA3herqyprtHuxLkgZZG5fEorBxaZw4CZHNuPmqGGShgcszH9ngLl/n0xuMs7kdAAAgAElEQVTEByWb55pC0js/dckcJfzmawp4xXMv6SMKLXkolO277+67wfOFSelRw26p1srO+ikW3TS0aWoMuQeIy4u5f1Kb9fbm9TwBdkq7Oewl5CtYYwxRWRdAN02/VBygg5FGU8BlM5CpcsAGcAaDTooy6djKNLApIE9NQ8VPl4q7cfOW4h2vE58h1p6YzrQFsjtcsyZlGs1AaECGI0oFeuM5TuUQCckXiA2SImQjxxglST/0sn0yUxrUjP0HLyXARK5J53o+7yAH0y7kAsGvhXsNWx9pC+I20hYXJickQ8N7jY6N6N4DJuOnk+5IaQoh5gH8ydoD5kvORedwl85LTR4WjyxlVRnXjgz0iWlNA291fcOqzXY7KbrXAgUt8eSA/Tg8KLAP1irnPvccmaT1tXV5SLmUYUNsZ9jvVeYvkh2WgU1LQ8YaAg00tWNNsWDzuaxlmPyjwZ/A+NXH5pkcmJqalgQQe1beHrW65CdeLi6JdcZzTb4GAK5zUAWU+wqxd9iPkxMXNEVLMwumLQDt9s6uXbt6RXI/Yr+GSR/uCfGZCRUxymMjOdelyQAagQDnTDgMDg7qvtFg4/wFgJLnGEA9HjvHR2L1c2YQR2FSZ1I5q0oaLCUj7GoF5j6SUof285//zL76+ms9F4BTTNnx2ZXT4R8Uzm0aMB9++GMbnxh1Gcx6XaP9xIylpWWV1/2DQ1qrV0uv5Tmg4j0ZpqSI/8Ggl7juxBjX1oaRDktubW3Nfvqzn0lH/s6dO2pwianZ4RNHPJNIXLBH24IcQRdTI/W69ff1SK7JySop949SrK+67EYBuUHPvYnHAuE4wzo7bWt3xyc/kzQD/ZyK8piamGQ/yVMMCY6qFYoVSYTw6GUzOZFqNKlWrWgKgecNRnnMsyJJQpPNErZ2oBCAk2sgPgE+xoKevUL8INdmfcgr45SpF/ig3k3tqcEBDNAb1t9Hg+1d6+7NW4OfMeJPwzY3d2xv71A5K/skepGpHqj7ZEkt5FXysgu5uhp7xFXMegGmg3Qo181/Q3Igdoj4JECXSb2GDY9NamLz13fuqAGBBFxXJmud7Un9T1rTxCVNJTFxA9t5wWYuXZIMy8bGVjiT2xVXRDgSkFwRGYZzToC8ZELxwXMwBeCPJtuVuTmRsHheue9Npu+adetKdcrnBnPqv/rLP7NMqt22N9fs1cILe//HfyBiAgDxo+8f2P7Ovr3z7vt2VCjbsxcvJV9WIkfu7BTgx4RSpcK+ZZq0bm2Nuj14/NCGRoft4OhETFi8KZYWXkkCdWSIafiC6g9qKz4n0pBM+mAiL1AZmbQmHgiQXYS4WjbdaRuvly2TTVl7e9PGkd3d2VejvlCv2THnVLrLOhKd1qy6WXN7psMuX52zmekZnfFkWvypHD/4OXGeeP4aJukT5lP6R4e2vLSkWmhoeEjycwD3nL3Kt8M0OHG0ra1pu9sbymW5T3pGE2jpF21za9e6e3rFnuazpqmtKhUZiEuWK5u1tdVVfUz8XRwcFAzpWULQ8/ft6M8MYCrX8Jd/9h/s6HBfdTNxFEliJiuoSfv6BzUhz96YvTxrKyur8nbkv6mluVaec/YIZ7KmKOTX6HWnS705CxjpYkmKMM2UybSmMvl9YjDnCc+8JlPMfRD5uSdPnnlei/dcmED1qWAn1EQ4zoHEps4GYowUFwSCZZR7MdHv9aATXWg28Tk8Z2roLNzadtIcORwkiyiD6gCwkxHIy8UQRlZW8lmuC8/aep3uZCBiDJ+L95S8oTzTfCqHuCqsQc8teXgwjrY2MYyJY13plHW0J2x6akJm9UhgwaanUQTp4fPPf60zZ/ritG1tb9vspVl5lbx+vWZjY8N2HenDF88tlzH787/89/bsy19bpjNhl67M2rP7D/X5L81dtfXXq/Je4ffBOo6OTy2ZTtnY1EWbf7lgt9//kbWx/uWybW3sWFc3ZDqzV0urlsv3adrrq2++U35R5n/e47F8d9byXWnFiKG+XoH/kBiQbxvDfL1StcdP5y2ZztrB8aklyHGZbEMeVfLRToJqNlSpSP5RDbYgH+rENqYLaIQXXFYWHIapJnAP5eHeKKdmVD3GMyFcxmt2B55pfiHR5goN4j42E5bPuZdoLktTv6Qax+On187gHUwzHxyXLd/N5JQ3ddT85ZwM5tuakK1X3AScyQ1yZJEpMgKL5cUgwmrRurPkE0mrQoBKuIY/IDLSRTTAuGbep2FtIpGclMhLxL7UZ/amBGeqk4wgHkZSkMBnmPNhollNGviyUq1gnR3adp9Wx680bRTWsFRGYjrKOPleDwVlS1XCm3aRZRq96s4mKsihHTuIkxkOWMWa0dUZYv3nZIxIwjsPlr8Ji//uiYpIRhPViskO4XVh8up3AJ+SrQrgfAuvCD9HHufYhl9frNPPv0xrPcLcRsyNfHLBsaEoqxsbDJoOk7wVU18uUUi9q7iCxLt8/8C7wKwivujkKL5ctcWnPNz02htCcSpFSgBB2lkTZQH3Et6E51/AQKm9dF6Ezrbi6//vRMWZxNP5dXiDWHkeCwrkSZGVKhX70fs/su6erGKkrvsH6affsSt/+Na/6hVA+omClWI2yjzB3OMBJIFylpLLenjB6Y0HCjeCkDp6A4Mt9opM0AjKAhoq3tmvMdZ3KHNc2DRixdMpl7ZeaEYgq6RGBUCa+y24RASFmAdjDigOtNhNVGKJBJAATVOizfg3bHoCz/kGC9cqgDXoxhN4aCTwsCMPERm1HFYy7RJLGgayGy/DaooBqAVsAwwHfwqKdRI5mKti2Qemu/tsOJOdQKsOe2ieiPEfjMIwku3p61NSRrGLrjgMO4Ht+R793tbWtsI/ZnmwcjnkGfGNzHESLwAHFkP6lDKf89E3AruMkIBPQ0ebNWV9KZoAa6K+v3t7OHDGdcVRQXW2w+hnBM51XzQ65zrakmQKxQwJPAZbJD8AQ5IMY99g3is2MSNswZwpMBic1cHBDuvG105yDPI7oFHk8kKRCS6JCXSiMV4O8j/np1j4OxJBBHHkhShOAQrGxsdtY33dC9ucSwTFJB6mHIDytauXxV6dmJiw1dUV7XkSj6mpCwLwmBbh905LAYQKZpqAhi4jE5sGnkDE0Wr2NiC3d+sFTQZ2AtI/ZyfSG5MVPnTRKpa03kEOS2zs4B/gyZUnRgI7kTqjGRWM3km8kBaJZ2fUB4YF2Eg465/nTQC+JIycNaPnEL4rMkuAtQ0SA5LCEzESYqHj+8CLHhI4KccGbw8MCNmTKqBqDRsfG7f93T0d9BQgjMqfwh7kfqjh5ckkBQf7N46Ys+YyRQymoIDA/BvXxb2LTTiaFDQfjylWAyil9Q4SRUqWYKx292gaS6ZxYjnHKQIf6ddUVbMpHWziGIw8NVqDZmjLcBG5lg7MXHtUBIuZowYFaxcmyGoA+26QCxsXkENG4IEFIqNo1q+JFApGdgUVenwBFIrpHDZGnFwhrpIbumGXgzUkZ858bde+537EqRIAP4peQBLuDc8vUxu7GPMeA5q6z0b8fEocVej4tRMvWFff066T7PvYS10V0JjRC4DzZqZYc8gpYQAN01H60027deum9iOa8MR+pnW4ZlgwR0cwcGGU1VQcw5IEhGIvwupkTSk1pE8cmEmxaIqFFbGc+0GDR75F+A0FlpqbUeI94kmuTNNgk8JY6+nRPhajDIP204LuEesCIMnrcr7Ja0Om7i7nQpMCwJDrIzEmPvE+AlDDe7PerAPLxaRXZAFyv/ksUWebBJ3GOe8DABYLRMBcij72mKaygseMzjyS+RKNEljNFQFOPKsAw0zIcd/cILtT3lI0WNVIZww+0S6mP39OTE7Z3/7t34amI0CsT5axrgBwAJ58CTDQWUlhysRImKqQrJNLnQFEKYa0BWk55RI+ISGWXjAZ5DWJ4VGzGlBbGu/hLGAyhOcQpv3ezp5YjzMXp7S2gDvcY6ZDWVeeIwpcsctDgcg+5P3E4K3CNGXyaV+sSb0n5sdWtqG+vF2evqCim+Y/Mgqr23t2/+Eza+9EK7+/1ch8+923bHxqygonyLXUrKu3104PDu3ut9/psxweHPl+Q+M50WaHxbKdwlqm0SDfmLKYzHrWaEShvZ0w68E7C/A0CVBYke8VZxiTCADvrDnnC/9jYmJjc8t+8+vfiLnL1/rGuvIyCCfPns+LTMJ95gxjIsHZWZ4PuYzevuIba8Q+jZKInOc0KpZXVlQAXrx40Z48fdx6Dc5psd6DHrRYkDSPMQhmOjE0WxWTy0hcNQWk7e0d2cjIsPX3D0pLP5JBqlW0uLnnTfvwow/tn/7pnyThx3nKXmXyQ/lqmMakuNzdP7JMpsPy+JkETXmeF6axOO9glsOkprmwuPBKuQXNNHIcJgHwwdFzjuwQIE0NP7ac7e3u2OjosACZpVcv7ae/+IWaub+9c8eBS030OtPU8xWAwgGXSiJPhRGu/CQrvw+ZpKfTWjskw/hin0ZyBzEl+kLhp4P5Mc1eQPMKTUmkRQFMAps01Yl8BqxhPkvRLs8hCzasfYfczff3Hvrzqt8N3lE0IQIJgXgm9l84owGdWE+Y0r29OfvpTz+zxcUFge7sC01CccaQM5c91si3Ke2Nas5ogHjJN5ETNpAMKdjW1qpNTAzb22/fUgyVBKm1WaFYtYUXC/IOYuLGp6SDpJ0aGk7koOETjag5byQpx+cJbHPACc4ETVoGkJV9Ry6kCVok9zrTAuqnZ2ft6YsXNr/4yiecLWF5JCJLGPzSgE5atjtnx9y/VEaTRM+ev5A3y/z8ou3s7LVqAiRsIAh8+umn9vTxY+UP1BWAndIMV88m5AnNpv3pn/yp1gmpNtU9TJdjgo5EGIBf6dT+6A8/tDQTUZWC3b/7rV2Zm1Xc7h7qt29//YUd7B7YW2+9Z422Dnv8bN72Do/tpFS0yYsXlTMdHJyIXFEsMsXRbblsyhvvuS57sfhSz8D42IgtPF+0i5MTlu/u0gTCxvaW3oe8HKCZxKvMVHc6Y5lMTs0KJmEAdgrUcUzaVEo2OTVhuwe7tvlq2Xq6sgIBq+0Jy/b2SNYmlUyZ4RXQnrSjwrHVmjXp+Uc/FNaYM4d7BFklTr9x1vB8SiaYeuj4SD41XNvVa9fUCGCaRcxrJBrDVAUZCLGgVDq2oiaVOq1YoGlF/KlYoVS15der1t3br2eqCkhLXdZM6Px3xj8TlTVdk7O4nVDlGY4TrzSjiGwNTSbtyYZdnBxX7OIzMF22f3iocxfG/dDwiLyAiHPEUIzsvU6t2MnxqXI7zq7Ls3OKC2vrayLeuOJAm2IG8VINCIzCYaYLLHRCEmd/lFF2QLmqBgPxgfyH2IHsHzGjUvUJMParwNUgoesAoTcrqZc1iVcoqBb1ycsOm5icsJeLCwG0CxNWImU5g5scS3Xo9qZ7xEnGGR11bw57nujAoPwf5UnipC2vL5mkdTINuWbMH2jwen7LFDVxpdICFVvkDkgriSCFS+2e7LAiOSMypMWi3bw+a4MDfXb/wSOdxRAMuN9MmnDW4yNCHjEyMmKra6u2soJU04Bdv3Hdnr94ZigK/sc//2N7ce9ra2tU7Nrt6/bi4SM1Qy5dvmLH+8d6PzyTmEJb29iy7r5eG5udtV/98z9aX3+vfG0gRGV7BxUHXz1ZsNerm9bRiXRtmy2vrFkKiVziPE27Rl1+XjQp+nvy1tudtUqxqM8EwY/z6KhQtI2tPTs4KVk75s8C38VF97otgMLFgkvkqRaPEk6BHS4z4qCQQIySDJsksmlyY2hOTgDYjmqAkzTBXoiX1GKSwGaKAd9SeR06IZXHhoYFsR2pVxosnLfEcCbmiJ86c5s0L8qWzjLN6JPn1N41OjnEHknvUjY6QRC5UccPILuQvxzqWsBFIL+Rf3OOl8npMh3Kw6kTM8hrJ8PEdZCARJqTs4g8VL4LbS4hrFxaPnCBIS8A3v0WJEsV8l/qKEhfrUYFrxJUN3hfb+447sL5x+Sh71PH888TDqP8kDCXFuXeR/e9IRumPcJZKWJvGO2PAL8mwcHTNP3h6hd+rjqm9fu+RMs6J/2k2xDr3Eh+C1EwNm/PDxvE140TB/yMJkOiZFUgAAqfETEjNL+CVLZf/3n8w3Mk1UMiCbvfKvloVAHR1AOxQpNXBZHakCbUZPUp57ET9oSJaPIs+FKG6XVN/ZfcLD6S7eIaRdyLeBTxpziNwXXFponjMH4ugBcQn6MksbC/s9GJVgxUHGwNapzzojg3vOE/E2PmmaelfA5Ds4za/vLcJWsmvMlL/vlDo+L3bvEf/uFf6wrc6Mccb9dliIJhKEw+Cs211TWBZchAocVNEtHb16OfW19bc3+IWk3GUMQXN9Zyc8/IPOF1SJZIOmHD8fAT0J0Z5mBqBKcVWL2fHQ5Sxsf9UHHwOVAMgvyNSxihXVht6bVTFAIiA+Lxehg/+WhpGBXzJr8OB7Et1YX1ziSgpQ4KLkidUAdinBjuGs4ySZUxlDOveX+AK0BRgBLJpkgCyPXIY2bmTOUzbT7AdTFEu3LOZgc4qFTs4GBP4MUA45LNpr148cJGh8eU8Ll8j+tOu5kafExPLiUXIk1Sb+jweUkCOWxZQ/7dZZ98rI0ASBIj9iSSN+d8Q/ie9NlDgRr3dpQq0uEYoGjAataXgAlIzMEg3W8aOBjPUvzJbA2wZdDWNze0NwRwhcVRl5sDNZgR8vpi0CVcqkoHdGBs8Hl0n8J0hczWxAhxYyuYRmKK1GoCATi8JCWQwajTmUqsozRrZdaGvJWbQlOwwJBC3mRmZsrmrlxRo4c1e/70mdbkYO9ASdDFi9P6PUa7MSY7Pj0RsCpZAKR3JFEAC8MPUh/l9CSHRoWzmMIKRMA7eHSwLGesgrCFBBA4C8bZMWcTFf7z/v/0f2LA+z3WQd8MCSvvGRpobu5FAslIJY24klXqFR9rD4wQ7qGmmcL1+6ij2a1bt+3+g/vSp3YpBgprLxzi3lJCFRIMCZGRtIREWI2KesPyubyAVPYrLFyxgGoVfxbQMI4m1jWuwRuAaJwKGC4WpafMZ3TAxMHys0QnYcPDgwIWHMxGy9qZRbGZ47JMbdI9J/65nI6bdnly55JgIolyvfl8yyw7MtFiwiogpVZTjKA5RCEgI2XkQHhGg9RclFbjWsRACjGN58T/zeMAQQqgkiSJgpaiTux8NY182kL6nnr8aRjXbXjEPy/yehTd+hnicmCJUOzxvjDPZXAYnm9iGMkfICjx0huENBBbqafeA7aaGHRJnheX6yCuqbgnCZRvTngWg8/P+ZFkAEY3Jm9YdzfnQk0MPZok0rCmoZbCZLbopnswwrI5Tf2gxc81iPWqaSamHErOdmrHA8T18dmLGv1tuBwCxThmycQosbySroMsORZY3kew6WH++bMqg2pkG9LuaSH5CRocgd1HfOH55vU0ARSSSTkAKQGnsEGyquya5ej0BoZNXE6ANWfE+/Mv/eUg1SCmI83FIJnoTaAA8ssrh4SUJNknBvni3nNviS28nyYRwhnJvtR/J4I2Lwz5/l6t/dj4pM7Azk7Mv/GaSTtw3Zm2rnyP/dM//3M4bwAcfNpP7GzOsiCbxb1XXCN+B+kY7lFkOTtAHx4B7ffgQxSkviJrieczToL5GccZS8MfBqhrAtMEBGDG2wbWKzGDCTFiNzISTLXs7O26QWSUHUI6MsibxbjK+8R4zPe8kGpaPpuyevHEenMpuzQ1bu3SEW5aRzpjW/tHdnRatuPTiuW7+92nqlK12+/csq4cTEGftmFvcrZtbW7JU4Fim6KVPUcRX6g2rNneIXk7pirYt6wVMQ2vHk4JvDEouAEUABp7enN269YtnU+rMnYG5C3ptb1pl1WBRrMCcOjZs6e2sLAgKQv2Ng2dCOZx73jW2Ueb21sCVdiLUWpS06nIKeLLA5lDUyXdAs5YeyZa1miCDA46QxEmsEw4kXnclcwIRsbkQpK0Y4pGxXrFjk+P5Y3CJAObolZD490LcAiKmHM26mWfxGw3+/jjj+zrb75Rc40GBa9PPON6kFGBrew5YNr2D/c8njXIGSLbkM+Rlnny2Oi4rh8iSyykpesb5DhhLwvsBkhAyoWJinAGEWMART/5yU8Up7797m5gWlJoe35CXOEZ5sGV5w5gBl49yaTuI/kv57BiQJjuVOxA3gxD6AKNFc8diK3ZrpztHRzacbEg9i8kHk1WBN8xz705F9Hx59kp2a2b12QuTGNifHTCPv/8jsB2pkB4XabDOFeajdgMCLJc8m0KSUSTeI4MU9V+/ouf2vDQoP23//u/2dUr1wRAAhyrEEf/PEiyMRnFc4rx+ObGRsgBmFBy5ujJCTJ2O3b79g0bn3At/k5AqODjsrq0FFiMgPowqt27xz1Xgv9VwiSfERslOvZCTGddmLJgLYh1TBb4RKtPDvKafG5M7EuVqvzsdnb3dO+I4OzT4cEB5RQyJG3UrK0zFUBs9y5yuc+mAGbWnedcecv+vvVCYDg+tLGRMcU6tO3ZPzw/yo9DXTV5YUrNU3JEdPTxIKGuAPSvVwrWlUra3MwFuzA2bN35LtvZWLVi2RnOE5Pjdv/uQzs6LNrHn3xsuwfHdv/RM9vZZ4+U7Or1GzIIf/Bo3ibHR61cdECHqc2FxXkbGfNmJteCzBV7hrP3+bOnIlj5JLBZBokqmhBMOeEJVMITLO/nMJN7Kdd+T3cwVXJima60dXVnLd2etIPdXcUtpLWYmgZEpWnieyZliWTCtnd3rKsrL1k8wGBek73AOc1kCBNa5Pc6UzRNJ3U2XYvyjXpdTVskcTkTll+91LnTncu6ua/8QmDVV1QvSqLo1IEoNdsTSa3Z3sGx1g0zXa6BmAqgTo7lBC+Xho1Txdx7B3OdFERj3mUq2zVBRV07N3tJ8ZncAW8bcj9iFg0IJrr2Dg60R5EoxKOCvIe8E4+fWL8wlcl7QYIqShXASVrsNyYJOQNg+0cyHHEGYNhjCXkBk5LXNbFBXcqGhHSBt+Hiy0WRihzkC7VgeP3IIo4ZH7n75IULui80bPnc5BJXrszZ/Pz8OQ8qJ8fo9WoV1X7ECa4/yuEpL5LkDhOC3u5hncmT3QvNz3iuS8zlkFNxDZHx7DVIZJZHz7QA4rWhIe+sfqYFyNeIoQL0eF8myKoVu3J5WtNEyCRu7ezb9WtzOrMX5ufVkMGvggmNi9MXbXlp2bZ3tm18dMymZ6ZscfG59eUz9qd/+kf2/N7XZvWi3Xzntj385jv5B81ev2HP7j3Q2Td9acZ2tjad2c/UT0+vPX76VD4aTBTd//57uzx3zfKDI/biybzt7UPIwdyd6ZsTeSY029qsXEMO6UheMROjw0YENzxe8GXTdG/Ost1529rZs8XlNSBlTWNA/tP9gpxGLp9wKa06Zy0yoch8lkru3SXSCqQgfEWR2kzrHoFzsI7Rv8tLSZ+OJtaT+/B7nBWsHc8lcm3cR7CKOKnnRAZwFEhfYEQ0LDLaC8gh1srFQL6idmdyMOHSi5oOT7txdcAFBFRj1t2VbU2GUysyMYU5OlOQmHbznPI8Uo9UajQqHJwuFlwtgXOEGNzEyhxPn3LVTgtlimFrynOiKRKXs/29MeB5op6yQAr02O4T8j4J/Kb3g6PzHkOit50D7trHmIIHie7zVWvc5/5acaLCGw0EaOXCUmrwRkYLEwiVr98m/z2enVhjRJJTK/eJD/obYLhfrwh2oUmh1o1GnPwXvFUb/vNc08ObIOGaw2ucewsnrAQ8gjWIeAUvFkm953oUYd1c+onfVZ0RVElovHKuU2dIfrtRV47FVM3RyYnIRcQUajveh70f5ZiijLSaEpJ29wlc/4yOQ1Hbxc8SsafA1Qu5o9cLkqtUT82vUZ8r5B2qv4KXrvRfgp+pNzSc4KfPxUQ8HiahKSYySvTmEUn3/2XvPZ8kPa8rz5tlMrO8N12uvQW64QgQJAiAoNFQM5zZVcRqv+2n+e82FKOYlSM1lDQiRQEEQAJo7211VXV5l+WysnLjd87zVBZASKP9tmIgGWB3l8l83+d9zL3nnnuOMUmT0cTUSt1O9p8k77hw4Uxs4ReVJXe/6ag4OvW++fsfwgjQUbEG2yuz2GsHAt3ZDPChIAkmKWHBwgBWctdWVqs/CSHJxOjQsME9ATwlsZOlz0qyVsSs0YxHkks077OUBEBcXrjSERdrO1tAZBY6TGmShS2BgGzCDp570uZHG3q7AhEWO4eH5W5SgpDayEnkxdBJG4r1DW0oDQjIvyWdQRCHFBIs6JpbE7WpKRi0TjuHN/ejttsWG+HC0he4opYvfudA8gXuCDCg1NvTq5ZzDlvGhUOQsaIFtq/X3RQ3b9+J1pZ6nD5zUvdJizxVYPSG8+a4vbMVO7tulWdzZDwB1ymgSLc8mWTzuRzEBCF8HRkkkn5vwmbhuH3QrC9VgZPxEF8HUMvgrv1ADESaQQmrHcNpsw2yFr/Nwv1c0aeFDWL9dLSDq9JbhnEmMBd5g1RUkUcGcg6JtWxwKbHnkg5+yhqiVnAjtjpERGX0KSoQr9kSDN299lXh2gBvJHlTq+kQ43mT0MpodB2dcpIbDFybVMxgdIaGBmITTXglSK1RJUmRHm09TkxOxej4mDKovYNafPbF57pWQBPG1EU4jxefy/u5LRYNfrc+ipV1SGA6YoqXNpXfL1RkkyfYh4nBiskc75uA9UYwlRKsRJ5gbeYCguSzkmwWQVsuQsB2hTmeDdi4NgVqAt+LAsI4zHnOzFOGXRrRJPf5+avoR+dAo6316DWpw4LggvGmS+GgHm3Fkpi8dPRwLcsU23KMprpMk+aIzcDNUGedcR/sPardpCDDrAgOdMDlkoJhjEptdOWvGTQ2aMv8YwGwnim00R4q5mhiZzAf+B5BbfZZYU1yf2JT8r5JXiK/rwF9J5es7az5ndcWgHd+8MhqABDu7Nicm/1UwWcGc1PRFGf1lpUAACAASURBVF14ABE+Q0XCxHrJhQjXVZsk5YDPh4p1kpwwO4l797/NEELWB/kABpVkhMSFNco+RAFPxZdM90jyXxRaXCQzeOlk1yBlDmDNMkx+PCT9Mp5nHlEotrm3gfsDMb07O7s17vZKYV7yjOlsYR2bAURiY2aQCyDap5OmuvZDCpfJq4g9xn4jB5ImGR09puILexAJls6iJneXwermPWGdEwxz/tDJIQ4RwW1t30W4JMVkaSYzd/ke8y935zFdec7uvKM7hi5ArzPmrjoHZIxI27qB/ezpwHppbvIeo4IryVsqjue1k8ea6zVzEYM+d+G4sE4g77mtjiexF+3dwdhJQ75oXWoZSHe0udOjXFa3AHIh1T32I362KnmjgdHR+KcPf63154IUzC18JZCEgZXmbj3N58Mg3HuGi2jek7NZnjwnZJ6X/E9YjwBh+FSk4qmYUZzdqeOF56xkmTgBBpoMWJvi0sVLsbK0FAvzC5JHZG9i3Hv6erXm7GPQFX3dPbp3AOSmdJ40jLSbtAfJPFLnzH4U0RzfrcTYSH8MdrdFqcieuxenXn0lXkzPxb3H0zG/sBE9XQPR09EjmY5ns9Mx92JWRrTI1AAow5gdnpqKzz76UNJuyHatrq/pzNpC8kTjbZkvFTB2duPb334rfve7z3T+wYBmnkxNTonRWdlYEdhEoZT5wXsyRjCEs2AHoC9riTHFKPMff/nLGBoc1Djcu3dX3TN8D33uoWEbOwMmjY+Na53SqUXxAUkt3oc9h+4qns2lSxdV7ODZ0921uLTg+AXPgtQNQkwAcIlZKHsI+6M6NVfRKm8WoHkXJnlLc7S1d4oRKdY5Cr6sFRad/jyQxw/61t/61uvx+RdXdV63tLpzFm1v9i9AHYoGTDPWImzwtY21Q/kwChQmY7gLl99hDxf5pmxARZ1uifWnPUrdJPY3YK9krtH1h3TLi9m5+OGPf6gC2dXr13WWW2oRQoy9JnZ3iMlqAr+JdabGj4l1rgJbkjvjfDVA1GYfikKTCi+A5eoWbm2NjQrx3Z46ptqQWJLvAozpugD57OMDQMTvKb7ZpfO2Q50gxCpNzcWYnp7V+qajEKbt+uZalCUJZC86umW5V2IUPwsK8tVobWY/3I23vnUx3nvvnXh0/0l89NEn8eqrr8bq8oqK+ezlRUmzWl4OeBH5I0BNsTJ5XxXerVXOtbIXv/Pu29HV26NCq3Tou7okYQLQBHkHkIvYnvkBAOWOumrMPp9RwZm1THwHAAeQBbCNpA0azYyLGLGJ1MKHU4ACZIfFWyq3yeCW62M82fPp1mxKEp3soxAlkBVZr1RicWUlhobo+hkQO539dGlpVcAbnW6sLfY7gXtRkAwRf2cdAJIDMvKsmRN0ZhDHU1zjecgPgfiRPQOD0GIhLp6ZivZiU3QWm+P8udPR0YZPxn3FHydPnYyH9x/H5sZOvPHWt2N2biHuPnqMMEtgX4t0DHsugBsd4gCm7PUwLW/evqWi5f6ePUQ4k5mTP/njn8QnH38Us7MzKq5BWOMcGhjs154LgE5eo06aAECkaNqjbjZ1xtJNoNPT5+H+LgXWLp0V7MeMm89RpICR06LIXYv5hSUBl8zxtbUNze/e/oFYWjFZhefU1dOl7kmRUJA8amnSmiQ2RB6ProDzZ8/IB+/6F5/F2tJijI0Mqzjo4i9zh6LflvKDrFffUizT4BFzGGzvVmNxeSPa5BlFccOxQfbdyQRfziURjJhz6kQgL7A/ivIQzL6Lxbhw7ryKzZhyMy9GRkd0RuNvw7mwvLqu4hzFOoonSAWiWuCCnP2ZxsbGdG4y32RILXk5mwvT2c36f/jgoeYw48+eQUGK/e/F3Lzm1KVLl+RDRK7HC9mowcEhSRJa+jIxlZMnpcC2I2Asc5NYYXRkxHN+eTl13rWqGEOhIhPeHL8AkDu+I47Eh4d4lf1WpDc6K+jqhdUuWauyc7Dks5FJje6gtk+A8jnWc44/c/HiiJ59BlQLKnybTEQRiPcHe6DLkf0cfz0IdBfPn1OsSxGfz0b2ifHQ/eztxdmzZ+Px48fx0qWLcf/+AxW18UObmhyLe3fvxOhgZ/z4R+/E3Wu/jWJLPc6/dD5+9/Enii0vXXktHt+8rZxmYmpKhVm64UZHx9UV/ujx4+gb6I+pM6fiH/7HL2Lq5Kk4fvJM3Lv3ONbWtqKEBGIt4tGTp7FDZz6AP+bR6uypxvvvvhEXz56J3a2NePLwQSzOz0ep1B7NFFTr9ZiZXYymZqQf92Jrcyt1LFVj8uSJ2Npl31qOPcWVdOd0KtZnH2C/UifthnNl1i9n++oaUoXNmm/MI+a/OmYUZ1Jc8nNX3Jr2esWJktd1AV3xalISkKwgZzXkMKkjFKKnsz1GBvtjB/9SeZhuSx6XF7gF0n8ba+s6F5hHxEXsn/ZiwWemqhycbimkdtvbME53bobdIiS4TYrlbSbYqWDKuR6FWF7esJ4/xQ86bzcrUVfhuxAHqbDDeLg7wcQ1EyrIt6304Hs30H70dZg6pUqn36dBlW+A/WTEfuXCgEmGqYMjfUMCXE50nWtlpZFEgvxS3p+yMSeJzmXy+3mN546FI9dz5Nq8F1j6yHiLeUb5/8W4y20Uus5EkkzvmwshXy7uuCvCTSKNezg6Zl/FOxqj4t/lJVm4Q/nnQord8Tbb1x6jszZ1TPN34lDNJUlfmoDWyGvTOGe5SxUb8o80PEF9P94fj167sIbky8czo+DJHuJOZWOZyo/J+ZJ3LWdm9jJRDg1ZMZGBMuGHeIo9C7lHziN3+dqLkMtjbUnusgQB2fjrqZNTeiSsI2E73xQqvrQev/nHH8AIXOwflMYzL7EdZQJWFhsdViCJE8EiAYva9zo7orO7M+7fuWeQPApxbPSYAg8OKoIiknIVg8VaLWuREVzCLKEAwiJn0QIEcbBrM4ABm9hsAoFSWzrsJlfXzQBhkcIO6e3p0wHKZlHZ2IixsREl1ix8knq6N3iJjbJrgInN5LANDlPBHQdh/J6ZMshC2DS5AY4BHDlgEIs2MWqyubJkoACCSpan4b4JHmFCkuxxrTBM0FVdXFpR4i72SK2mcRdwXY84c/aMwIObt25HZ0ermKKqX8vzwwxnywLUBRTAuCIopPjDQY42HvetVn+BQgQNGJ5Z01nM8MTCkwyUQCOCjxxoOEG3riGAl4E2AoZsLksQIskdAEdMFQVK+uBhXAHoSAgEGMqUvcvgTTKqpkBB8gLAhTmmujASu8wmVdaD5BkzJ3geYh+nw42xUsKQj3dkdVpaJKMC4KRCV70uNgisK0BbWEsCZQuYj5PMHajIBiOLZIB5QpIAACQNf0ll1eLEieNquxVbnYOHQGkV89ZRMUIAvlrLxVjfqgj0hD2FGS3dRAZMDzQPkCOT0XTWdUypnYDtfLjnrx069n39xqI2cIBiDjOxhWDIpKKA6h7pMM0BUno2h8ztxABnHAn0KBjA5iX40loU88WdCczFXKjIMkAEWCSAHMjW9g91ISD5IomWxHiRQS1+DznJkLyELLXdSkrSC8CjYhPFKWvc8h6LaDyyd6jrCQaPGdwKtmBat7sAQTu6Em408ZPxJxrKJChoLktSQ622re5yEGiSNSjdYcI8Y19jj2L/yp0LfI9/k5SSYMk0NZnKAgITxOt51ugWSsZdBOWpkNnTg1fOpooPYkQgHyBj1bRWxJBnn+p195n0XGHvUOjyGiC4yfsXUk0AiCRXFB9yG6o7XBxUMc9Ym2ZYu81ecisqJNG5Zv8S7osXhsO71T0Bvbwo8K6trCkJ1/NP7BmvbTNN+HwSYVhYgMMq8qh7jA4B/w4BFHOzr7dXRaJXX72cfHAs60cAzLgtS7bBBUf5WtCmvwPIvBGdHZ0KwAD16NZTVx5gJF1RlS137lEsTeuTvdn+B412XJ4rYyZz4YJ1R5WAtyS5HTF0IjY2Kon9Zdm13C3BfZMQAToxlzOjzL40yeeoGZZtMolT4Q4zbSTkqkrQ8jPNQS5sQwMmVRVZOY9U5EueD1k+JxeOHVy7g8b7oTtBWooAhC5c5iJkw/iNMaVAQqDM3C/r2akturIVHd3tao0+PjUVYxPjsV3Z0blUqezE3jb+GWaNnjh7Lv77X/6FgEieD8m/WEkpEHfBzJE932ODBXTT8z2SWGStVuY/zPG8D/K8HHO4y5BzV/MwFfiYxyIeADZJW/Yg2kou6GA6imQcgDzGlRTMiRe0pxVbo6+/34ar1f1YnF+IU6dPa97DtBaD8uHDuHLlsoAIinrMxxezMzE1MRbri/MxNtwbp6dGo721EAuLL6KjpydmFpej2NkbNIjUay1x8dLl6Ee6Y39PEh+WtCnoHOFa2aMA3ixxUInr16+rEF9Tokv3DevGviFrq2tx/tw5+UyxJqQpXi7rGocG+wUc29DSslvSJxfYbu8b5gugHuCB5DSqe5JM4rwjGb93/75AXu4duUNkD1lPnFtilO3vW2f32DERQhhvCht4cIjJe/KEpNd43BQzZmaeS2KKuc8aw5CU7wOG8kPsaZKwbHbxAnCUa5qbfyHwubmVPQJfBZMqDiAw0I26X42yuqFctHzj9dfiF7/4RQwODes9AfaRPkLe8tSZs5JxRNebQicFlALAbFCgo9PKCSOyFaw75rEkrJ4+FcAtw2q6tnboTDHDk3VLjGMZzw5dh7yN9vfjwb378ZP/+BMXKq5eOzzbMsNarLrkoYDMIOv7xOS4QFbOKultH9h/y95rZraKEEJhcGBA88BLCi3umsB7unm2dnbVYcF4W0rFXZCAfsQakkStrEdfX2d0dtAdVZHc1fom5JyafBkYa0zZ8S8ohFmIcglIhRoRTehowceCBt86XTKlePNbr8XlN74dv/jLvxZZ58qVK4ph2d92tirR19cTezvbklbBi4N9H4IT5+7yIv4adPK2aEyfPHsiz4t3Png/agCINYolbQKvZ6fn1CFJzIA3BFJ6JaQckfhoLcrYGpIJ76X8IRWt5VnXRKcVZ/am4i78uCyLZkIHk2IbzyPkBDcrscvc34DF3CJgizYcun8purGOO3uRKS2LVMP7MQeIDfALooivLpwmZKW8fysGS0bM6ozEm2hrS7JZ165di8fP6EyH3XsgxjOzFDkvDHZ1ccz3g4i25oN4+/UrsbG6GBOjw3H+zAmtg6ePHsaJs2fiN//0YaysVuI733s3dqrVuPfoaWxs7cTOXi2GVVDblARKX2//IVOTLgZ87ujcZr4zXyCiwRyn4xR/qPv370alsiE/myJ7bMoJyPWYk3REs4bwFpudnVUBlPVBXsVcr+7vCODkPSTVSR50AAlrO/r6+wS4Q/4i3xLgxnkmqUFylYin0881B2r1ggzG1f2ucTWDnjwKPyrLG+0LnGS9DfQPxB//+IPo7+2OT3/zYSzMzkraRdJVdOC1NItF3VEmBve6osBZaC3F4sp6dPT2yYR4bmExWkvt1rsnD1BnuOePvfMU2R1Kp6iT7JB80aR1Qbc1nX68ZqanFSMjZQWABgB+4+bNqGwjp+M99NmzaZ3B7PXkaJwdzFWK3Hzu9PPnKvYA0XHmsV9PTk3pTHzy9Knj3N1dxbnaBxQv+iy4cOGi1iD7O4F0/0C/SGp3792331wC2VQgOCohS25xmM/VtZ/L008dWRSmSjGF9NOjRylHM2nF571zR84z7g+PIGIvOk9yjGovOGvIc838Xi7kEVNyLTlv17OigzR1aQrkU2xhUh3fcw7lbk5yIoDogeFh7YeKtfl61GN9dVVnwmuvvKQ9987duxrr8+fPa9zwHmSfOXvujGIK5EivXbse8/OLceLEZJyYmoj79+5FX08x/sOPvhv3bn4epdaIi5cuxJ1btzTGZ86ej/u37sRBtRYnTh5X1wsx7OTkCZ2hT56yJ7bE+UsX4qPf/CaGRkbj+Olz8fjBMxnVF0vs703x28++iKZiMSq7dJwgodgWq6tbcer4YHz37Tfj1NkzUdjejIf3H8Ts7FysbW7FdhX2+JaMtPfxw6ogq1zW83/5yssxv7wU08+no6XV5w1dT8RHjCNnlhQadncllZS7oyXnBFO9uzvlIc7HJfsn8p3xCMVudPGm7mOKQlJoYB/e2tI92KvQ+QF/p8gHwQVyQm8XOAaqGPs6JykcM0d2dg9iaBDvCszTqzo/s6eo5i2kKOnxN+ssWFtbdyETTAACFt1yhWbJzbWWrdrBOmXfhixLnEO3IXn8YaGC+CwRZYmr7E2Bj2gqI6Qu+y/Ft/+LQkUDsDdIL6WIlGEdLRvkgoXi+a8pVCg5TwRT40Ksu0aB5GghxH0PztuOAuyZhJVzmXQhaX3mfwkOT/dsPDBjDAb1GoWKoypSvk+v2UzW9TtmfMgSdiI0f6lDJX/u1/+Z8wnhSyKTEmO7s1LdbEkdhHVMnK0cVB1UVe1dxgDAI1zw0GcngqvGUAUAJmdDYSQX2XJspJzlKz4T/FsEleyboTPTxFphGS2txk8422VW79w553b5uu27Q87g+cb+NDhI3E6u5OI5sT1znOvlfdTBlHAqniVxFzdIUZ4Y55tCxb8+p7757r/DEUD6aWEBkzjrRsK64+Ai8IQJAiDNIYGskILc7i7pnT588CCZ6B7E5Nj4oRkxYDgHpJj9yCCJIelNBGCYgFkt7qmFnSHz5m12PMk716BFL3klsywtq1KMsfExFRYATwApBWigC9/TLQDROuoExTu6djalyuaWEiWSZRY5nwEgxp8kPhxWBhRTS51aIBPwl6qxYoRID9RGS+qsSEkTXSRmuraIAUoxplRqiZLaxQkcYFYfxKPHTwUWAIK/mF84NPHkd9GThWGzWVmXzty2WrlgB9FVAfhOC3tTrKwuaxPr7GrX/QGScK0Ac1w/AYaAWwXXSMLsu33+iP5k3ngNEiV/BElWOQnkPdi8OfgJ8Pw8cjXcwFk2Rs2Hj8YOwDqxrK2VvqNkggIAz5DCyuz8vLtuEhNfwJcYfWbrC4xJ0ieMt1vuk96+GMG0Z5olDptQlWslPQ6YeE6SUtjdcbs5BpWbG2LtMya081K8AAylLdsgNkblgLzIYJmJhXa1Zch81CqA2tlVm39ne4cSbOSeltZXLbsFsF0qSUdXgVQyISbAzhr+gAU2doRBf4TFlGDeXNE/DBm+8oXMUtY8VJnfAYsCkhzppPfVIUvykDxepJWcgHrGm+eh4gQsqHJZ8wM9z6zV6M4L2P1uG2YuOFF0uyT3ypRSi3wKAMT80tpwUpfrLlnzsY4es4ogaf0EMkwtybjVMhg8W2QDGCNLTLil1ACx9wQzdmxSbRa8u6xcSLSsWAbMGQcVWZNGp5jhOYhLhSKkDegogamsFllJQvE+SZoHAKd+oCIs12Xz0BSGZYJKKhawXpHHY2xJ1Mvl5N+SJNkUrKq45KIPxSxr+RvwUAAmaTMHi2ovhTWLee2Opa5yAJpBX2ll0p2UClg8X4Aj+wi4WyAXavhsEkgKwBQJs6kwax9GnuSPkq9NDohzYJ3N2jkPSDRz94SZuHR3eR3m1uS2UjHeeP0VJeKwo2BvMXa58AObMsvykaisrK3E9MysOuRU/C23KXmSATQBMIXLWk0MZJuHU6hzpw1zw6aMliAD/Gffk3F9NTMlI/brsCIdGPLenFcuzJoB5nlmsFPMrxaX2NR6m4qn2VrTnTNOvvN6kRyJG69sxJbkWmC/cE0qKlEMx3BQ8xlQxt0ijAF7j6XNuCfLe/l+DrQ2DCK580I+T+i7pjVucJa1AcOcorzBU8ZJxtqSVLJ0GpIjJ06eiOquTQmRf9rZomtknwsXUPf3//MfXbgRuMH4e+0cPf9yIdedHQZV/LM52XFLvP2hPB9ddDFDT/eWwBJ9DYICyWQ687NmP2cGngeAUFOTkzEz/VxylMenJgV2AOpOHZ8U8YA4YGRkVEVQSAywydkzmXesDc5nzOmZj8y/XFgv8az3d2O4pzOOjw1FbWcj1laW49vfeye2a3UVK5qK7YiEWFe8vVMFA62L1HXCmLMOYIJTDJRETqEpPv/888QCxHjRzwnN8fkXc5oXdBhxdiLfonlYLMbp06ejo70Uu9ubOoMp8qsQzryWRi4J/W50dfcKVACwJ0ljPv7ql7+KickJzRHiO8AjYiYMXSnusA/CpKY4AbjAeGiMU0HX8h02f52amhIjlHEjNrl581YMDQ8eJoHIhwG048MAMMccAMSFIMBaYA9j/3S3HR0jmMznbriCnuvE2Fi0CoDcj62N9Si2NsV7770bn3zyiSRkiB3mF5dUhGLfqmztyP/MMZHJH6C68v0S4OJ5yMveW51ig2PATvxinzNLi1niIflhpZiDeWZ5TxdTAXZ+8MEH8eTp47j6xbXEiDfzV/N7rxodbSWv0xokjU4VXdjLAPYBZ6y73RYLiysCrhkngH1AGxtAAtJCoAGkqinmpjBDv4LGD2JI6s7VGpMuf6t0vGGiXrpwGj6oQJjOrt64c/eRyBOtxLKwc4N7LcXeDkQgNNDN1DRTkc4Ig+bNBXwv6tHRTjGlGO+/90E0lcvxy7/9hYyWLbdgSRX2YQFNeztikh8bHdG1Q8JBCkTSgJJiocDcIrD0yquX4/SlCypWUIyorG3GrZv35FPRWizJhBagTZI2aKJLIiligE4aMWsr0hMhgWe/hg3LmcVcZ1wA5dhXLl++EteuXY0b1+/FSy9fUHGNQkWZAjHdwfsHYsJDdBno7dNeivkqoGeHimuWo+GlLq8dd9VJdhLPFHXZ7elcZt1zv3yPayJG5MxDh33uxYt4+nRaAL0IEvvo8tOHcBAt5WLUkI3jz7396G1rjePjI9F8UI0T48fi5MRo7O/uSEbryfR0rG5sxZvf/k6srG/EtVt3An114NixiROKNyjojAyPKLY9dmw0KhhlLy0prqPAQpyIlC8x35pY02aub29XRCyiqJg7Bom/mJ8Qe8g12JfHRkfF1id+zlKYFM4oQhAbs3dRBOrp6nJHYvIPoluXa4D8sbIGqc25GX9SPJidnY8X7DfKI8zkpuNHZ4+60u3RxXOQXGdPj7p4Bvp6ohs/H2LRnUpU8Nja2Yq21pZoI34EOE3+XxC6FhaXo6u3T/J70dwq+acvrt+MW/cexdDIsPa6WzdvaZ+FeMBn5a5yxQwAW7UDkTygpogcJYJfPc6fPad9GIP2xcV5rQOICYzD1IkT6pCiS5uxR6pwsJ/u7nXvXfhh7QJsT2pNP5ueNrCW5DzYw5Dq4ppg/Xvf8nmqXE9xof+kMMIaIO9kzOka5cx/9OixpbvSGZ4BWM7EDClmEJHnduwYBMRN5U98nbE/MTUpr4ujJIoMmPLZzDG6kPAQUS7Var8M8gRJLuLL09WpWCcXkzm/OUNzd7jGOZEwVLBK+ZHIKSkGOVqoUJe/ukvrMTw85H0/SYZRAKdohDH8Sy9fEuGMQgtxAuPEPKLDgmtk7CnEXbn8cty4cUPnGV0XkxPj8eDB7RgeoKPi3Zi+fzM215fi0uWL8dnHv1UR88Tpc3Hn2nWB43RLPHlwVzH+0OCI7o39kPGeOD4h1QQ6iMZPn4+n957G8gqF9t7Y3t2PT3/3OUmvChW7ibTEcx3q64rB/t64eO5UnKYTpNQq4tzc/EI8ejYds/PLEQW6v2vyzCCmY98cHBmKnequItitbXuqkQ/kYgLPQziIiKE+ZziHsvQz45/B1OwLyHNSDIesVCKXsO8RT4mcqYJn0V0SFXAJJNga+SDPV0WLVLjobMNs212m7CmSBq5HzM3NR7lkpQPPFXAjx9wUKdR5T15XKMTaWiW6Oj23WUvqqkhxZ1t3u+6b/Zs3LpfaVLSAMkeHhgoVFM4AhkmrdRQai7CKgPNVd/6an8OfWU425+U5b280KORczSiCcrzUhZCJXblYkUmLjUIFbqLGHjiW9WwOO5QtA3Q0D/xqoUJ52FcKFV7bX99R0egaaCiZALB4iI90UchfKu0WR4qQGar4aqEiX5cB+oyLeJ/ifXMB4MvXb6wp5z98mkjAyReC/VNdtPKas7y5uuSRR97dU47AnGUPdw5Ws/RlIvXoGeTiA5+TqmiZAJgLFX5WuRjbkGvK180zUBe9sEHjgeo4T3gbewrrTAV5+WiZDG38wXLgWQ4rFzHozH7pwjnlsVILaG4xWaaKT5K71uhOUg4IZlZDHm7NReqDejx79vSbQkVeiN/8+YczAhf6BsTGZ1NgIyZZZtETFMI49CFhPTwWKAl5a6kYCy/mU2FhJ8ZH3a7KpsPCJZGQkbVAlhYx3QjmARasPe3kiE3GG7MPosys5iTgI21e6jZiDK4ICNh8CDgb1U719MXm5rp1D2VkA9PfjGkbPbuVFhaRWonVLWBpnkQdVgCINiHANQe3WOvIgaAVKXANs0VLi/R096p4Q9GBA41WSslUqDIKq3EzdhPLDOYeLBmu5fqNOzLzOn3mdNy7/0AAPu+NpBbsR4KDpiY2dOuNwioj4QDrIFDV5txWjr6+brHj0A+FSUjgQfVYP4M+rAA7mx/KGJxNLQFcPA+zXwzQ2XTbjGM2P0ubGAiW5E567g5Mfbx6o7aRm8n7/prlE2CwMY7lZJBJ8cIyYJ3d3eoAURCQ2G5iRgiss3STAhIKF0e0mPmQw7ZBkhtazl010nwrtVgjXya9yVcAJjmgDcESAC5VeApcBKY8NxiksDCyJAmFOcAMBf60q2NymvwGtC6amqO7HV3NkhgpTa0tYv8j/YSZMXOMZwzbk7Z6d38w7oA0zOcEaiRT8Ky96Aq/ORD5wMy7S04aPMSplTbJPHH70l5OwL/glBQIZYCS9+N5qgtImvIOOngWzHUbkWOM7QIA2uEyWU6HqdZjYs2I9a42RUvB6Gw/Egghq2ZTNF+9/UwackEaV+4wyXYxYIUkcURXAkk9hzKAJs+XNaiwikKJABrfAwEt65wEb2fHAIYLZ+6a8gx10l4udgAAIABJREFUgMW9sR4AtTAczQd97mISB6TJkg3SjZYJnAsVaGtbe9I+Nazx3CZNUs7vcd2MpecqfSL2KSAo4gVDkWJW7kARqEt7aFpjjC+FU+aH9LFTa7F0T5PHB/Ob++XnkJhzrOlg0vPG18d+S4KAYaPMURl8q/J4zabomX2X9yPRplNBHW81+2PQQcea4VnmbgdJVKTfZV+isMTzJ/EUKJ2kVwzAtykgk774diVOTo0J2EBO7ezZ0wJGkeLgOfL+BgddrOJzHj99IjkXgJS1tU3JGWjepvuVd0qas+zNJGvM1yz9hIk1P0+RCeBNoJ6S3ro6uGB/R0sKjrV+vNeR0LWXKY7AxHZnF193gMgZkOTaEosmbXnak9SBJumlVJCqsaciUZQYjqm4wtzUnriPtCCglyVB1IlEYpTYUbngzZ+7u6xZwBCbzjHnxJgRcx+Q3XrZ1rHOerSsaRsa856MAcxXxptiicybZVLp1Ag2t/cZZBncGQOQRtKGjFIuTLqQXzuUVOQsMoDjlmxrXiOvZ4k9FeJSl8SXz5lUeBEI43WqGCD7JqnQjSygz4yckAlMqdWiv79Hkkh0Bsh/ZGBQc51z5djYMUuf7VIs7FMyyvfka5SYxPwOhQykFpmLnJGcFei2V5DGaa5HT7kYYwM90ddRjvm5mRg+Nhob1WpUqvWYPHVW0jyFerMkamBIcxesT+at5HrwnEArmQL2GsxFs/6Qk7hx61aKa+oxOTERq2srSm6Ibb77ne9oL/vdb3+r/ei7330npp8BNlf03pxHxBkUUHcTgAqozTqmY+LOnXu6jlOnTsfVq1e1/zGuMC8pPLhL0qxXJ33u2GHv4fcAJYldKMaeOnlSck88R7o7Hz58pPdTV8KzJ2JKb1eIPzrs74Uejkl19nrK5056tujIW24TAMN+GirM0l9XsEdAVzvdfYXYrsAE3o83Xn817t69J9kKCip4TXCdeHtwzlCc8lmwKQkH3o8CSC6GUagB3IOty73CLMfrhv0LwFQmu5kMkWTHmOPMF3uvuMDJMyQ2+v73vx9PnjySGavXowvLOUmUXB37RpEu5NboKJek5e+x9nURGywur4mJzrrJxqYGRWF3Mmfr8WR6xmxykuzWop49cQb7BePMPejvGI0WAMlb49LFs05wWyhqDcatW/e1FyH5gbwNutsL84vyBVleXYnO7g6ds8TmEIjoj44anZZ1dYK89ealuHHtTlw4fyKuvPq6ZG3+5z/8Mr7zzndcnK2iSY80LJrgZstyCvI1GN3Zq4NnlMkFdM3hd/LKG6/H8ZMnVFCv1Zvj899dj20MulWgsM756DGkDFfS+d8cgwP91sgmNpeMpMEMirqMB/sP319aXhRIy/PiOfz1X/1tdHR3xp/8yf8ej589i09/95mkcJhE5dZSzE7PSNsczyMKFBtbm/pM8h/+HB0d1f3S3ffixbziWtjWxJDcW5Y/4ZwErOcziSEBOVkfLAqKFfPzC/FYzGoKPS5UBAUj9rZ97/N1pBk72uLM8fFoa4oY6umIsycn4qC6Hfv1eiysrMfY+GTMLS3F7XsPYnWjEptb1Th9/pwKNqx11of2QNZzZUt7436tHmPHRmN1dV0muMw95gpzDBmyyrb9A2FwK1bv6pR0antbh8aG/Z2z1V9z/Dw2Nh6bW8hrYHzdkDWE0GEDZuT9kNFFriXvCc0qMJKflDCxR8a3p1fSboCGOouSvr5ZpJwvnNk+KzkX+CwKJdXqrnTva/JJq8v8e2VxQRJ++1t0R7tjX11N6/ZNpAh2IKCzIMN0OlHOXbgUtx48it988klMHT8er736irqm7t27r3sgT1MxL3lFQMgy0cpWhvLmOjiIs6dO63cAy9kzkT/iP3LW7u6eaO/sUiGXQgPvS67J79FFkHNfpJ+YR89nZlQo48XeytymA4NzDP8EpLByp7ONpW1QS0p75sxZ7d2QSSiCcjYwdk+fPUuefxylDtS5FxVApaeeALTEtB8bHxdYry5b4ru2NvnQ0A2icz6RlnI8RBzCelA34dKSci3FAiKWIYfpPE+xCjmIyHR+UaRhj2Q/pTjJ+cm5lAlxjgGdUMjTMcW9znHMeueO6FLO3kqW+mlRngg+8Mrll0VOmZ55LjyAjgr2X7oduTbOvJmZmbh44XzcvnNHBWN8QSYnx+Pa1S/i+MRg/OQ//zj2ludidXE2BkcH49N//k30DwzEyXMX4v71W8oJ6PxaXV3SHnRs6kSsvFhQ919Pb3dMnpiK6zduRKncGcfPXYxnjyBcrEex3BkblZ2YfbEgj5c6XWJFm1PXD5Coa4m2YnO0F5tjGLLG8SmRAOvFYty/ey++uH4rogn8wax3ddCBgdCB1FzQvSyvrKvgz3zmGrkmd/E67ycPYO5ZMtTFAM4lcmgDyyaTqrOa4q1iXEsvEo/0dnWpUEH+AzHQHn2cLztaA6x5S7o6VKB4IZyH/BxiitZ1h0inyteQSdzadldzOosVLyLRDc7A9VBgaW5WNxndhBQmeRFr86y3ICy2mbAoWSXINJyzyG+3lt1Rsbcfa0g/pe4JdVVkE2nFp6m7QiSkRkcAc7EB/ueZ3FAXynlTzqdzkcJFNCgFjpca2gpZIsmdF0fLA5ysxkq8J5hUasKP3uZL8k1JEjutiXxlTh2PMBrT2nNRIMsbpdzS2XcDdzlcqY1ChaSc0+fmYml+r1wQcZHDY6ic4whmIFwiEUTy+xy9j0wM5r3Ze/iTvR/8hd8T2YRzhMKWvC4OlLuQpxNTQ5jWM5fsWGYWprFJeQd7+levKT9XX0sDVxHR7LDQk8fJ2E0uQogQlrAaF/Hsocm6kIxY8ltRISmRtlin5DdcNz975swJmdNLEWFvT4VfcD5UKFgrrBMIUJJEbCqIdL20gjdlKTaRO/9G+inN7G/++IMZgXPdfQK52QByIEClEgALppyNEnvFDCLZO4ZJWHUvXszOmmXR3BI96Ogmk1oYb0tLiwIcWaiwlTm4OLSR+xBgniqYqoiK7Zu8IZImvnwKqEAiVbJeiSuvXNLByX/IFkw/e27T0wTMkkj29HZZHgHtayQ4EmND3QH1ggodgJvXr98QwAPTWQDCIWO0OTFzvWGT/HN9tIyj3UoAyGZC4kuAADORJA8AYH7+hfSyAcOmpiYV+FQ2d6K93BrtnZ1x8uQpBfYw/9h8YII9fvRE90dCwEFMoIkMy8rKksCL8+fPiN165zbBcnP09PQloKBHbcGtrdYDJZgHfOFQZ6MmyGh0P7iA7kTRm7wYeElOSZt06gTJIJOBMwN4R6vvrghzOPp0NbjkjTwHkQTKBnDNggD4INCFAS3jvTY0fNvj6fQzbbyASDnAdEu/pTNsouZiiM2NLEHFzwsghQUHK462SxjuO3ti7JFAcV0E1pbwsi46Ujy0LwNO8HuPHj5UQGTz0z39HvcAECC2/EE9+gb6NJfoEIBpBuuuur0rphjfJwAk+FvZXHcrrNqa99VRkQsGgNsYbDuwsHSZAN12S6DkToSvK1QcLVLkRICv5SKSCje5HVQP3MW+/LLJlgtIh8UnGCHpmTP+2TeEA13SRk2e41yXAVODhSr+pPeh64BnRlu9ryuxwQFUGK+adeRdLPHV5G4eAl+CLTFy+Lqwdu7CRVCSOIBqAeDq8MAXxF1BSB4J/Gr2tSDZY2MsS+4wLzwXHfzy/HluNqEmKDWYag8DJKOKlgtL7ZmMF+skm2llFjnXlccVo2nNscx0J8AApEs9sDDD+FlAxaXVFfufwORQIcDFURVBxFB3IYUCaDbUyoxQrklJBuzgg3oM9mM2vW45rbQ2lFxS2EjvT5GJ6yep4HrQ+JYBZdJez8Eq+zHMUti6BH82fnenGfu7isMwn5NOcJ5PXLs6PVIycygRlaQxsnlpNkbEl+H9d96Kra0NJbU//elP46OPPlSxgqSd+6AjDtCHseFJwgJEI5zEH5A8fz8zmyzlYdYs64B1xHwiyadzAoYoLN+unk6ZiTKXkKtgnybpVxCNZBJSXKkoivEl4yi2PbIEdHGowONuB9hgdK+hz01nSO4m0NxP3hAqFiSmL4CQioap04J9g/kCOEyhVM+2uSnKxTafPS0wZoqS2aFIpLnRVNA8yz4Yma1DgYwkkyIIgDXPVPJ5u7v6O0khoBrzZm5uIcol5BXdraZaMAageErQtVSke5G5KOUTMdj36DwpksQhoVRUIpg7zSg6sEakRX7IanRQngsdLryY6MA1A4ASB+SOKhfQLV/I888FPUnmaJ42CkQC0hK7391jB9GJ9E/9QAAgngG8F2aXL+Zf6DqHR0cUY3B9gCTIp8GchKXHONMJ+ujRQ4Hec7NzloJE7qu5OZYWF2ISE1qKmvWdeP+tN+JgezNezM3orHr9vffi3uMnsb69G+WOTrH9hodHY2NjR0Ab5/vA4KDiCzohtE+nIid7K0VL5DC+uPaFANzhoRHdn3xT0NLfhP0aceL4Cd3Xnbt31NV6+/at6O3rjvPnzups597EymauirUNe9fa8sQs7EdLy2sCRRlngBgACSVLFAhlZN+lLhTmHGAUsRSSF8glshcQD3IPdNRyH8RcFIY4z2DkEu+wV3OdgNLZx4f4QIVP9ihit82Nw5hDMl6FFjEWmQ8wLZmvmS/L0TXU3yfwm3VWWV+NH//oh/Hpp5/q3H74+HmcOD6uPWppeSVevnxFzG6KtxA9APSZ2/JyqLGn7MUPfviDeP+9dwVKAY7/8pe/FIBGXMdcK5ctxZa7YUS8SOedOm3FpjYYzx702muvxZPHFCquH3YZ8SwssWY5CcDciWMj6lhCsx9/BoBh4iB7vezL/4p92iQSktmW6OrpcZG4uh89ff2WvpP0pYyojhBV2hS7sFcRU1liGTm9XZkqUoykwxT98k8++UzgF0Dx05nZ6OnrVizM2cI4yGtJuuNlJfsbq+uS4QIQqx/sxjvfeT0WXszEowcz8R9+8kGcuXAh/vov/0pjTRFIIAsFqB2kTttU8GP/Qg4KeSGKQsRnzC/mHGcI++C9+/e0Fr/11lvaA/f2C/H5Z7eiuaVk8LOVvadZZx6dXfJsKRZVKBBhASm7XYxquZ+61glzmXlbLpbj/oN7IpScPnVaxVJizj/787+I7773dly+/Er87d/9Qt1QsJ8BwhbnFmJkaEixAu8rtny9pqIceQN/wrAmjudMx5sGU+27d+4e+p15j7d++y4EpJ3dmJoal14/XkzsZzdv3YrVNUtKirxCN8h2ReecC07N6q6o7W1Hd7k1vvfW6zH35EGcnByJl8+fFeGrgq8DoF8dLfVm+S3gu0HBgjOHeUMORpxB9/Dzubl4+eUrut4HDx7qfBO5p1Q2WF4uxebGun2VkN6pbOiaeVa9dGolib/1dXc/QoZgzjOmdFq0dbQJFDUaVVf3EHsvXgFIRE1MTLjAnvZ+nWUAmJXtKLU5LwE0b05kI0nZAaDLey+D6HXtlZA++H32M/YxgPhC/SBmp5/F3u527FGoWF7Svl9ZRcZyP2iSo5gBts2ttHdyHheCUwgpJsbw7Pmz8Ud//J/i3sMH8bOf/TymJid0Rly7dkOfq3yQ4ujBge6PdYofDgCp8hRikjiIC+cuKL4hz2PPZ+7wu5KF5bmt+4ygkxFWPz/z5PETqwJgohrOU9njMaWv1+1Zlkld5J68KHQASvlsdf4FKKzuyqZ6HD9+Ul10dP2w51Oo4L3pFhDRIf0OfyJdyO/nHMEkP8e8eGKwT8gLp1DQOXpsdFRnqFnHxKBZksYxE7kea5qCFmteHlM8jyTDQswpeZYkx0r8wnzkvbTngQfsWdKKs0ExMMA9nQApZlOB1tmHxoZzT34chyoHlsm0Tnxz1PeRkqvE22+/JTnIGzdvxOraVrz55quKmVmXdMvSaUgnC2ft3bvIoVVUcIJo+Lvffh4Xzo7Hj3/4dmyvLUZ7ZzHq+3sx/eSpzrGTZ87Fneu3BNAPjozEnS+uajyOn7sQOyurKoCMjA4LP7l240Z0dPbE+OkL8eju41hZ3YzmViT+qtGMEkGtLpN3QEpIPphpY6I9OtQfdH2uryxHV1ubJBlPnD0bCyur8ZvffREFpJ/23XWLAgPYxebOpvYbSUbuQmSs6ZwSAQtQF0KFgE93RwACS3pJ8mfN6kKU1AyKFkh81kPnM+cG5B7mizplKHKCGeGvRL7VzHzpMnlUPhhNGoP1yrbeA14DsYCJkJ7/nMVmijfL64pYj+thrt+5fUtzrqvdEs/IvrKHImDIvrdZ2YmeHnfP8LKBun3m2jo73BFBjigfGt8HBXHydqQG12Q8n6SfEoXGXTuZSAMYbfmx3FGRwf1DhkaalblmcLRQkQs9mWiWCxUZ+M69DhlXYbxMu2vMc363Aexn8N8+EaaspXxbuHyi7B3xqMj5evqpIz9/tFChjTwRgRu+GIe/c0T6SYdWpgYekkmtpnCYN6b9IRd0GkB/vtbcOdEoejSKFYmw9xV/CPaQQ+Id3dfJU5J9IeNDzEnkbtW5njGHhDs0xikbWyfD8MOrPjKeSbVCxN5MrFJ3sOXVmSPgCBRZ1d0hcjBxrbswiUWRTXShwp+nriAVBrMyRMNbcKAfqXgIULvqCmcflYy7Pq9ZaiDdHZ0iw1SQv1ZBDUnDgogVxPHfFCq+9CC/+ccfwghkM20OZS3PAubUnQrOOVisl+fNh4QOxhGbKpU7GZByuHV0Chgk+ePgU8sVoFaqyPPzqqqvrx/qy7GYsxwFO7+Y/rwZqAksyNSue/bMGQV61kdv0vsgCYIxHwE+ASSMGwBMNglrigKYFBXMmhnXpOCWjcbyU0mPWBI4xcPCCQEVG7yMmqTRaDkkki4CXLE8aW2GVaQE3f8mcORgh8F08eLF+Pjjj62lK8ZKq5iTBtbanZwXCpZ+WqVly9IlZ8+c1e9MTz+NUrlVEgsczBvrJGkEBAeSsII1vLe3HceODYv1KvaDWL2hYhIsBTGak1cEnyWWemIrCWxMGrBscmI1JGaaAaUGcz+3veWWvSwNxfi6ONGQL3LRIrcV8r50npBI8jwLClpnZ2YE6tgQdEtAmGUXDJ4JtFDwTMDtIkoG5nV8ApQdkWPgcBAbP2lM58CWxIi5QYKrjgHYP3hmdHcrieDZ0h7PWEgKqF4XyMmcVOW+VjssVCgYqtWiG8NLgpwWd5ns7jtxgrFRVedQq5JWujRyUULSMGr7c5cLLxIxQA0x5o+2Zqbhy1/7l/YWzW91v1iSovGydNDRQ97r2QyCrLWbx9WM/IKeEQes2Ae0xSZzVMkZJCY+95Pbg3O7pYNT5OKSbFfS7+RZKjnQvaXrS39k7wl9NiyVzARxc4DAvPX1Nc+ixGYgFjKrzvOW++nsbD8it2OzZX4JNiYMA9aITLthy4itbGZXBuoAS3ju7sJo6OxyXaxj7lseOkkOjHnB3Ovv79Oc4mcoyJDc8CwyG02SZjJu7ZaMlLxtUjElF9/yHOA+YIgyZ8Q0ToVY6e3KUNv3rCRWXV6WUVBxWDruXmuZWcNgwjLkuQgEJpinACBj0SSlkzrYGFDer7vH+rPsD0pqq/sq1DlxdTKY52Nm6Gu/T0BnluXJQbKKngRgETEyNBivX7kYz589EUMKIBJzUdimJDzsURRYPYcLAnFhhdh/hWeF/rUDTxX+YNKlYqa9HRzscTZQ1IChvFdFd95ms2K5iLHjvcgt3Jil1rSXy2SaBC3J3wn8lexg6VDGSeOWOvD42dzZxXrIc5xCh9nSPjsVnNIlgm48pp4KYmnFp7PMewDAXj6r1F2SpjvXyQtWK+dbNlvjugTcyyvJDFMKEHjD6L5gxKX2bLpJlIClWFtdXcn0j72TTiHtpRQVihTagGwKAhT4ey6mccZmzwneLBd9XSyyXA6faZnAxK4To94gQQY/cpEvd1/w2TqTk1QF60NBuBIBJ64+AyxHoU4VnVdoD8NqLchEFekngMnjk1PqkCC2mDg+JcLA3j4SAsgvFpMcEqBcs5jFSEQAGLO22fsAUNjbYb5iXL23uR4jfd0xQaF6byc219eitVyKvrFx+s9jebMSz57PRUdne/T0sn4xA6foaKlI5jRAFmAdlV+A9iwxQXzwfOZ5LC0tRHW3KsCKr5Fc8JwAAQH3KLbcuX1Ha3h8Yizu37utLgkARAAvGVgf9V2BVQVojSdEZSu6unrji6tXE0mhXexcyfsVmnSfo6MG0Og+ETCxZ1kOroU/AacAqViv/M742Fjcu3dPpAxAB9i6FAnzemd+yatGOtX2HhsYGlTMxXrmhc49RSEBusRvq2uKfzynYVo2yzcKtiQeQ/hVXDh/VgxleVlontj7Yz0x5dRhUsNckCI1nZhJUqDZYMrosREVq3PcCZCO5EqWGmWtm1lpWUPiGsAWxgNmM9eR/cdg7b/77vfi8eOHAjDzvOaMpzDAGi+1cuY0q6CmMx5CSOoOZl3JWJGYUUUsYrdd+b1xbwDnRYqs3b2xuVUREAyobTkrS3wxH9zJUFWsRwEFM2E2hZ2dzXjt9cs6/7if1pZS3HvwJD76ze8kpQhQjPTixuaWpGDYXznniIW0VxaaVTBBfisO9uJgbzumpobj3Xfejk9/84lMjz/4wQfRNzAQP//F/4j+gcFkIm1fGWT+SJx5joz98akJrT0KeNKar3qfQQKLe2COUxh7/Xvfi8XnL+LadYzWLTValawj0K9jGliSdBxL1o/CCmzhFsgKG4eylCqQ7+9L+od76+nqkcb+3//9r+K//tf/K549n46/+tnfxQ9//IEk2ZaXVqKt3BGVtY1YX1lV8Uckko72GBwe0h4CmEpszpxDygY5N56dCxKhDr0M5Bok2dPcoWOtvVTymmwqyNvijTfeiE8++VRdD0iZSa4Po2RA/ibWDtJeyTRUrOGdGFE3xVjU9ypx+dI5dX5SuMFLCpP1clenzLRlAst+ANlmYzM+/Ogj/claRWaNuOj119+Ij5FRQ1Yr+bFRtCBvUkwCQ1mSosTDlnHk/HWutB9/9KM/0vpm7n36yac6LyTxmIqmuZtVvnTVfcVKFNtPnD6tvAAAVsbGdUuw8DN0zTD3DqJJXQV5ntPpRlHexcxtnaMUvIi9stQiOQ9rgBgMkJNiAVsNkmpbFZimTkeYzrUqRcmiOgs5WzBwh3iO8TDXReENH6M33nhdhf+/+Zuf6fzMxRz2DxUV1eGET1hJHdfWPgd4MqQ4NDigOcH5AnmOQhrjB1MWiV6eO3M/SzFB1GGPlN8Xs6F2oKIwL86qnW2T8fK6p0DPHMVnx4Qzg1c5lyB94/xn75qbe6HYhpgCU2/ioLk5FypcHHL3egYOOc/5ej7bmQyQ7jD7tgyl9166cjgLBLrlbrk0BuzldGbxczwznhXkQABryY4lrXb2MvlIJN80xlAF+ES0sqya5VS4vxyHimUuuZMDAdUQWngGFGLBL9j3FNvwfhSs9/clvSdPta1KvPzyJcnkcf1cAx0VfAbdgjCVOeeQtbpy5WX9DLk1uTvm5198cSMuXzoer18+G88f34mJU5PR3kSHeEE5es/oaFz98GMR2iZPnIg7169Fd2e3SInMjidPnsbAQK/O89t37kVXT18MT5yKO7e4lnq0lNpjZXUjKts7USMGammNpZU1k3jqNRWPy61N0SdJwWbJwVFwGBkfj51aPR4+m9Z70InMuSIJbPaW5iYVO+hSB8xvaSkqf8rYQ/Z1FIif8kGK/8QxxOrE2tL+R04p5SMi3EFQknqFlRgYR84+YlXIPVllqFiyb6nIKyK8NQdelcRfzmCs1sFew5qXZJPOIDzJiopPuA5J/xzUZSIOk1wFMAr/BMRNhdjY2I7uns6oIXMlElRRZ68IXSK9mCBTQmouydGV2zpU5NiCfV/Z1rNUj49SkoY/Rb6/RteBY/38+iqp0LlAurdE5nOhInc926cxuSN4fuf/xLj3Z+dChWCxJN2cEg29vzs1Uhvr4dU0Ppvryt0gxvDypzSuzdfqMyA3HVjq1nJ2itMPb5S/WGrZr8PvpMLGl++Zn5PvVXpj4UzJR0f4RVLryATMBnbha8rjKhlmESFdGFahCjJSV3fq8GtTPIpiizBKPCyTQTsEjFzcSQ/FBNGUazSuLXeKNAbS+IUzVJleJ4KuCWqJYCRCHZ0djm80Mqnwm5oDdc0m+jYwDOc0lis3YamoeIHCaE9PR9y+fSf6+nuFXUAUJxbR3ix1DLC1zuhoY/3tu+M3DoTZLi0uflOoOLIWvvnrH8gI0FGB/i6HT9YoRGOTxU4QZSkNG3DJgwHNdRlGbynJ4QAY7HdLNmAorDtAT206km+y8SkBP9JLvIfW8iEj362DktnY4xqQ7LZkDgvv0qVL8Xxm2qAT7BSBNq0CBNvK7Q5cVJhoBFpqM01SPFwLTXRKiI+AwzDPAIvYANl4SEglNUFw3m62OYc0GwkGc5vbtNHaTDpr9hNMSm90YVFABeAEXRWYcymooqugH2Mct9hzUPH7MEBIcGDZyRNib1fmlXQgVPd2xG7KVflHj56p0EKS7vuqqXtEB1Xy42D8SMKl5QsBL4F9ApVq+9Y+T+bHZtgbtMs6eT4gfOhktoBb3hrHkTZrsazRsHeQ+3uv1NrHRRDMswETuDKukj2p1WJ1fV0JlEHC7DMAoGi9ZQ4ngWJib9vM2vPFcmFigAMws/kjt5XkidDPVqscQbAkiMzSlVQGZp2dHfoeQDgdMQBCvORnsmVzPH12qobzTDq6YNi7WEUSUUOSRJq5EVs7O7G9txOVne1oSl0ozDVY04lkcGjInoMLtf1JOinpuJMUZo+WBNy5EyG1ZUsDzI+mEZSY4ZGleRrhQuampqeiFmsXKXi3w2QmBQdmNqcghaBBAUWjjVTm5onBb2kmM2hzQsG4krQ5cfM6AqwS60lt3r8fQKGJjfSTAN/UUdGYQwUltwqFEhgKc7yl4IRWn2PIAAAgAElEQVReEi6JoeB5ShCKVFNmYhuQZ+4hccGLOUfClOWbGhr7lmsSuLC3p+KMO8osYcB6ADTInQ+8F//GeBKDRCSnWENOUg2sZ71JxpwuKbGfYZwlCTOYp5l9m2Xv8ErILH4B4UmaKwPz/Duz03W/6Znl5+ZA1GvIRVZ0jvd0DwQ0WVPVHRKWVCPcQsOTeY3JIkkI12q9bSfj7Au0ucLCysGjix/4wpilrcJ2KjAr+Ew+CIwp74fO72BfZ2xuWPue4pHWYbf3LvmYREGAPJqxsP0A6EioOAdIZJSIqMvD+tZKPjkbWN8UMyg+pc4vwCFLOBXlQaF9uupx4aWuG5yQk3SVZKEAMlRMdACsomUq7Jm1B7gIuOF9VGGoJOp8Zpg5Y0M2JJQciONpaGN5kj2eex5TDk72OZYG+qKwpy1jkH4v/V3riOJYCubzvpGN7iVzwrmcEnft4+na3JFGcdWBs+a81rYLvbx3Lvx5L6cobMk+wKnsAwLIxDOgcKazWuxEy81AFjgqCcVabkh52TcoAwo5ERBYlRhIBkqcZLHvZtm7nCzzftnvJO9bYg7RCdLaGidPnoyVxSUBlSeOH9ccArRCogmgiHXHuiG4Rxsaxj0eNPIISp15sHFhYpvRV5CWf0e5NVoLtWg9qMbYwED0tpXi+bNnouOOnT4dhXJbfHr1aqxtbMXYsWEZYh4cEHe4w0dmoanzUAzVgwPFPBqDQgj0ID4CsGZeA4opqdqgRR3G466Y4bCQ6cpkvPFp+Pjjj1Q4QEObmEgeDZJjaIr+wYF4/AgpEUymF+L8ufOxu1eLjz/5VDEBcdXTZ0/NaAdU2dyM0ZFRxWOAFRQteM7If05MTupPxpVrYE1yH7B8kfIZPTYqRjaa3uwd3Ecu9lCwI56hSCOzQ8lkGlDiOjG3VEeO/DcAgDGZttcYz5ZnDrgPiMcYsOufPnVSn8X4UUSZnp5RcZUxg52sTjskHg4OxB4liVa8I5YwYEWLrhOZTsYSCSl8eMTIS/t/Lka7KMp69rkFuMb+xvqAhENB693vfU8eFTdu3ExJp8kCzB86LVtaLFtFBwWG9RUVekLgFesBaRpiDa6f/UZ+CXRqKmltigoa4pxfwV7P/6fCp4r/FNfsm8M4GaioRX9Pt0yR6Xx4+ztvig0poHhgOH71T58I8CxQlAVgLxflD9ABkz2xArln9pHsUdFEwb+Zc2UvuttbY2JsOC6dPxe//McP49jEsXj3++9Lou/+w0fyWmMdb6yvid2OXwzzer+2J++K7s5OFSvkY1F2IY/9Q2ulpVkM/8vfei1Gj03FZ59gUF5QhwwsV2SgzKx3txxFNQDf3JGlsia+Mzz3ej0qFcBPTMwNCgBOvvf++/HLX/06zp4+Fd9668347OrV+GeMbIeHLZuJ8hL+PM2tMZTnXRGfrVpUD6oa8xfz89ob6XamwEZcxB7E9yhcYJadvSooIDMerIvjExOxuLjgNdhWjj/90/8zfvWrX0vyzKxKpADxYGiR5MheLSQjx/rUcy7UoqWwH90dpTh/aiJWFmfjzTdeU/c6slOAb2OTU9FSxDS9Eu1d3drbYIL/+sMPte9znxRCtpAuasYnELYzcYaBH9ah5pvkztyxCsPeHhWW1jh18pQAXdY+xcB//Id/UEfylVdejfGxcXVUcD+MBe+Rx4bznXvBUFxrWEGL5V3phpU/mvyzKFJS3LdRPD/EevK1mLBk5q4lPAwwEXv55wA0JTcpXy+6H4gPSpo/Yq5KbrNqAoUMUQ2WUfBxESxJ9u7vS9borbe+rRjlw3/+UL497Ev4SjCPLS2bPK3qB9rreL4USghrkcJ6/vzZYYcse5V9eZpU/OKcouhB1wHPmHyvv7cveU7UBK5xRnDPSIyxj3O/jClzjEIFa4did+52VsEiEQPsW9EUp06dUjcc8RwxCns5YyzpJyR2lOub3ctQ5u5Sx0AmIfDizHnx4oU7NmHMt7fHQH9/PH365BBIzJ3vilmR/Wst6ozCcJzPtq+BpTGzFCtxkWMyk77Yj7OUS85/IH8wRjlmyUoMisey5E4Bzy0TKrjuLH/Lfm0yBDXcfRUnKHRdvHhez/PWrVuKDxgn5gRFCfxqkCdljL71xuvx2Wef6x74GeLlmzfvxKuXT8UrF0/G/dufx2Bfd0xOjCl3L+HNUj2Imac2UR+haPH5Z/JIOX7iZCwvLMTaykoMDQ3G0MiQ1kNHd3+MTp2Ou7cexmZlV2buSDNdv3U3DiBbqUmezgGUEGoxOTYYxaZ6dJbL0UOHL/H8HkXdeixvVESgGBmbjBfzS7EoDySTNsEfltdWFNdCYOHZcuaA3zBvmBfqapN8mv3reG65+5/OSXv82adMkr0ivpkMY5Nzx8KcexQb6KYGrxAElEhmYC08E87x3LHBXk8HMoXCUoli03bqEExJr7wC7YdIxx6xRrGlKRbnFw59Hjkb6BhZXdmInt5OrUflWa0SMjRWIaWOmovM8tpBzs0dXRSJKeZWyBcMzTslTYQZFRCPNBY0FIQaYL0Bdc//LLWb/+2CniWURFpUx1J2XTlC7Uxvp8KCxq0QBfa4/DGJLHxEwSgVB/IPNDJp/80FH3dI+dmZlNUoABzm/xky0L5KPpnkYFFkOFLE8F1mQaoGPvTVT1b+nLqfVADNOI48sRrdFl/9va/+OxdWXNBIfhHkxHTkIXnaTteMlT8gLBO3stdKWWBrK3WwNwqdGZHI2JXUPNKzO/rZLkK5SJGJWzkncT5obCW//DfndmCNh1JqqVM8P0/GgjhJ8tAU+JPCiUhdCU8bGh6K7p6OuHfvrmKJsbFR5QnlUkf093aLLLSN522tKi80SNTuSq2m7sjNbwoV/6uJ9c33//2NwMW+AQVILPzM2iKxIlhbShqtsAI42FihsPr2MF+jdR1T7Oam6OtGXgMT5xZJAiArkgGIrM/MoU+Qpo0ysYaJwqzhj56/N0eC9zpAdRMgf68MvWDKwvCGSceGYLCB3y0qUdndRe4I1kw5HTLWPzSTtWHSzDWiTb29a2YLG6iYcOWSjCKHh0dccEEDGgmgCCXzHKiVrU2z7Jtoa7WBNQcvwRZ/5kSSexDjF6MmgKcCYNyKAlzeiz8xxYRRRrEidykAYBDA7nOve9sCNBiT6enZ2K/WBc4PDQxJNqJ2gDQH4FJq2d0/EEjA5ulCjn0RXAE2OGVtvIbhWjZgzZVt7jUfqGzUWffTGvHp6Eubs43MzV750qvgYgI6xLSosaFKK5I27a1ttdA+euJWZzZWm93aMJjnQWBlfT9/TRt6YhSaUW62IEedTKnZ6BPjRuyw5KECeAHrExAHlh8AWHd3p0CKiclxAZMwaGjJg8EEyAXAxfwk4xgZGpZBES30FOUUtFFUIfBPiTHXv7G1FdU6GtLIZbWIrZkBZ3ejJFpXOvSyOacBaxd9cheJxl/dJ40uFZ5XBvGOAv8GqK3v32Bz5OPyyAGqruwj/07BV9a19DM3GC3mchxoTXPYyxQ9yymlBI/ESqZrSVtSknFI98AcFePdAAPs9nzQH50fKlQ0SBhfOuhZ9zkZIajleTNOrG8lIXQGwP6rk5zAsGV9s4aTdEACnkl47dFQ114FaGNZKHuIGChBR78Bwvf3IW1XURJPvJBBayc+ZuVJpq0zSRWocOR7BuJxhwAaqzbPUjKNBB0SDzCPiga6VCxgvxEj0yCY/TKQXDDTkWBW5tCpCAkLD9CLYIXibAvBZ9L2zQmluo4wKexo188oaZfHhecJryxzRSeTNIuTrif3sLKy7HmbDPK0F2sqsp5T9wDJPWtSrJZmnQeZVamuKHRjq7Cye8SOfOe734lnTx5Ef1+P9lK+TsKDwaf8gGr7kqeZeT6rdY23C4Nv7eVabG5say0ye60ZX9Lf4cKw7wvsTsxPTMn5HvPEBWhAF4Pu8gCRxqzN1DQ/UlCoYpuY1HRduPsFsIR7R0+4iiQWUkskjKm9XWsvsZtytwzjSxGd4pCeu8yqMeTeOjT/4wKZK+4go8BmNiNMc5jg/Dxjm9mTjW4PB8zyhUmBs/MJ78sKnNWtwV6auicOjjBkde8UKsyA5Kla+q+xp/OMYU1KCkYaqBAH6JC0x5QSHsA7SdV4AWuuJu8bSzI06xok18G4Jq8ieXgkiT8xJAX0OIFVFyb6xgBUKQHGl4Q5yXgDyCtGSHsOQBRgJefI8sKiEpOxY8f0nGfnZmN0bEysW4gXFP7Z45GfOXP2rPwoOBcoNJIsyEdBXTZeH4C39f3dKLdENB9galuO4Z4enQ0zcwtsOiyiOP/yy9Kv5p4mxickW0Mx3mNSUrFABdbmFhE9kB8jruDzAX0kldRCLLCuNf3OO9+Np0+eaP4id/HwwUNdL9IfxB2XL7+kZ8JemyUvmBt8JsAgTG+kn9BF5+dtal+Oq9evqYhDhx/rb2BgUGNDwj44NChZT/Y8STjteayJjYhV+HnALc5Qkj7ABaSyuMhjo8di+vlTeYBUKhu6Z841QJlctJOHlEwu7Z/D3tZWatMeJPZcOk8oSNSqNcVWlvcKGaUTixIHIW3x6OEjsVJZx7TC0xHLZzOXAK85A0hciS/YSgHemYN71Z144/XX4oc/+kDscp7j3/78FypW8FE5djMwZ+KAOqMS69DxhMEiknV+/4MPPpDsyc0bNw+723Ii+5233lSn1O2bt6Kzoxj9vb1JhhONfMehaP1LOkbSqu2SvlDnK1IUhULMLyxGuaPd45OS5VKpTYxYdcuhy8w+gPTk3o6AIQy8hwb7YmtrM0qllhgfGxHgg3Hqk6czMTF5Ih49fSqPCtYFoExXR5fmE5o4uVuw3GqiEO1BJWRFS4WYGBuK6Sdz8c7bV4QVf/jx5/HBj96NYntbLMAEp5vqoK55dv3qNRVrYJUfHFCUpqjSonhexcNEhIL5mAvunAdIs3X29Mfc7JKKzuxDAEbyi5J+uCVk3ZlAx09VXRq8r/d59h3yjg6tHwolYjjWavHd99+PlfkX0vRfXV+L//gnfxJ/+zc/jxu37sg7Aj7DqRMnNXd3t3f1jDlfpmdnYq9GzNilIgPAK2c24wMZibU9OTGprpef//znihtZ94BtSDwALPb1dKq7hTyBufTtb78tyRlk9SgYsM7Yu+Zn5yU7Umgpyp+ktdgm+SnmXk93W2ysLsdAX0d8+61X4va1G3H+9Endd7e6uTZjdHwijp04HZvLKwI1/+nX/6T9CYASoJnYjK8jXbi0uKzPJkdgMSNph6STjdydB7Efm+hRUDcSHeKs8Zs3b2pfZ0+jQ+z9D34gUhaa8HQlaO2njpKcW7G/4fVw/cY1y6MmgDNLexI9qZhPB2JagyLloKsPyIhON3tpkTPIZB35NugAccc1XRpey+QD7mxEMq1VflkUXPYVf3FfGaTn3OVcZw3a2NkEpCrEu1ot/st//ql0wT/66KO4fx+fl5rWH/uDPIeISwXAO1ZEO5x5OTXu4m5m3LJvEXuSS9ARhDcH10F+TDxIUZZrGhkZ1ucgQ0axmL2OvZm5wmcLWN3dkfcE58TcizmN96H8pkB/5N6Ksb6+GufPI0E1q/nB79JZxPgilccZSC5OkR5pPoGrh3mI84Hc7ckZwB5NwYk5R9GFWJmzjPgcUFs+GTrLvberKF3kOta0BhkzxWrJT1Bys+q8yx4/7rbnWjJQDj5AIY94BqlLPk8SeCn2oms2y6byfi5Su/vKKgvMZ4iJ+IxBUNlRp95rr17RWr1167b2k5deeknPkLGn4MW5y3n68qWL8bvPPtP1051CZ97Vz6/GG6+ei4tnJuLx3Rsx2NcRI8OD8fkXV+PCpZcElEJk2GJ/7+mJX//i71TcJEZYWpi3D039QF1ks3Nz0dU7EENjJ+La1TtR2Sbe6pCfzLWbt9VhROcvBVsKtZwrYyPDMdTfI9P4zdWV6Olot1xYS0usbm3H84WlmDp5Ou7efxgbG451AON7+/vUHQbRiqIc+yYvg710HllKjz3N3nENEom6xUVqhKTkuFW5azJy9rN3IMl4cz3EVvjF8LtMLmLrzLYjHiOuZF2wV1OIooOEPYm3ccGJThkX0WwczPUZ3G7Hh6+3W7JOfJ81ghcO8cnCwlJ0dLBHO2+URxj7nCR2LfEo0gFeUOQvu0gi0uXhjooVSefZHDR7B6ioediF0ChMcC3Oq11Q+dcKFZn8y8+aQMo+SCbgXqacDmfxgTymAucTR1+fpCKIcw9zgBseB1/CYPQP4vWkUpKC7YwZOB53sSm/vvw3PuPLhQpdZ7pQX5VJql9DVT18zyzZnQlyrGV1JfwrhZKv3kcee97j8HLrcYjzKR4Wgc8+FYxoJpYKs+NcTaoDh4SnbGie1QIOu0MSfqKBdlc3L3u65mKu5wOhWZbIE3mYTrskM27ZbK8nFfCTRDaxQMYIMyGXIqcl+3ze8XWINcNDJgHRaU1MxDrZ3IDsYRLe2OhITIyPxdrqsp4BsUkpkThQF/lG+un3V8Q3X/l3PgIX+weVSEifdXvLZljtmDMOqe0eZqWZxzYXJsBvKbbG82fTSaYhoqu9S/IeYpgCyAvIb9c+zsKWDM/mhj5DzF+Bowkklc6k2zlZcJiMdpLE1Wpx8cI5Bc18/szMrJIWsRar1n9Wq+dBBEAVRng6bJPGMEwBPs+bnY2eM8O0WtvTfRDscL8CUArudlACF6F2bQzYSCho8+VeSPB5P65H7GLpkx4owOd3zQzZVysoGyb3ScsvAADB07Pp5/o77eWY3vFZBHUEmASSoyMjMgJcXsbo65w+m5Z7qqkYeHOIbW1XolajBd6VYwAPxlTa9JLiMDNbwQVSGUm38xCkgn0jsA8mqCvcZsP4IBWQkKWF8qauPdvf1xgKJP+aiV+wTBIbOQERBS/mVm4RZdzaOjoE2AAoECxZ890dFbylwAxJUtmsje8BTmXvCq7ZBYxmJUncOywJ/mQ8eQ8x94oY7bqQBkCAh4Wfa5+YUgRBzFmxPJOeKWNA8jw+dsxfAyAlKG5rk+4wnT4YiBL4wlTcAOjppo3cBmO8b/Z4cBcRRSPPu2ykpHsCkE2AuA/h1BIp5kWj+KDDkjWUTJ0dIKWARQei/55LFPk0/32+hn8xfxZgOWOYWWaZHc1ay4GhW2VDHUO8sm8FBzedDzz/7ElCy6UZV21KajJzzYFc4+XOiK+bOJaPoICHBFeWUzKYbzkaQDleJIi9PV1HOgAcnIg1Ila5i2UAiQ7Wd3QZanOXRI6ZvoC7ABS8ZH6ZZMbE8kr6kTx3QmTJ5KgYZXkaQFjmByCzEpAUyPi9rZ3K/CZYJBgBQQOQY53jO5OZ5KwRJKIMCKe1Jw8L/93t/TUxsZZS9xYgTZ4jvD/zQaboHe3aS2ArWnrHMjp0g+HhYgaI5wDMQRem/CzoCHNc5n3Ahawvm7N7jD0ftU62ttTpoMBbuIHN6viP6wUkwRCXTiYXmmzmnI3NeD/YxQ536/HixYLGDmmQbIrLHsy8U1dcWhcNjwonQtwDgAjFbG5BMjY1S0DApIatXq2SKFPcBATJrczJ0S+Z+dlc0jrjOSEWKz4nXEnii+vXHpQSKOuNpmQuP/9sWi+maslt3hTjqxhIOgmQp0cyeiZJzV02krejkJDGk3FyR0yjQMV91uo2ftc5U+d+AYcdDFNUVUs8yUwyb9Ma1uNmTdk3ws/aWquWgvD8sH6/JbQo+Gcmlv2fWlMCagN2nreemZhEX5YNBDwR/pwSIz7XDFGKHPiCQAbwPGNtqJDLmgc8Tl4dWdZQRAjtMaWYmjoeq0sU13ZjYmxCwA/gzclTJyXtN7+wFKfPnIz6PnNsS+cAhbJF9MtlJNuqPZ31RUGAc4p77KBbdG8r+rs6YurYSGyurmpP367uR+fQULR2dEUJ8+jd3Zh5Pi3zTViM7DMqdG9sSsObsV9f24il5SUBXuMTE/HRhx9JRoP7Hhjs17xYhWU5OBiPnzwVqMEexJnPvgqwL6Z2dVeShYwL+5e6WJNHCEkO1z0wMGCtfKQQkTGqheQV1H0BwQN/JvlkdEvHlp/nOiRPglQL3Ul7ALPdWpMAQ1w33lwqtCZjU/mR9faow5VuQ7HMCk0x0NevTgzAL36evQ/Phbn5F9oL1WVBR0Waf1maAWmpykbF0neSCvXecmx0RCx92uAhFxCncT95jGC5nz13TqApZ4/JIpgwEzMwhyC+7Mfrb7wqTzHO9NWVNQFUFL7pgLE/k9njJrMYDMHEk3VJIYhiIC/mC7Hte+++G7fv3Ipbt+4IhNbZIU+f/fjxD3+gc+lnf/036uoCbAMI9uEZhx0GkFV4P3V0NTfH5ta27ruCsXdzAR9UAZrI9dDlw7UAwjPOAJPEbXQOmCG6H0N0tuxtK7mdm5uRJxCMWfTIu7r7Y3t3X+xcuj4VOx6EClMUt9A1Bqhh72M/QsKKYmCxBYAo4v3vvRFR24t7127H9z/4Xvzm4+uxtrUaJ86clEyV5jm+O00tceH8ufj1r34VZ06d0rj19XUrfmatY9YMaCoJlu1t5RfZIBiAf2bmRTS1FKO9o8sdaZKFsUmqCCrEcAlMZ37ArGWOqhst7RfMPdi8jAt7F3sTkglI1fYNDMaf/d9/Hm+9+VqcvnQx/tuf/XeZW7986SXF/RBqiB9YD+uVzZg6eTxOnT6ldcrXWJOcBRT72MtnZmflRcZaBOhnbQG0bm6uam0BpBKbMmeIPS0rNyJJ3NHRsbh85RWdIYBm7Bt/8Zd/FU2tJT+nFgw0AdUA4Lk/wDU6oXbih++9GU/u3Y8zZ/DAOYiOzm6DfMT56azCi+XBo+l46aVzcfz4ZFS2nMOwj9G5uLRM99m25ntbW4fjVXXOwvxHRhVfvh3tSyqYvpiPhfn5eDr9PParxON1MfthmiNl6y5iupsg8diYXR1jGG+vrSnO5JlRvMznA7mawUBYz7lrOMeKJlOpo1rdfABDUGgMoLpj3PF/NkrN3UUZ9tPZh5+egpVQIYFnxUseW6mABOEuv1j37G90PXD+vvf+e3HpwiUZH9+5c8eFm+5uyS5JUkn/HdirLYW0kxPj8Xz6eeqgo2N1wESe1N3I9bLfMl8AkUVQ2dy0p8fQsCSFKWzzb3fyhAkl8s/blBQT8TAF5NyJ6VgV4g1kFcdoyAjjY2jgOZzrltskAUg+z34rw1l1D5sgkXNay0lZHjHvfSYBmggGlktuTzG74WOGZKqJZM57duWRwftoz4LdDuEsSQYR3xGvcDZw5hO7kvcddpozl/bwqLTqQc6POJu4FjOM2e/xh8MLy36W7JOZRMXvqgMf370kWXbmzEnNAzpS6JChU4jPf/zkiUgmk1NT8Xx6Ol5++aW4dvWq4ls6XOgaenjvfrz1rUtx/uQxFSp6OksxOjwQz57PRHtHZ4wcP27p0FJb1Pb25EGyU6noHF1fXtHXJk4fj531tVhcWo5iuSOmLlyOLz69HtUa4DEyWZW4+/ChjLTrKuikLteDWvR2dkZ7qSX6kHyB1FUoxOb6arS0tcf6zk48nJ6J1jYMuSHHmDQlIJTclecsmVRwD2RTLZPNn6wxzn/2TA6iHH8aTE3HV/IcUF6QyDHqRE5SOOrqPjhIeTYxHTErxQ0XHJiDWRyArjHWDD5GxBXqVqxsCTPi/emwykUKCo4CmhPpgWvjdzvay5KEYt7IzwrSxeaWYn5IbGLzIxeEQkciVqmbISkxMG+lytBSdDF8/yAWV9fcJZnpg2k7ctx1KOzQAOxTB9FXOyi++u/fL1Q4lueN/i2FCmdlKe9P/j1fKlR8JcfO+xkj5w6OrJzgPOurhYqjGbqRBMeZX5V+ahQq3J2h/PJocn/k71bscPda3pvdvZVktVKRQPd2pGDydW+Xf5/nIPxCRTYbxSehJRffKOAl/Idzib0te+sckjnTTRhXyc+gce40rqVhiK18IRWmc07tLjTLCLpQYdwr4ynZ91UYXAtFs5IlpRnXA/xv2T/dpUYeDmanTsDWVsnPIc8LBjg4OKgzhvid/T8XRxh3MIupyXGtDdYR+SX7D7/zTaHiX5iY33z53+8InO+xmTbBBUE+LFkCO4Iy2Gt5ASq5grlJe29bOZYWFg4NPWGbSO+/ah8AJDyyHps6KlpapXdM4Mom431aCIarj0m2RGDUQURfd1ccnxo3Iw/mfWurElKqpATTMiBs8UG7vQ1LGqkMm9I22CEYNiKPYG1wghqujUOMZLu1BGPcAR5BY0dHl5KSygYMo3YFKBRHeA/YIQRC6C7LgFPFFwJInyKw7NG9JQGjSwLQANYASSYJE9rTBFFm61LYKIs9B3gO6ADQwe/ShVCpACq0apx5Jjtbu7G3W1MQwzXQmt3T0yn2tMajgGZvUSwNa/dZrzwHnBkUM8Jo+SiZq4qdxNjCVrIciCV3MNwyCNY41Bpgk1kGyTjg96Z9Bv1hO9Vt1ksRAl349g7Ngc6u7kODVdjNmnOY/qolef8QyDTTPB8IFIXcJaMDMAVQKrLAtCDxTUA8Y6RCBeaWSGu0lxWA0XUDi4OghuQS4zSeay4wMXcliQM7tFyOzq4OBTNIPPHCk6UVlk91X54sG1uV2KnuRrmzIyrIFTRRKKkogRYbHgmcZOKsAy4xiTNwKNaQGMyppfZwLB0sHj3Ec7B0OOHSQZ+9Kvyr6cBNB7+CG4GdBmAyi5y/5xbvXOTIBy5zCwAtt/0KaEzBUdbWBuAE3EF3FHYkCSpr83BOKdFxF9O/VKj4cvnCV09Sk83X8zXr+QqwKKh1W9Iz6Ka2lcS85PvsLTDyXPyhg4m56qKn1gvmoCTftBknTxq+zlgy99x15d/PibQkyRKgzLWRNDFHXaiwvNL+AdI7lifzvuWCK3OYTjACCzSQYU8TTFDQzAUhAcSYZA+w91pSTmstSShleQzuj2JkZquxF2U2Uy5A5uIT9834mLXCmnNXmlq+WQ8tLvTwM7mzRNtKM2UAACAASURBVLqeKysC8xkjwKQsu+Ul3nhS8heBja9rahfrWWHtkc6t/OMAuOy1FFzkKZMAVgODlukjcNvZcbDnBMWa6WZzGjij8AXjkj1eSc+RwqqeOclIKuLxfQWC7M2tgCMwoa1DDfjCM2WNGwBpFGcNdpg1zXrnDLHEnueRWtwpTqSChQrsyZTeBSYn4U7iXDRDeoIEifHJnWcqAKOhrmfoYj3nA/NUUiBKJC1XgeSViolJrkISGDzTtJa1vx8WV/13Aw3J3JN7RarqiIdK7hzgazZiz94s/mwBVV/q1nEHSmZByYxQppbu/MrFhywh4T3ZRQex7BJ71hKPHl+DyI1DgyJafl+kxlSoYm2m92C9imHGPkmxUtJTLTE+PhbLi8uagzAW2cc5uyePH4/FpUWdi3QN7e8CFLbJ+4SE49D/pU5xC+NfZBDKAlp3traiq6MU+9uV6GkrxcSxYT2L5zNzcYDm+M5eHDQXY2TsmFjYt65di+6uziiwnqqA0h2aqzwHAEnvG3sC89BG57kT++QCEfss+6j8bqpoe3ek7tK6gD+SLMDQwaGBQ1IHsQfrhD9hrou4gbnsyrLP2STzhZzCzNycGLs8W4gBxDwUsNY21lVEJKkBuEJzfHtrR+ciwJoYv2trh7Jw3A8g2pMnT8Q+Zj7Pzc/p+6wvdRjW6gIp2Ec4Y1W4QzYAyaF9zK1ryWS1RTGBC++OFdiz6VR79PjxYbGAIgHa5nRvEE8pZsGgdc0GrawHtLbZ2zO5hPXOvs6cqe5DVLD3VXMzZz/AeZ98d1ZXiK8A8ne0p1sL3WeiOtQSg9JFHkuUcM88v/fffz9u3bwh1qr9YdDHL4qJfeHcmfjpT/9T/D9//t9iGXZ9sVVAF2uCmAoG9dDAgJ41gJtJEGUxZ5F4WuAMbW1Ocd+emLyccerKTZ1UPDNMFFXIVuxTj+4u5g3nD6Aj65ICBp0lxJmdsbJWiXpzS6xtbsZulT2X97BkDV0DXrMm/8Be55zFxqa5gCnvcHzrlZfj+YOHklg4dfZU/Ozv/znK7S6y7MjnibnfFd//3ndjfm5OOvhnTh2PnW3PBYoijBPFbBX8W+hotDq34o5M5JDPAom7JUJ3dg0ysYbodNCZuO/OK7E1k1Sni/N4Y7TonOQFUE6Bgj3u099ejf/tv/xx3L55Ox49fhJ/8qf/h4pDf/GXP1eB5szJkzE/N6/iEFJJ+/VaDI4MGa5Kkia8P1I6gPAUmui0RT50atJFMOYKn/m3v/ibeOWVy/HwwaMoHNREhGGfAkxzMYy9thgvX76s35EHUIQ069k7unv71FmIr4tZmUjouXuT/a+5cBDjI0PSaT956rTkGdlbpp/PHHr84fMF0M0eNDY+Evv7zGHYx4C8TbG6uq45QGzKZ3L+sNewT1HUBRini4IOAPamu/fuCSghVtL+ks4UOggt+ZnkmQ6pwSnqU6eBOzAFlmUCDnH84ZkKazrL0JpYYcKIJV0zc9VMCC9N8p2cp1gO1h2yInokWVo8qIivfMaJu6JrZY7wUueyZMO2U/c5cQRzeV/PxKb3NQHZeIvQ+fn5Z59rX6Q7LJ/1FOcV4yRTYohmMqxubVX3Gh1AIjPRJQWjfRevQBd7FaviRbG0rLmhzorh4UQSYYzcPaKuQvkPVnRGkGe7Kyx73GUQ1fsR+yudQBRx3aFrny3L5a0rvnG+bbBLJaBEapDkZJLiy/mKGNHVqua5jenL9ntMgDX3rs5dScnVpATA+URcy5qQP0Lq8Oc+dL4naUfDon5l3XmBfMnM25Ka7pCSdGFi8lNk4LlSHBHh5qCuucwzZR6jTGDfLseW+FMQE166dEEYBNfPmj537pzua3r6OTSLmJqaksThK69ciS8+vypPkUuXzkd/f2/cvH493nn7lTg9ORjP7t+OrvYWyT/evXc/BoaGo39wOK5dv64CegedM4VC7NAFWSzF5x/9JjrKpZicHNc1zS8uxfZeLc5cejU++uffRqG5HMXWNhFsUI2oocZQKqszCJIRJE9MpDHvLjZFjI+OqFixubYuyaKZpaV4sboe69tVr+NtOiUoQIPnlISjqFteWApjaWla+ZdJ9cEEHx7qoSyUwH7PS8herC3ybGIi+2GZtCKp0EREwucHc3ukCYnBuPbD55DOfJYecTtrE5yjp6dL8z+bBhMfMe55b8xeEJng59qjpcG5D7r4XszNqhjOe9OJyf7A+cvaYY8vEQuwfyWJcd5The7Wss3Lq7VYTJ1SNO58Ke9JRZr8tUPA/t9QqHCunaWfTPQU2Jz2wv+vhQrn1D43M0jfWEGNuJq/IScoyXARMYz5mOTlOD1F6/6lw6JMxu+T90XqaD/aUdFUSAVgfcjXkw7zHqviQvK4tWyf477855ev+F/6l3+HvSn769h70DJe7DGal82eQ0hKQlrIHhXsD+whLq4cwVW+VKhodFCkspDPCXV2uaO84ZHh++B7h3nkIcHP8sB8jjvCLIdtGTo/f+JsdxRCznZuaRlc55vsQZABpqefqZsTsgVFRs5l1mG16q5fSOUUxqefzcTIyIBiaElJ8txbRt/6l5/Mv23Uv/mpb0bg/1cj8PLgiNo7DfwlmZBym0AiEmU2mq7ubiWJLFDaVJtaW+LF7KwOKFhSHeV265+jz55aSs2shw3vA4SDEYYeAaPkPaRpb7DEJoOlWF3bjDffeEVmUfOw8fC86DbLSsHSzq51Rau0Q1mqpLWV6ipmfQZ2Gv8Z8CDo7O7sSRu2Ow729ndjbdPttwS5nR1dYutR2Z9/8UKthEhHIBuxIhC2OcrtbTE8gimZGSf8HIw5Eg5YNrxgU6GJjT4eBR/GAEkpggcOY4JYAoXJqUmxstCvNrulTa3FfT09SrKppg6PDAvAun/vUZSKbRofgDSMsDCoErCU/A64T5iSOaE2eOsKtNkAeSM2QJfZg5KEyiwjnWC5jdGJewZvube8mXpDNZP7a19KKKxvS2LX29OrAJ3Ple/JyqrGE9BSgFRixcm/Y89VZg6gbMjaYHUkM6+mFExLHsqMbuagClIUO0icpG+7rwRBVXYZhXYrGKO1F0YYiTqJBwPAJk9Rg2cA26uXghbJUpkOok7dL4BMEeCFzooIdcpUD/ajhIan5JIw0FvX5xkwtOSJzG5TF4WLPGnsCKQTsHg4jkdYHLkIpvE+0j6bAUKzpV3Jd5dCI3RhXPW/RHk4fP6pdVSHcFqfh/NBE8VzhrUp47TkqcJ7AbKpgJCKLnwGiRjgENJBBmSqos7wTATs/h7b4+ulnxQrYZLd0aHfgT2ZWdzyYREb7/9l7z2/4zzPNM+7UAk5R4IkwJyULbeynCRb3bY72NPu7tmdj7P/1J7dc3Y+zkwHd7u7ZcmyLcuSZSWSEiVKIsUEEETOKFQVUIU5v+t+7kKRpt371XOEcySSQKHqfZ/3CXe4gjc0kQWIIq5TyEl8vEEQQRca5XHNzEGC3H20dgRr+ywL5g/JukyIyWrF7HHfCu1PuxRxWoROIvDeLIEm82vGzJFgWIwBeXTUJDMGzVqsFOky160FZKwCKk9Q3XPDi20gnd2EzudEfIm+nHR+o8kajQfNqUQ7lWyTjCQdnRRNGK1bJezME/AyXpSHUSFT0tZW7RsgsXn8akoj3aamTgqeUirJvgsCl4DNadtexIuQlyKXJDfqbuCYpqTPUXnW5G1zk30RYzufs0La4f8AKyOxYUAV856u0a6IWwmNGh6wHhKjQ40hNW696MA+70mAF6oYC54P+73kadL9hO8KRQs17OQ94fR3L6j79/h9Aku8DfaMoNR9XFwW26+DQhFfUSQBY+b3BWPA2SMqFkgvFlPcihJkl75KpqXyMmA8HA3J+DvKxqUUec6u9+rNBN9LfMxirsRzk256KtYGndiTBWfY8VAkicWfeL9IZsObA+E9o2CepnXeE90wnlNxCE+NXGqGNK4LuS5PBP3MYH8GUesNKb8HZ3GI+UEwrTPcUUShE+tNUR9LfW4CA8j0HEkR2HNJLurEsWMNo14QSBQppqan7fDkYaGH2ctBFuUyLba+6qyByk5VZ7jMvxPDwz2OMMJzo7u2fIuV11dtsLfLzp4+qaLF4vKqZdpabXGjZJ19SDau2nD/gBWzLVZC+q62K5YgZxdxhNCLzNG0d7KWxLSs121+fklxVbGtTXschUBJT5KElCuuK01xgeQZk/itkhotSE84U8iBFaBiQRR60m6iiA8MDroUIvM2X7DfvvuOYhPWAGscNijjDquDIiTvD8qaYg3FMi/A9ikOpLGJBAka+4wVMjfoevNzkKyzC7PW3dutghJwyfWVdRseGFC8SBPzoYcfVszDGbxVLmnO+drxA4nPJqnkrF5dXrVHHntUxSPMhiniIffJdVIIvn7jus5QChfsgfIW6e7SfKMZzNwTOjlJLfKegBJogiEz95WvPJp8FDbto48+seWlVcsXvHGdx9OAokmas55U+1rBlwMZCYFZkuzZC9/6ll269KF9ce2GGhW8GMNPGmY9XZ32o//0Q5u7M2Nv/+Yt96BhjeYL1t7qjV3R9BUXYSpcF4sA7wgOk+W1DckOIX1GkRkkrgNJfC8AyBJm1dLir9dsZGhI0nqtrXnb2kT/fsUb1GrQs47z1t7VpyYIzbosRtZVzjJHt1d2OXMoAiCl5zKUrAXMULvbaNrU7MGzx+yJhx623/z6LTt2+qQtr6/ZW+98aMX2nO1hSlrC46lVjar/8z//nb356zfUNBkdGRQLlQIkBqYUOWGjck9xbpNPSDYtk/ymWrIqrFWQRNzFY8Q1z2WK29WpIiNzHAY1cwsgD0VRzjjFBEmaUPt/sVWeLv/9f/yDfe1rz9qxI0ft9swdu3L1mp06d07NmZ/868t2ZPKIPfknT9jIyJg0Hs9/eNEufoQR/Z7AKcQBnHc038kJOMOJCfFIYi0gG8M6Gx4Zss+ufCxJhnfefseuf3HVnn76KRVJXn3l59bS4ucCTcHevn5p1w+Njtj7H5zX2qXh0Idn1KY3KPni7OJeib0OHzxkV65cJsqywYF+K2GSnS1oDbBPdHf3NGRyDh4+pEIHhdnu7qIXXHI5W5hf1jVgqL6xXtKc0HlBwTIV/MlxHn/8q4qTP/jgvDOq5MVQduleya/SgHOJHz+PXJJT60dI3n02Jvse+7cKM8RhoK3rbh6q4o88xjynkpdEkntlnYj9B3I1mzTBkaTNgP4H5Uos6IxrmsRxfvK+FKZhGYi909amswAZRwExEhOKdb66tqJnRxOv3uJrEQndiMuJycjpnnv+OZ1Nb775pt2ZueOMWApYuh7WjOcavd2wzW47WDdjyiMpPAM8kD/Qxqb2bZlNl7etv69fzUGYd/yc4v6xY8d0LnDfmxsl7RPse65q4AbRIaPF+Ee+yzUBsGOMnV3puR/3w5mL/BgxrvxPshiRE4u5ZFWsSYEYxBD2uAbpp+vXb+jM4VxmncOWxXyas97zRS+w6fMSOM3ZGg662Np2A/SQ1oyCL+A6xk+FxCQ5FDEPe5vHKgksAQOjtagx4N4AmjFn+EzFmjX2kQ41OuVT1o4nkANFiB05H8kJHnv0EZ0VNB0Zi4ceekjxGI18rpUaALn8o48+onuk2Amgrbu7za5d/cy+8dwTNthdtDs3rthAb4f2uPfeP2+TR4/Y4PCI/ebtd8R6GTlwQDJund09useVuTlbW2HtZdUYWFxesbbOHhs/dsbef/s8Dh7W0pIXcKfe0mLb1V3jKfBvCv6SWc22WHdnmxXxQ+rssDbOhVLJ+gYH7cPPr9jNO/OWQQKtCHisrnXCHBI7ITEbFMcm2WRJNPGeXd2K5XfwdMnnJCdIHsskBuDDMweIxnkBgE8Ag+Rj4qoM3jDTPiHD65oNDgw480XyOzQdnDFZgVGs5ogDjPwIRYIZ/yoa65giu58nACP5bqq4nhDwkjSiruSKEORVfd0dGp9eGbYXBRog96TZgQIxOY4ksWFSAkJsa/e1uIU/VLuAJlvlim2Iee9m2iGBvc+O8OtMte1Gs8Cjr98v/eR5bdRLXFZVe54kuO/PqIjit/ZQJIgixwr/z5QrNyShf0+zgNOc3EqNogR2UH7elJPfXcPxT/Lv+TMN6d1oVDizwxlyngDd328i1AH2AZe+o6gpmq43mgaR69777/h+gEgC0Km5l8Cd7KWsY+UUkon2vQ0ACOy0MIS/6zNT7N9oPO2PcHBX/DsCeTo4L+ovgCSZ12o0qcHrbHOxYxJzXNK2icXOPbHPcQ9qZquu4YoakTcyr1xi28F5YwfGBK5dW1uxpeUV1RwBNbPXubF2t34X8ENXV4fdvH5TsSBznDoGNawvGxWNEsqXf/nfZQSOdXZrUYcGN4kZBUN0LdFOFpJJ8hO7XnDHk2Kgz+Zn57ybvrMjDVC0FwnCMTGScTQoaPQuE7qU1xL8spFwaLlJN6ZGFesf6JXm9JNPPqFO4frqshY1i5Lgjr8TgBDckZBywJCQI+8kmYgWilm+WTmqeccPprprXFKEkQZ9pWyHJyYVvM3M3vYmSg0KdJsOMDYU7oENkA2pHVNtaYrXhNCnaREoSQIaNg6CTZoO0o2l0dCkh0+gOjc/p6ANuYqLFy/oNZiuoakt+RQhnV3aBkr76uqyDhdMdLh3JCRIqkjo6K6urvBzkiSCUdDRrs9JwMWXghMFAX5IOUOgTd8jgWezVQIg2SRHiUfjIqiBjgJwqrUjtlOhKx2Sfqj8bqcizi+efXcnhrslFbeYT1wfUi5Qmz3wcEkFDpEoevJvl+FxyZwobPBMpUdLcT1RGrlXkneS0vAmcW1VNzUlyCS4VVKciokgVQ+MH1BRWIawtZqSLxJOBcUqFiKphZ52QZrnFL0kt5DLq6BT2vQkiGsRFpLiNEX5lqzQ6Y6acmPO0DeMojvJnYJ6eRi4/mZDMicdoLrX6PyHkmUikSggbKAUnH4p6RcKe82NiqBUpkekAuI9ptr7jSxnNvGQGQOuT6bCOnndm0HFpR1Hg0k3NCGwKSggz8H4gfoRUjublQzI7zIqktBQc2AVU0jorqLmCcmqow28OMt6p1gcyRPNuuGhAQUoq2sgKWlOUsx0ZJeYQfI5wKPCfRF4T+5D7ImEbHBKsstnUbhnHsCUcJRtVYUoFXRVzMZY243mxMBKTVGSJDVeQRcJucEe2eYyPgkNTpLaDk29SjO24LrCLdCZPeBDM5/nx2e6gbx763ixkgLtroIX6VUmHxcPGPfXH3+nZo6pKkkF6DFeG+g4GdtLZ7ldifP42JizYXZ2bW5uNiXBLgfUKIyrIODID0+8veHAnEAPk/VDku1hbfgvYCDNnsZYkyR5gM8eRRKhJoGMYZ3VwP4i+YSC6+aCbnbvHU962Je5HzaLoBPrerTP+fwAjcyzVdG75ug79n5nwLgeK7+P70IEh7FHB8omGrr8PLRFY22S4FqL+6A4kglEL/Jc7Be+dkLOKnww3KAQeZe4Nm8AchYxblyba/E6CnS3vqP156aZrLOWJPngzaNARVFw8j3Zm1kqLIqZ5c/KkUeOKudcVhM6TNDDj4bPVIPFTcC5DxXQytu6P+YlrBaeEc+MV9LQV1MuNSTcYNs/i/PEEUvOnnGWkxvOhskl78U1KqhPyV0UP6LFytwPJlcUL3zt+XsyZh2J4kwBe3V5RXsOhUbOX5pgp04dV9EB6RQa5Dyb9ZVVxTJIInAesB6DRYcmOHEDa5vCeHdb0Urr63bq6GF74Nxp+/jjj21+ecVaiq22sLFl3QMYoq7L0HJ7fU2IYYwvSfCRrfPrdBNLzquFpSUVORkrNPLZh3r7BySXw5gppinh4wQDB9kdfFLqAjdQsMXPYKC/TwV3yTIgc4NmPz5YNMiTHw3Pm/2ZAhHztFqri6EAQ5MpSsMBtDjXQTwCI4V1ePPWtB0cH9PZzF4GOIKGBdcFupemD+PF9TCu7H88WxrTPX0UODijMyrEbyN7NTJsPamoK63/mRkbHh1RIZA1gaxNNOhu3rqp+JJ5wRh9/evftH/68Y81306fPW0zt2e8YR6sInmeuGQTe/WRo0dtZmbGQQn4GcFg3KYpTaG+RWyIF178lj344AMag1s3p+2VV34mtgH7HqhnGAhO4feiG/PAG0VFxQCsV+ad0NDVin3jG1+3ixfP27VrU3otX8QJlXLJOtuKdurEMXv2qSfs56+9ZrduTkkfPJOYbDt4qW1XVBhlG93YosmStzxG7zs7Kl615LOKh2FzUqCKM4W1zdxQY5umcr1mR45MqOhVg9XZStzkutfsxtxfPo9US8FKlR3bru6oGMO6lVSQ+T4thpSAK244rCRfMlfb1pZrse7uVquWSvZn33xWZ/9bb//WvvsXf2FvvfOuTd2Zs7r2NxC3sJU7bXRwyM6eOW0Xzr9vJ44dETCJ98P8dBzPGNZ40hDnUrkeroNYSExrFZ+RgnGUrQy0YUkk7yTmPv9mr3LZUFDwGCjjW5dTM5LiBGcbRamvPvuMLdyeUZOtu7PbnnnuOfvxv/y7rW9u21//6Af2yeXP7c1f/cb+9u9+ZAcOHlIjCBDWL15/XeN9+sQJ+UgIkZrP2+LcgoriNHuIVaJox95x586MfXblshDYZ06dtP/3//m/7cmnnhAi/+ev/DQxHijKdSumWVxasRKNlq4uMYeILVnfw4PDdvv2jEBNw0MjAj2JwWwZmcV++umnNjYyJHYOkjU0/SlIMUY0CcWI2li30lZJxb4nnzgnJDefx544N7+o62fsVpZXbWV1TbEa84BmDIURZCZZW/JTkTym5yfkI6wDzmWeH8wP+fxQqEloX8WMKTYJvXCXHwE4k4BJGTeYZg8Cwa3fRUu+rcNjIOJPS2dTYiZRVJdEoZDRnImcUa6J39ndpXN7YxPGVbd8GjhbkRFlf8UonX2KXA32HXssLB2uS7r17R22a1l5o3DWwTphDcmsFSBUR4d95zsvKc9489dvyvxaPmMJuEM8Io+IQlFznq/wAOOzXGqqXQV21jRzmGJwT3eXCktiDpXLajrRlOALqTsxphkz5PUGBhXfCUyREMURBzHXGQ9iiogd2btZC6xp1h7SZMh4cV2sQ/kTqYHumvmeD3jeF+wymrU3rt/Q9TNOGLl6kayUgESuF08sJrADuV5XV0I3u+wysbviLOIC7bn+XsSOxHIUbTErV6MsGTRzX+4h57Km/Mmzljwk0intNPldYixkwJh35Oh8BmcP64B8H8S9GE2ZjD3wwFk1H2EH8vuPPPKwzn0YM0h/wcKEnXhkctIuXLig+Ofo0SNC69+49rm9+M2nLFfbtvmpazY2PGCDA7125coX8vo59fBD9t7b76rBPT5+yD78+BP9Lg1E9g7iinq+xTaXFm1uds5GRg9ad9+wfXDhsmUy1C4KNnVrRhJEm6WK5ITB1gCCQ0oQRsVgX491tSGpXLCh3j7FQPSjMdK+Nb9g2QJSbCV5XEimsZt6BGoPeOC06JyHoUncQBzKHBZQDSN7znIDlNqlc491Ljmt9nZnARPrpWZmsKNC+iliO+Kh3WpF4ArAZc4ArSrnBwDBcyRXdqa1e5twNre1OrNWIDVYQ4B7AIJgcr1VSrmUA5d4vjSBVMBWMwVzbGeND/f3KSbTOU6cVK/b7MKqGiGKj8WK9riZeAmZLprta5uoI9BCzQi9fndB3yNUl87dJxH45XqDNvbn9M/0Im9iOBDQ15YadsnQOvLZBvLd30pxngCcaQ9tNCpSU7DBqGh8tjMU7v5K0kxJijal9+k+9n3ZGjCzplKOx0LRqOAVrlEicE9DDtj9NZVaNWoV+9yOkPGOHCXyo/DhuF9T4vc3KprH3vMu9mPV4dra9Nw5o9jLnbXcqjOEOQyQIZrmqnMl82y/D7+6hnn6vSyT9HjxHpXEdWKGkKMyIvE8Q8bLG3YOftQzTjk6a6BQcFlyz9GSwkXGzc65EM4o3p/7Yf8gQASYIQZcsai6KWcp7DRiUwCRE5MTmufs8+urqw6mlaff3peNiv9divNf3sf+CJwdGJZcgqOUXasaxB4ocw+eXVdN9CUxJNgU6ioui/a/B/3cER8ETCSzIMKcHrXnRmi5FhWKlhYXPehPUhAumYLZLMn9rp0+fUrBB4WaOAdC7iKCKT5bxWrQV4lS5WhpLwyAYmOzIEECHUDwiCTB1PSUDsDjp09IIxL6qAKp0raQLzRFlAgmk2cVOBNqK3QcOdxAXUj/sQKCslObCxsg94y5HJsKgQDvQxAnw7vRETf/UnDQqk1paWkx6cuCyKnJuA7pIZCFjJfTyd1cSkW/OkaDFDXrajyoiIT0QpJvYmPmUBcalcKhNkJv2riOqdP5JA+TmhOBtA+EaUPiJG2yamDc3XZvTBySy1CAEjpgj2DSC4MuS+BmfARHBOYKugkusmhxbsjnRAe/5EWcTcHzJOD1RpcX1xUkpKKAAujUTZd8SirMCTmtTZoQNenQUgTeRh81b51CaVT0TA4dOmifXv5Mz5vf29xYV3EupMF4ZnSqKXbw+RpzDJykKb7aSIjQkGY9SONXETX3hYSa665zIUHtAx2oYl3yR5AcSjajAhXPS3qZSX7LkUk+fkRy0tTVmZo8AJJ0ExfVOHiTfI4X/5oSmXh2KRDxPxztJm35JI3E7zA20axweSdf91p3cZwnyjz3wlsrEc3ntCZIwkSRFNXa0fbNAZQCkTRHGglRGGCn62YtsY5IVHnmIGZUUE0FGLEcYBVJm9QZEF4wCqkzL+AKNQcTDOS/EDYuWdCA+SeZJOn8gmKX741TnaV9nNDcJE7MSRUTkzE2gTLrla/wG1DBmMaVfGG8GcXf1fBJUmnyXAkUWCrQ00jBzwaDLOZZSOCB1Cde1Fqo7kgvmoKCMyX2dZXj8Wrt5fPygwCVRyOT4kUKrbUPC31HYpgCPSFXq1Ul895M8OYI+6+j0ZzpxjUF6oPnS+n3BQAAIABJREFUEE0ZnjHvp2ZIYjm4t00yZEznhQf37v3g7AVnS3jR2ufQPgLTg2Qly+xf7CdpHAO552gUL9C7DJa/P/PAEwJv/oURoBgBqWESyD+egy8pf1Yypfc0RWcgiQpnIGtbSUsyBwxUz36y4eyKaKS6bBrnlyfM8ozgXEzsF85YCiuscdD+3mTI2V4mGjgUq5MknAJr9hD36iHZjUaFN0z2pfr4d6B0SOa5Pi/gOX1ZP0v32pxsCWmV9Hclp5gaJ8xvzn++vKDudPowfo9zIxpbYrIkGTtnf3gRV99Pkmr825vezQaFwfRwBBNfnBUuS4hsgCNp+YkaIJzrxbziBMydiU9AMJKguNnySEPSiEIuxWoK7zQq5F9Qq9nI8Kj0o4lT/Fx3A3YSkM7Wom2urtnk+Kg98fhjdv78+7a6vmEblaqtlXdscPSAGh4DvX2W47lzwTmQ8zsqgonZUvCCeaCtKAzRCLpy5YqfjSrAgmROhu9iPLEHeYOJBg/FnWCedna0qTCpsyTTon2CQrMn0/5FUuM085wj1zJZu/jRR7pvPhPddfcV2hOLEEkoijckTyD3QS7SxEfOiYICE8fZiFtaf0g+McYhIbK8uGhdyL/t7FhHF4VXsxIgAOSoNrbs3OmTdurMKXlytXV32e5exqrlXfkkUExm76HgilQQ/gAUzP78r/7KfvmrX9l2pWSDw8MqBlIMBjgi9hCNvsQ6WV1bVUFSRa8aspjuy0CAIelFMTrdmJCklrhLxU3MgFfWnNFEo7DgsjTRyBfyU/GFy0nyJ2eOvEJoVHz9a3b+gw/s+s3blkvv0VbM295O2Q6ODVhbMWtnT58WY+HVV16zInIUFOHZ+zB3hVmXySqxpmBDobqto9Pml5eF5iaOiJKD2KEUqdqRBcnrTBNaGtQr0pSdHVaRQXxe3lkw1pgDwcZC5oqClVDcPb0yLWWsKMoRu1A8krxG2huFItVeWrNiQiOjwc6J2pbbseefe8o++eQzW1xes6MnTtpmZccqSK5UK2IZceWt+aKdO3NajRsKVsRUvV3dtqzi3Kw9eO6s2BqlJDXIGsfPgeIQzT4Ycs5i9OsWixPmR9l9WYidWQfEWCqy7vJ3fDwAJ+TFTGEfAAzEvKXoy9pg7rz809fsa19/zopt7fbyT1+1b3zja2IWXbh4Sc36b7/4bRs7cEBxQhRiPS7mHHZvKcmKVXc1hremplTIp6HAWtILM2ad7UV7/rknbaCf4rnZ+Pio3brpsmaFQrvV92iuZ+3lV35u6xtbYlcjI0XsA1ND976+KY8Bml3y4Ut7JsXwfNYkoTo0OOReBnPzeobONGlLQDA8/WbSfmL28EMPqAEhBjngrXI5oZ23VcymeXfm7FntSaub6zYzN6ui8ALFzxaeBZJBzMFsg0HAh/I8dBYmI14PWSmy+Rnve76bJbMeZUgOQCp5FrjEpRekQ8InzrKIDxRKE8+k8yHyGoo2FP+dneNxAnPI398ljbTf1vaMJiFrRk2JVJyl2bWJ9K5YiuQlFPDxSYIB4nKmgJR0Pragfd9uzz33nFg67773nl27dtUlcFJ8Q77G3oESAONIbEX8yWcKZKGz3ONCxoNnwD2Tt5E3xj5FbM09AaYTyEA5BgCMotQMuCdkvAD0CcTQFA+ypxCnjo6OqtHLnGBsaYTxOmTF5PWX5NPcQyqZ8zaZzOpYy+WtV0BBZ4B6jOUSfDyLLeTrEiOfeJG4NHwLWAj4mvDMkc4l74uCq4qEGlPP5fhivHkOHtd44dxRyvvSMcRpjAHzMGTKJBWWpGSicOy1U1UflL8w1qUtzMAL9sC5c8q7Z+/M2Nrapj355Fclo8VaoU5Ao0KSgyMj9sW1q9oHzp07Y4VcwW5c/cz+83/5gW3N37TVuSk1Cvr7Bmx6Zlrx2+Hjk/bbN39rYwcO2/j4hH326SfWP9hvvTR38N+heZo1ybZhfJ/Pt9ro2GG78NFlQ3WpkO+wxfkVuzk9bTt7GVvbYn4U3fQ5YzZx8IB1txdtr1a1XMue9Xd3WzaTs+3dms0ur9it2UUrtHVYdZe8g70cfzpvSpUqHnMiNc1+qGZfkuEMWS7mKPss80fzI4HOPD5ygAFrT+stxeXhCRp1BnnubWw2ajo0jJHz9ZzY5EOxBZg1R6PCA08xKQCzIikFcySflck9fk/aRwBn7XpDGxUNmBhiIu6m6+Cs7miz9dUNay3kBCJpL+SsF3YrTV487GBZwu7LITflni/MX+KQlnzBtspVWy9RgEaykmtzOTsH7vk8jJhX9ZQU33oO4efyfky8LzEUv+dNQI+Jg4HSDDRrBHLe27gLhKafkd8l03Mvhu+vE6/ZOQM5fN3EUEpvGtcVcXiAUuPa4rriPgOYu8/Y/v0qCH5tnuV7lB5gxCYca/p53GPzWDbu+w/8RaDOJF3l49zibBqY4Hn3tVNum8u5tHwRz1eUBUKiz9ltuv/E7r/74+6VffIILK7T7yw1NhLjlp9HniOQYBr/qKtFjurNWRrYDiKLJi1/B+AVqijK62v4xLSK/UeMDxhneGhQe4B71TmrPIzn2VtRBgGsJc+jckUxvKRMv5R++v8ztb58zR/TCBzv6hVCiQJKFNpAuKHzBuqfoIJCPgcFARNUWJICgnuKKmwUIPe8yO/oE9AbDX8DqMJFaI1lSQ2ApOBA1MJNZowcZF959GEtOgIw5FcoJpFQE5REIRCUGQkPhWz0Q0lICBY56KSn+sVVdeR1mGQyNnnosK6fZPj6zRvyExg6MCJmBAmHzK8IfFpbHdXYkvXPz4J86rBr168nn4xd6cWxIaLXzHsKCWbQjju1qRCQIVmAmR3mtEJIolPb3W2DgwNKpEFd8TUxMWm3pm6piMImxYGIyTZSOkJRE5gWC/qdz658ruvjnqF2ib7Y2qbNmgKJy+H4Qc6JASo89Mf5LDY5FdgSMud+h2wgx+Mwi8MttMj/0HxuLkrJMCnQ3gSJaBQTwCZDbyFZKRxsb6v4LN1witTJYD3eK5gTcWBEgZdAX8VT0DgJmcOfdNFDuz8OLIo0NH1oSLgUUU1IO8acA4+gn8MMZBOeEzTgRB+mSNPZpufCXOUzYRxxncGAWVpedqNSGXLlxN7IFYsq1qvjng4l6OEuNeOHVAQqXhB1/U8hwVOg06B9psTLNY29aRA0Sk/+vJHH5zTTGqMgH8XAu4KhpNWb4p7990j6stLAF03UfSm8gOz+GXofFaODheBa/6wZ+YAg2aRgzGn8zs7yBkdILpE8KrFJdMnQqAYRyNpinJmnrOcYL5legw4SSpyEz1F5Qfkk+GbfoVERRVBPWpsaNngqtLt5VXztM4gcBULQwLPl3gkS1BhLjAtHpyI9tJsK+bvav/aDmX0dUiXXSGJpv8QkdsebQYnaLiZZepb8ncYkc5DiYATGIb+n4L+6q4akXlfCxN3XMl+e0Du7RYZxSJ9JLmHf/FvPhCZgSrjFNpMGs+unIzkQfgXyHxIqeVt7ULNPCnPQpdnwA8oJuUkhCQ3lQBFFs0EyL0j0gDiUJBceIDSV3Zwv9GzZr2MMHSXkqD7dV5KECy8GL3j73Gpo1kouwpkZfIVMgPa6tDa0nwny5Kgniidq2qYkLRo93iR0BqB8GpDXEVvLZRFCjsjXnn8mr4umjEsnMT8cZSk/EFCIWgcg45jbiR2g/TD5qagSn2jEib3Dmera3/67XDtJvJA6qRGrpKWJneD7ge8vFPf2GxWco4lqHAitVPRiHOUrlSSkmhMynj30Y/azSNacbefzgOfgbBKXahKiLkkAhCxAPBvdf8NM3Rl8sR/zbNi31cxJBqWcIJLj0f6xP19IWrlv9LdhxSHLSNA+OTmh4gPzaXJiUvs7hcSjx47Y1pYbTPvzdWo4Eoryf0JGUg1LL0xzM22FnO1VKlZsMXvmiSfsxo1rtrC8bOto05erVmzvsly+KGmDFopCrJcdCqV+lgWClbHkTR1pShKVtdnZOYE7KgI/uK5uNGIdeJEkAjVebvIMeGP8wKgdGh9VoVvF22Kb1qcbJvsa4tpp4Mg3RvM7Y7emp1KhtktyFqBhWd8zM7Nia7LPrq5u6O9IWK2srghJuri8rGcCo0KAk2R4ShKls5yG/NqqpI7Kau7mVAiiQDDS32Nzt6btsQfP2elzZ2x5dc1qNH5zMIgcLLgNwINiCWjm6o6VtxzdeeDguKQW33rnbRXS5/F5wL9ltyaACzEPrAyKHTICTSABb26v+7qswcT0MWEN9PR2q6At/49CXrItlYozKGLf0vxIkqFiBontmFWRTudoYp+iLfzSSy+mRsWMiprsJ+3FvNWr2/bQuRPW2Za3pYUV+9YL37BfvPZLm7p9xwrteCq1a63QwGL+eRO2IJ8rGpArINWTFCOxtTejHUjAJgNzYmCgz6rlbTWj2UtBBtNMApxBIUuyL/Kqwf+Hgg765G1aI7wnTQrmHY03Cto0F0ryd+MzUlOR65LUQV0Niq6ONnv80Yds6vplO3jggB2aOGSvvfq6tXZ2225L1jYqZdve2bPuHlhDNVtZXLPJQwfke4IUK3OM/f/rX3/e3vjl69bV2a734XpZs8hMIS+yQzNaxpN4xrSpsMWZDWMyfLbkd5L0+jUmCXCDHKz7FTmrEqY1zxDJJGLmzz+7an/5l9+19z+4aAtL8/bSS3+qeO3ixQ/13J955ln795dftrX1sv3Nj35gg0PIIubUhEDGh/MfdsLyMk2JWaF8yUOIW1y6DhNMR5O7aSaNzC577pmv2okTk5bZ29U+wvsUiu1W28vq2f/iF2/andklzXmtfcnxqZ+s5zYyMip5WfZD9mMkdavVshpWSD/B3mUeA5aC7SQ5IcmZeaGGXEONLYBi2Zw9+MAZSUzyWRRmOaNUCN2GVdauvfPCxYt2e37W6hmz0ZFhAXOkqU1xWuj2rLz78POZujWlc8rPLwccqVGmeGwfEMXv0ohRDJQkngDpMIeJe2i4BViHfYBcU2j/5AXIe8PCqe95HBaEXDWFE9tXsmI0XJIcIQ7KzHfAal2MyxasNW9ycf/ESeRYvGYL2Zsaxt/4c5BHOEuU8wxE6+YGBS+X2aR4j5H5U089bZ999ql9dOlDNct5/hS5aYzNz817YYlzhBgI1qJyNBjtAM/c5F3MlNY27bvsMzAmaCazx0smB2BVkh4FKOA5y4jWAN6Jvmf5ua+zl1hbRcys/G1oFLB3uq+Fy0kS71EEJkaQRBLMmPSsYizd984LgpJ5TIVYcmVnwcD+rYgJrOK3pBSdGcv1qMGeSf6QlhH72BsVSRIssW8j3mWsiZ0AIDa8r1JhMHIbccXSNTH/YeYLiEEuIVa0s07F0k+sjZCTYj6xb7Iuzpw6ZQuLCzZ9a0rF6Mcee8yWl1bE3JIqxABsx3XN/S+uXlFeffLkCTGer1+5av/H333XqhtztrYwbUO9A9bX22+3bk1ZtpCxQycm7N3fvGPdnf129OQ5++zSRevp67XBsVF77/0LdvT4URsdP+DAGBj9Vdgn/fbrN9+xTBaUdJvNzS3ZjVu3VTwvVfAmybpEYKZuRycnrKW2Y92dRSvCTCsz301eFksbW3ZtetaKHV1iUdmex5ecr6zJ2h4ShFmZSzMP+I/1pTkmIGOL5iLrLhg1zEnJKpZpCrdrT47YnP1IMaAAV55r8TP2ZDU+yb8SIK6nq0PxhDw7xehD2aLSkO4OLzpyJck2qyDvzYuernaxw8M4maaZ9t4abSjTPtWSb1EdaGVpVXK8BmMj0yLmSVuhaL19yK9tqL7VWuRsxYwdWdUW7b3sr6sbW1aqAhRo8aZrPYEXUkzW3HCIeDny4ua4+ffVSZqL8//R6+9tejTes8HccBCqAwUD1pAkaJPcrPbi8IMIxkOTR4Pi03tY+XFdzQ2V5kbN/e5tv5i//9N9IFKKTJsVFJre5N5GTfw7rq1xjYYcrqsm+B7Av10VxBtk5F0wZtxHjPOGvZ7YNbwlFEPQKE6+PnHv/hn/caMiLltlkFQPiXUSTb3mMQ0AHL/HWqNRwVokR+BCWEucGX5ewzLz/JX3mJgAYFXRGU1Nir0Olt4Qcs0pl6eJTTw7cXhC8oxd3Z1qphMXKBf8slHx+5bil9//Yx2Bo53dSihA25AkqGCVyyuxJVBvI8BTMODdQSWAfX22tLAotAeLDWotiaw0JhuyO1CGXecO2An0cIKAatmRJoE45yDCvG19dcUWFuZFb6IgykKenDziBSFpX3aI5kTzhIT0xIkTStTU4c+0qEHx0ceXJG1CQRq5lYmDh9SM4N5IhDp7uqy8y3Vwv9BNoQlCu61og0BeRQg0jPjyeQX7BFCiACftRTaeXCarAIX7JkCdoaGTCitC12Lw3OaUSTZRCj4gPy99/LGmCQUBqL0E12G2xKZEQZKmBwkXci8c6NBU2XxAF8JcYdNGczqSb4IGgmKSL14HSk466wnZSjBJ8BhJngoPTcW9aE40H1zNh8jv0gp9pjfMgBKFLcSgAnFAEXtzfUMdYhIQCgoUhxR4SauRrr8bGkfxMZDobOZCcifDoUhKHO3syHTmaBzqYmJIN9cbM8wFAuxAxINMBHkIipDr45qYM2ru0OhIBdo4ZJGfgUZOoZ5xB41B487RimUrlcrWjjF3actaZV5WJotLxVtnv1AYc+kGR74SUwTtzwtnrnnvyCFHFEexTveGzEdCtwtBkHwQ9g/NoKL6gc1YhHSKIytIfhPNMBUx9dxSIYbrkrRW0gn1wpib+3pskYpnSImoOeR0TyUDKnAi0eTXTJGEn5H8hFGqBxSO2ArqJNcpg6hkau9Fd9fxlxRFanCwJiIAoR7rppLQgtvV5ArES+hqs0a1n/ggK6HXfpUYI8wfFdlTYhsICAUZKgIkczkVmfFP2VETJtBqgZpgT2TvAIEdRtz7wSJSZG0KgjHZpeEppCNa/TQoEgKEoIS14Gh0R5FFcCiDuVS4YP4yBjIblTQWOraOS2OOR/OOZM1lryiYYOC+LZSeZN9k4O1jQgwfJucHxse01yO/Iv8Gyc3gy1IT00xJiKTWgo3g8yGXA6VFoc1RRBTdXN7PpYy4F0eAoHNftUIrmpyuP+2mteHVUG14MMjDIDV4gunge5E38hxt4gg7NTATZbe5UBG0ALEokiG0Gjgxv33muk5ymMsntpYXq12rmfmjzwQt2tqqwrJkqNC+pWmRkN1eh47153I/khVLDYNiodXPPNC+qYgglltTQ4ENId1K8tXxogP/F7VZKG7X9iUDE6tFmsPONhEjSqbhqQGaDGo5h4W0BMGdpP+0vzY1KtIO3mhUxDrl+3EeyABeesSO5qRooqZXxZtqLhvobECxykA8qtnvDadoToTPRvOa49mwz7ifiOso8z405+N++LwwUIyiJMXP7p4uFdFpMHO+BgIpCkN8DnOYOU58sryCLxYxjK9zziCdkWpy5lTg51xA638NA9K9unW2Fuyrjz5q169dtVn0rfEf2q7YbiZnPT191k/xo4R2/o58Lyh06PlmkUfwwiCJBJ+BnAl73ueff67PQT+XgjFSjhRStSZ46klSj8Iz+z6TA0YIjYo+ySwhtVbwxmKLN4klA0Kxitfiy4BMkeK0gl269ImKfoyBTLdTg4g9jOfD+1GUBeHpxYNt6aNjzsf+ijY3jX6+eFbEbiSDgCZoHHAusrdIEo5i1E7ZvvH0k3bp/Q/s1LGjkr0odHbb9MKi5VoxFMfzqU3jxLpgLlPMoPlAIkdccOz4cXv3/Ps2v7Skz6OZM3XzloqxfKaKjWmNYmjMeGpv55xUzEPhhEaEIzGffe5Ze+HbL9rq8rJNTU3byy+/rGKhF2iRHHK5R6HFk+SD9qKUYPJ3vk9jBY82GhXvv/eeXb85ozGmkUxzq1Yt24mjB+3UscP22eVP7eGHH7aBwWH7+3/4R9tj+QJowYuhznyPJnpOTatVQBA0LuXhs+XSN7CMZU6+Zb09nVatlK2vt0fztbuzQ891aXFB+5n2h5S0ywhbhR1vlAKk6O7C96xmre2dYqH8609fkxSBWJQ7NTFBJZWXd2NkCoHyUwJEsrtjD5w9aY8/espe/slP7KGHHrHp6Tm7PbdAd996R4ZtDjPgLAaWHULTqhiWz9nqyooR+rQVW+y5Z5+Sz8krP33Zzp4+peI5jXyMwfns9q5OnWGSEkvMONZAV3ePni8AJ85F971x+RhiKNYYbKFLlz61Rx97VOelGG3sx5WKZL/++cf/ZM9/7XkVCs9fuGiLC0v21FNPac3+y09+Zt/7/neEQP9v/99/kzzrX/7wh85qKm/bK6++ah9e/CSBTbiXYpK6cilDMSxk9ss1taiRii4666m3u2Df/dMXbHxsRI0Knmlbe5cQxbu1jH3++Re2jpSDNNRdzgIvQPcByotRgc461+YSUBRhfK1ItqRQsIsXLwrgxFnO/sJeSCGPWMDNbNHsdqQr43fq5El5wCDnwxwlbmM9wOCYnZu169dv2q452lpAKQp9PXhfbCsHKm1saVy+8fWv2xX2M6ThYIblYBw4YyGY8H525cSqdqBGTc2n0M2XKW9iaQU7jHMVBDz5aHx5PApDkOZue8NPgc/jS95VFOZS7CqWAHKhNG25GhpgeCHkHIQBAI3COcX/fCvMolVbZ93RQMzCVmr3xifPM18Qs2JxcUn6+WK1l8t24vgJ+/Z3XrQ7szP2s5+9pniLJgN7MnkfORuvlWxOuhfFqi2eb9Io5HP7e/v0fuxXzBniQmQNxW5OxXn2oDjHA9zBXuS+bZ4nsZbVoGrDmyGnZ0bOQhzDmUdszX7NWAFu4wNZb6wtMTYTA5P57CACP4Ng7SwtLQlAyBwF9OUeC8s6Z2QEm0AbwWblc7yx4DKFNCpUUA5wDXudYkm/bsU5xP0JdKOCaQKaBHM5QDBeGDX375EsqudWhDc8L8Yp4rTIWwf7+/UZrBfmPw0c4l4k+2ARASCAnQk7ifulKIjc29Wrn2uMz6DyUKnYZ598an/zn160lt11MSr6u3uto50m4YIV2lqsq6fDrly9bgP9ozY+dth+/cbrNn7ogB08ddIuf/SxchfQ3keOH3NfFhml1+299z60bIG6C01OJABX1QiGDQdj3L1K1m1kqN9st2ojgz20pqwu2ciKmACrpZLdWVoTE6O6w1pwBQAx4rMcOw4GZE5wdkRMpnqNWEjO5HTgiNd4QhmgUZBN564DKWE4IrvkKhGc59QYkN5iTbMHFPNIMu76czf3choaHPBzZ5fmL0Au8gAHMvHZSDqRscKqcJ8Ncr+Mrpm1QuzJc2dNlbYrlsllJNUHOGN1DUlDYhVYyZ67MG8Gerpl2I0kFEw/FDTEAC1tWg654a4em19ats0K3gc52w0GRfhINBX1I58MUFzkhVE7+UMNgHjNvQX6e+uGzU2NBkgwMTFCEUD5lxRLPO8NNjLv1XwN0Xz4fdd173U314D4e3iAxu/fe63Nr2++7mYgYPzO/Zoa9/v85s+Iz3V5ZwCI3mBhzpJThky4wEaWUXOCdc1aB7AkST3ADanGEYyPu5tMzQyWRGlJF+H1oLvvOpoVASKNelr8GXMj7tfznIzOTf6ufBugXAJx8u7VHVdnYc1xtvBz4rHPP7+ivJyGufzq2vGrapVUddQMrly96owKGsa1uo2MjnzZqLjfRP3ye3/cI3Cyt19JmIKZTpJnun15oQbRUmwU0ZK5MkkAmqC3p6a0cdApJBhQd3N3V0hzOt9qbmCiWnTzbH62uLgomR0V20olySWMjA6rYAE9XIESEg170HFrQu8EnRl0OskletT8HU8MFncU5DdLWwbSvbevT/dRowCCt0QLOotuZokW8Mb2lopk83Ou+U6C0dXRZUcmD2sc2NgohoDqA72nznTqUNNYAAEEFZSxIUnApwJtUWmtpiQclIzolQldDlqG3yPgpbHBhok2JpsPRQzumXFCPxIqt3xA+vrcLBAGQqVsu9VdBSwKJHdroqmTqPLZfqAQ0GwKIRDBRhykUcjmQFNClRAQQUOMGdzcLW4cQkk26H6zPMzsHF3sBXehKVqyGnMaBCQOFPwjgURzV2jbhA7e1210ZR4FrAlVIYmkRMEMhIx+N6Hvo8gbiHIOqGhe0PBhDDGK5/kRrKDPi8EgHWmSC4ouBFYwJxhDCrl87dScTk7Ep6IbqGqZ/jnFsgcz0p2qtIBBViJZQLGNZJL5E2hnoUNSYUk6wMnYygv0jlwM4y5v1njzgmAsAoVAbfO5gTIOI+wITJoPXn12QqaHJqSeZVOzQmOEpAPeL5WKEmAF/VJCchM+oXWStA4/Z36F/RfoSeatNGVVNHAUDPOYf0eRUhTVJGchOatMRqgz11L3sZRZqWQdikqgPLlO3gd6f0f1MK/a2vxARpeU8V7DgFQySd7wiSKpa5+C9HQdddaJIx9c/kzMn4Tc58+BocHG2nf2xr7htgpYoPeyziRg3tKoIlCXtE+aOwqgJL3iwT6fR8NUjdSE/CDAkhyeCr6VhmQSnxemhhGc8Wdo9Id0iCPcvdjPfahBE082Y9bf16sxwWwuuL9hkqwAmblc37ORoUFdJ00XNGmhjILy0x6yuaW551J/jpLiuajhlsbVk243a/O57mbdSpwJDmWUTHGkXe8p8+fEPgp2DIl5fKn4mJpaLqPEMwp2j3vTBNPBmx2wHkDguk9Eo1jfYER48VF1Co1RUmNLhrH802UDHAno+4i/ZzSzCAhBPUpPWUU8L7YE8jDWpYpAyXhdMmU0bije4NFAwTmkDEDiMGeSNBYLTJRimn0JKaTgds80zzhr1NxiLbhzu5JWzhjmhXt9JG8OMa8Sqo2Ek6Zlah5oLqd9X/fd5EkUKJ5Ys0GxlnyGJORcUo9YwIvWjm7yIoo3MaKhKUlBDITFxklG7DIW94ZyNA4jkNc+u+N7pZ5Van6z98mHp0nmz9euG3um2B9tAAAgAElEQVTD9Dh0+LCKJzAjuTYxQksl6bsrsd/c1NlcrtCIRrqF/c0ZL8GQElIY4MWem/Nxn625FturlG2op9uOHhqXLBpJbAW/ifUt28lkra9/0MZHxywLe3G7JDR4GMVS/EIOheelIkEyceQcunHrlq2srGlPIKFCdsYbq+4PQJPHgR8wSr2vRCx2+NC49Og31tdUFETCinYWZwmfhVQFr6UIR4NBTfhczm7cuCUmpwzDZaaaGlj4WaTGRciurW+SCG3a4OCQ9lq+KJTrWiyjmAV5UL4nfWchM0maWBdVa8232NbKkj129ozl6jtWq1Ssb2DA2nsGbGlr21q7eqyMVwLMsZwbJkvzGq8V0Jm7uwJoTJ44butbG/baz38hxO4AniDLK4rjaD6xr7qcJoW6ViVtSD1RjeEso0jua9obZydPnVDihy49jS2MYfEycR8a16tmDjMOwcKloMGcDfQwrwOkwH714gvftPMfnLebU7dV5JDZMU3ratXOnpy0nk7kiDABrdi3XnjR3nn3Pfv48uXUPMiqacV9CMTQ2mqFtnabW1wQChYtemcQsid4cx5mBPrd8mArIMXS5QWbcknNBmd4FlSowfja4z2f5+yNlQrjYFZTQ97leBaWlvUsnFWxJgSpziTAEYodQMN6wx4pDe7vpReeVsNoY6NkZ889YK+/+batb5WthIltT4eQ6T1d3dImX1qYVxFKbJjQI69W7Xt/9pKARjevX7fHHn1Yz5A9kHFlrJFMc1mnioqGK6urQspiPE4+wZxh73f9a5djUEOgr88uXPjUhkf7bHBgyJaWF5XkE0c8/9xzkuJhHeP78fjjX7G//8cfSw/+u9/9jv3LT/7Ntrer9rXnnrGdes1+8pOf2lcee8Seee557U1T09P2yqs/s7XVdR9HSaa4KbZynyS/JlAG4BPMT/cAJpiKggcPDNiL3/mmrS8vaf+isEmQlc0VbIf9IZ9To5MFrDgXY9fNLVtb3xC7YWz0gO4RNHIreuppz+XsQvsemdl33n3fDuET1toq8BM/cwlYj6vcFwJQTtkGB/oajU2KvXwm0mqwRGBoeOxsAnQRI9MQhslBPIU32/DgoPxueNZf/epXhfqcm70jMBpIdmIi9xjz2BKwgs6qxLR2Ob+6tXd0qhkQwAU+lzVHzKGCvXwP/NwN6ULYcZw9zFPGgSYV76+YpO6NGAcxuewlr2PMKMQLbAdTEY8D5qSaGSZJtAwsXYqzgv0DFGm1Dy9+aBSAyL3YJoi72ONBi5NbUjiamDhoTz39tNbcG2+8oT1G/kS7rjCAxB57Cmwc91ZAcosGdYfQ4uSIwYKRJCdo9O1tNYjZV2Bxu28Ue3GbTUwc1n2ruJ/8zuJsEyMBiWAx3nIe6dMUrVYbniKcD1w//k2cU1F0VTx8F3jDwUw0sZAsvnnjhs54rrF/YEASm6gpsKcoNlaMvm+sTZPE5SvRid+27WpZrxVAitiNfAFEeDrvo+ga7Mk4+wMMk0I3911MviaMb0i6CgzGOkzSYAJOSErKPRB4Leco8tKnT5+xhfk5u43UU2vBjh8/bqsra2IcUkvgnNvc2rSx0RH7+NJHmmNnzpxSLeHq5Sv2ox++YO25si3NTll/F0bZOf3u8NiQFVtzdvny5zY0OGqHj52yC+/8xnr7e+3AoQn78NIl6+7tsYHhYauTy+/W7PDxU1bZ3rF33zlv+SJNJOZf1nbqZvnWdgmRrm+WFMvs0jTq77ZqacPaW3NWr7pvYntrhzwqPr1+0xZWt4zIoA3Jo+1qkjFt0Xqv7FQ0z6vyEur2GC3FnNEMYpwVDyKVtA0LlTmZTWoayB97xTZYPoy5iqtqVFR1PrEGN8sleeAw9qQh/KdnT0xRyCtvdLPtPc1xNSsEUMM8vKL79hg3xZi1PSvkAAy2a49ry2eto60og2GBzwBE4kNKUyelPYRVAvdp065ZN00imqbdHdqnkRafnZvT/WTzBVtd3zKyGNSo3LPJxYabv5prI5FveCHbX9kM+LznV/XP5tc1//ve1/6+pkLk0f56z7WicM/gBYu8WYjp3ve+u0C/nzfF6/bBV6khkPzu7nc/WpcNsNbdo9XcjGlucvxHTZrm94yx9RqQy1mH2oDLETvAkS/2ei6F3LWdGJUmeGoQC2yYmBCJQNFgRUTNav+6mhsVd3tjNI+BP/L9ekPUnJpZFrFXu+Sy1904k5nj5B0wPiNHoJHK+UcO88ADDwiUI8nyTlhIePvOKT7nOon5OU8AHND4p/6HRCN7P+c46/BLRsXvm7Fffv+PdgQm29DRhGWwoQCf5BTUCUEKRXOCDeSN3JyqYn0YFhWKom7TwWMDgV7L77I4QSFIr17IqLr8FuiQs0AJ3oR8qO/ZkYkJdQuhsBPktWQofLi/AgUaEEvQnsKfwIvTboQZPg8x6CQ4JEthXqrEgaB/bV3+BCTrsB6AOx04dFBB+cztO43giYCRpomM+pAlqteUACG7JCmTVEwiABobGXV942SwTNCL1ASHNc0DCjqz83Mu/4GsU4sbobHx8B8bqApR22Ulbh4kupYmJuWiU1Kko0vc0iI9bQoDwtpm9rQRg9QRImlzK5kz1kVp9ZAgIX0lN+KarSomJ4kNoWhSZzq6vryXY45d4kf037QR+/d/9ys6zftFU0ci6j0VaED57hd9XB4VYlKQUO8pWFYSlTwBnH66L2kThe9mIyS9r1CwrpUbRrYh28B1EDTJnHaHZFYXo3uH4gyCCXQX48rzoqjLnOUAoPEV2rA6+Cg+1Hdtp7LjRXXQvulzQUDB7tmpgUjygiAoJRBXHDSuke1jGU00BTHJ7sOlcfxA5HXxLOJeJRejQoUX6x2l5gVNFfATsjwKk1EEVKLbaBh4QbNxAKdmUzQrovkoBkfSwZV0W63qnhgkFLpON2WLJhHoY64ZNKTQzwmlz5oMVozLG/lciAPcfTeEk9I4U8SQCZ/0PvelepCoAMHFdbNWKDbABeCZctjzPYJsCjYEqSAOQ7PYG0FegGb8eDa9vd2uTZ+Q9G6Q7CwSFWVTRVAarOw5yfSaOcJ9U6gOuYGGf4MasjTjAlHvc97RaJ5ci6JJQpKMgDUdItBPng4UgR0tseHG0Ike7waU3oyLZJLkmLFi/2VsVHwX2ih0T0ES5ZX4ssfy+cxZ6RHLH4HC9p7rmNdp4IDsLDljI1FOQQSybwergWTZpV725xXPk2cruZBkcBpmY858a4TRer7opIPc4/e8OedjJSmDZIbZLH3GM5PcQJovKiSnIqLPp5Af8qaCmFlJziGaKI6MdlRqrIe7fD08xnR2gwCX3uzhs4INFujMeK6BRvdA2s817/v4Gg6UjCMESdqKKry5ZIM3XZR8JUNpee9ovibz64ZnBoWuPSHVeJ9g3Owm2YMw5lQjOklIyUovNQS4PqdI7zMaYg9iUTSjgSLQ5ne4vyheRyEEZJJ7jtTFNpxGO1kyaPsSLGIXpiam/CvCSyLJsgSLzxkYvp9FE1P7l4oVJIYUF7zJKZnD1Nzj3pjH0cDOZbyJg647Mj6wH5F+4nOQZTl+9KiQwezDFHzKVdhvGGmmQlCprGfD83KfAzwQSgI9gMzuKGZtp1Sxsf5uOz5xSPf64UeXrFSr29p21bJtHTL6RSqQu+FM2MYoXqardRVEMVBmDwApLj8bGjHFolC2FEV4LUwAGhVafy00YjGodWR1metFumS3KkNfvDYAguDpEAVlCk5HjxwVogwJSW+m5WUG/NDDD6vYF3IwIB0pYIJKZCB1PUlajILbOIUxjRMSQawBRziqWJ+S9ji3KTIQt7BkuEfiEVhWtluxemndRnu77OTkYSutb1hbZ5ddn5m3s1/5qt2cmVORXsUjFaXT2UFhMF+0jbU17fGco21dnXbp8ieSd8AXAN1hmpzh1cQYcPawt4TsCM3Xhq+TWDrO7GVuERNwX+y1zK/NzW3NQe7PUaMuj6dGqsA4ngCzxnSWyQvHUaZf/9rz9uGHF+32zKzQy+yRFFFq1Yo9fO60bW+uW4ECXaUsL6zxg4fs5Z/+VPO+WtlxAE3Nm7qMBQXSlfV10fZVrFHD3VlhXA+NecAeXHt3Z5uYCjTp8X9QwxDGXvK2oDhILCpmUSsSA66trz1HHkou50iR/tr1m5YvtkqaK19oUxzGnBLKObNnxXyLUMS93R1W3d62yYOD9idffcRe/8Vb1kcjrNBqRCX1bE7SaLAyWMujQ8O2vbkpWTYBCtrb/T5ai5J8eviRh+z9d99ToYk9jvNLPhUwJcvua0VjSoaqibFVR699ddXlJUEmCh3trE8Kux6reMwBmxEwFGPAPnLu7GmbmDgko+JXf/YLsSdoWL373gf2wre+qfG+ceOmXb92w1789rdtbn7e3vz12/aNb37NHnz0EUm4/uM//VhG7Gp+VNnbWxsGnKwProt7UEO4nhG7CKmWYsGf5dGJA0JAylNOZwGoZ5fhosi7s0fj0M9Il7rxQtn09G35SjBnvJBPrLqtNSwG6raPl0vKVezIkSM6U2kwMB6Mo9iBMnF1BjNnO9ehIk+R/KpPjQXMoyVJKQ8F5Ex9PTAfDh86pMYT+6QKjAkMQMHvueefV0F3YWFOwKRoJDAXYONwN1wD0k2Mn0sG6sBREZH3PTA+brOzsx6nw9rADD01IF2mhqam68ZLsjKxZCmSOnDAY1I9B6RwxWorCCTBnCBOQ9aGJqbyBpr/NNEUR+/qjN6VLIizX9lfMF8n76IZqv2m4N5oir1oUKEVvr0lBvxzzz+nZwS75dbNm9ofORdgwkgSmHyStU2DFzZXER8+jw20ZydWCeNPXEyO4h4ZS43mPj8DkY+cLQVYcnXOf8WXSTJRLEoBsnq07lAHAD3OXnLkyFGNsfyNJNPIfYaKved3jVwhFeGYH+S609NTWmPMn7ExJAh3bGFxUWsx5PNc/sy922DsSYIQMGK5bBVYoEl2lteLqeKVQ2/OEesl78I4Z9IFNfTvazusEXJGrzcwD0O2yNn3HvN5jOWgKWIC5iEsEGJxmlVnTp2x2dk7NnPntmR/jh87JklVzOupebh3SMlGR0bs0qWPdL6eOnXSMnt1u/LJZ/Y3P3zBOoo7tnxnyob6AAHsaZ32DnRZX3+3Xb78mXV19tnk8TP2zq/fsPHDYzY6MWnvv/OeAAQDw4O2Uy7b1samDY+OWzbXZr9974J19fSTGcnwfg3zaM6+2p72M+bCYH+fPf/sk9bdUbTZ6Ru2Mj+ndT7UP2y59na7/MV1W14vWT2bt51dzsLwaXSDcRmmZzO2vel+KDwX5ZUhIQyboQxLK/nI0LxPMqmsK/YSAUZhZ6YcRCAaSTbHnlWTvBRnOPuI2M0KCB18IzZ4Am8g90e8wzoXsx9GxOqa+5mkGgSNXBr04bVHjgSIoJDL2NjIYPIx43fzmo+kRGr+kuuw/6R8gfnRpnjZvQ2Rf6LAKyWLPQyKy7ayui5FhO2qSz6lW/Jp2PT/yG6CDa88uiGlejeis7lAH3lP8zq79+f+3vsNjd/5d2oKeN0gJTFprNSASFfa+L17mo9R62k0AJp8N+69vshrJFnXMP+Od97/0/dDB3M2agpNud699xCNkvvdZ4xN82s0fZI3ithbiSWjnFyS6Z7rOIuZBq4ze9gLWP/UgfSVmhxRyYpr/cONimamxd1/13VJzns/B2yAgZs8S5zplhcgg7UWn8u9APARQCkxr7lv4ouzZ8/YzPRtrW9yaOT+HOSVTdJsSAhuqz5JUxjws9QWkCDfWPd65ZfST787Wb/8zh/3CBxubddip4snDTXJLLUpCAMxI3OrhHgh4ZPcBMHOzo6kffgCYUNRjEIdQSEo9X20K4EeB0XN5hfmdYgeGj+oggMHmC9isw5oyFUSD0eWgThzI+mEyleQGaZGLgvCIScE415dNHdRP3cxTFwxgptadUeBNoHi1O1pY9s6mUweoYapeN8CVb5Fup50+EnYOZRBQHx+5YpvNAnhSADIvapYK6mlnGiioG9INg4ePiT0F5/PocrGRBDLjtbT3SPjPTZ+THDokkpHL0nAsCkhMSAJJ7Q+QdwVC/bZ559rjGWg2NFp3Z1doq+CjPCuuhfB3PQ59NjZzJx6DSqEAN0pcCTAvnlTROHr3oMoWABKSESpu/+Xb/JefQ+0vDrbLY7c49lK4isZsuI1whwbGBz0oN8rsw2qMfcbDAOuIZKOkKvhfUgIuS++F3Rvvh/NijDKU4OMIqZ0g1uVZDEOSHpRwOGA4HlL/gEJqK2SDjmeEWO+WXJtcz6rtxu5rbwHXRQ0SYyEfC0L8STkdUrqSEpoRDH3VYDCCK2BBvDDXAVbIRw9USDZ9Tq2G8eFREswI7QmU8NiX0fWqbxil6RCrg70e8y/omEQD1HrLZk/Cfm+u2sHRkbFBCGY5fVRyAomQxTZlXCCTtirq7AgyrbMMEGeu7EZhSWakrqfZGIcrIpGQAMasKdLBUMSRVCGJGtCC2PuvO6soRgbkG40FJyd5c0/CmZC0yU0hSO9fZ47vdPRXt50q0lSYV+WYF8Si2tSUTuxJpgnJKUk1FxLBDLBChDrg7VWRl4hPcMIwlOSRGOE4N5NiF0yi++RbLspl6NwQGbC8qH4QMGGAowjRdJ6Swwlxg9kRXifBHtITAo1ZL0YFY0rLx47CyXui+ANBhFrgsYzRQ/t0Ulbm98hcaCII+3osks3yVMk+Upo9oM+RDagypi5XA1fPhbelGX9hHwANGpnl3ijQkj9BkrHm6esc95FDTExV5xt5fMQeRtHcMd+o8ZWQg5zDkUDM4JreUGgnU9jSwUtLyyIrZTQfCHv4lqiHr5KZ1wNjv0/vVCfGopoTWdhh7lhvPag1BCI5qOktzC4VTG8oIasnnf4vFCMFRoyL/iW9rjExgpJJxoVQoLW/exzxKHr5ssAUa07CjdOVQ8av/RbkVGTVIZrCDugDETRPoU5kF+8Jp6J1nYqxKjgkJ6D318q8CTJKT2jNE8b8k7xO4kVE41NPos1E/tKzFGdOUmyASQcXxSpgo3h+79fP8huT1IoBNLQ71BRDiQjcxzWJcnzzMycHTs2qQAfaYCR0VFJhjBO7C8gkPcb/l544ZCKLVdN2GrZ2rNZGxvst3pl2yYnJuyTTz+3ueUV29ypW9WQeOgT8rKGNj5o0nxOTT+kfUIKhhigo7NLoIX+/gExu5CK5PsUkUuSYOjT2pdsWNnPajU4y15ccl3dunVzv5NHJO0CY5J4hwYHMQS/e+PmDU+6k3Qf4+GoapdWkIFtkmHhLKSRSXwjHwLtkV5FYs0TU3DGSoJMxd9dIWtpwNDEFVtMBSnO/RY32d5cFYuiPVu3wm7Fjh06aJ3IIVZ37eJnX9jRcw9ZPYuMTJuad1uYwCZZviJMF/bxJN3Cz1c21uzazZuSYxkYGrLrV29onyReY90wR0ZHxnRvaE+DNieO8kDDpUYBCzBvDk8ctscff1xzgHnxm7d+I6kbmTJHjCDfG5cwFEIvacrHOg1mGWPyzFNP2yeffGKzC3Py2pIETzZvLXs1OzQ6Zn2dHTY1fVMNBQAQ3/nTl+z99y/atWtfpGZiweWr9kwFEmQj5xYWLMMekIqFrqOfQBbSM2Q/oECTte9/789saoqG17JtrrlHBQ2HFs5OFZCcIeKyRG5+uo28mCTC8NLifGu1O7OLKmqyxkDwUuSBAca82d7esvZiTgX34YE+y2f3bKe0KhZEZ2e3vf76m9YzMCQZtM1KxbaqFevs7laxYO72HTt57JikYWMfIVZVYW5oQOuGeAETdTxAXPKP2NXBHWosJ88yrk37UIoLKMZL0jObbSDcKWoxj2n+Lcwvqvh888aUdbQXJHXDZy4tLdgP/vIv7ZVXkLzK2Pf//Pv2xdUv7Isvrqlg/fhXHrf//j/+UWvtv/5f/9V++cvX7f0PPrK//bsf2uLKqv37v7+aYhEeikvwcU2sV2JupJVY97Bk5PCBlBhFr+1N62yjubFjhRxyNQNibepsEggka/VMXSbnIH0PHz7s96r9Nicg2BJNm/Z2NRllTu0qjn5egd6v1RoeCsS3FFhpuFKMlcmqZCF39dr9ooozIBl49NuRBiO2WFlxNjlhOYwd4lpJJ/JZOWfwISdD84wchDVDLP39P/+effzRhza/MKf4mvyPr5CPRA6TeDs85DizYRKpGZ1YgMw71jH7I/JJzAX2KGdw4dlBTENVyA2C2e99D2M/ytk2SNI21/9mfDZghYJgre8JCEd8z+cjVcX32R9ozgqMUUezvqznxDoRUzLF0g4Cgs1U0BnO82Ff5d4BKhEPcQ3PPPuMfeUrX7E333jDPvzwQ+2jAtok6UearV64d28hngX5sMfMzkBkPpF3ixVeqzvjpMmLitfBquBe2O8arLgUi5APeEOjw0aGR2xmetrzg1pNDQ6B4vb2xBhgD/eYHdlNj7UjDorCLPOOBtvt6dvy8GBtUmzn5zS+eS/5qkjqOHmM1fdUN4BN5PJ7u1beQe7X89LmRgXrOJ5/GGmLlZN8N6LxwJ6vmEvNCpd7UnydPLxY/45k8FntaHjPpbgnGj/M7/Zim50+dcqmb0/b1PSUdfV02dGjR+Upcnvmjo0MDYvtSF7POvr000+0j544edyye3t25bI3KlpzFVu8M2VjQyNWLdfEqodN0dvXZZ99hlRLvx2cOGHvvvm6jY6P2sDomJh8zAeKjotzs9bfD6O5xXr7hu2371+09s4+MXo+u/KFrW2WLCNPIW9UKPbZ3bPHHzljL7zwNauW1qFa2qWPPpL0025Li82vrNudhSXLt3dbpUrcuCMmrgAMeMO1eKyZ2XMvivCh47kzH8OzLYBB/qyQnq0qnoz6DzlEsC6UDyRvIwEcqlWXtMVfzPYEIkHeSvuHAEXOcEkpqKSt2opZG4DVlDFbXFrW/FpYXlE+LaWFurPGE8RJTYy8SJgZ62pHQrhHeTl7HsABmk4lPCLJDzLIUiamW82lbz2uBRyRs8HhQbEwuL8bt6YTiMIZJXgeBTMhZWOeZ4ThfKpbBJs42CmNfKhJXjt+J/IIjVsjyYt33//zfj/T76YrilcGePG+79swot/P0QI0eNdab+QldxfceU3sSc2/d+/VNgO4guVwv8ZGY29p+rzm6/jdUfAx8npWGncx032/CSaFNwcCvEYTzSW6vRYGW9PVOwLEps9puoYAqe2P+T6jovmaPdf2a+K/Ro0sPefIpeJ3YszEMm8B9OgxgtdvPK53GWdkn8h/vdnK+QIojFgVcAa/Mzo6JhlIQJfsyQniqkY13k/sZ+yleNex5+k1XzYq7jelvvzeH/MInB0YFg2bAiuLisMNjXWKe9NTBP0djohNiEgKWgS+S4tLKsaxMfV19zQKPHT6kEziSwUcnTIuC0OwRGMAQ8zxA+O2lxZvpeIFYxasNNlTV9sT93LqRqI5TiDppqiBdnY0kKN3kAuQ/iGF6WxWKIqjk0cUMLLRFzDtbckIdbW1if74rhJHPpuGA0U8JJmguBIIEywS7HPYO5LA9ZoJnmZnZqX5Ozw0pMCNQry0j0Xt3BGChy82TTYoEDagUhkT/CdIlkJbkAIrdC5kWAhCS6A6RvGocGPmQKRSPCSQkgb32JiCUAUUuzsqRFLIki59MloNFHNoeXqCdHfrofnf9x56wZYIuRwlSvdhWNzVzU+GyxTr2DgZX9BygUyPgFL3RaCuAq3rwktvNjVfAqHrxWc3QtLBInNPl2vh/mJsXP/Pi6QKghP6g8IrRY7hkSEVaShuEbhDPwbZyjWuJvQZ4zg84vRfihCSDkMGra9fQZeM2kg4kLZJMl8ETyqcY7pIwb8JRR9NFqHx03zQeFOJSI2KkOaJ5IGf6z5oGiTkpxcevUAYxVE1NZJGrw5zodC9cx9BgI/ZPiNGRU0V6JAschTS6Mio5hmFFSy4GE8+n2LOyvKqP5vwC0goND6aOeVUTC/kegyQ2jkJaRBSFmE8rCQefcmUlPE7FPhCbiSaaLw318D7Yl7LF7dFwcnZOR4AeyLtXg4uXeFyc0I4ylgUySpPxFgfkktq8imIaybBBskXzTxJLiWEq9D1eJNUq6KRM0c2NmhSugRPBB7RRGUoKKbyHNc3thQYax+rUkByA1an80PhdLkCzedEdaYRJu30JNuAL83G5ob8aSSTkQIcBWjJ9NuDHZee4jWSCEoyR7wGGSGxSVKQJWSvjAh9vTmSzD0kGIPw13BEjY9fIEIiaFYQltgFHtR641NrtQ59HEkWlxFzJg1sDpcJiD082Bzu3eIhmCMYvQij+Z6u05Gmrs+vRL9J+ul+nC/GKRgO3mhmfTg6OrwsuDJH6e0bqgXrgf2LecgYxWfzHl7wcWkWNe407sEGc3qv6OXFohqAKta3kQBvCqEpxLoYFbyPF4u1B8ho3s3nYQEKIZmaByRc/FzFO8YgGay6EbSjksNbxk3LGX9vVDl60veHQIJxzTHGMc7BJuFnanylBhG/783WfS8VrjP26gYDJhUueD/umfnNvIiGH9+LhkgUGYKR5cXv3Yb5OHusN8lcGo7nx14Kwo71T5N5eWVZc504gkI6Rfyx0VHFGJxzNMlbVSh0GYO29g5Ro0lOkZSRFKFYNHhhMEa7tkuBbq9ukwdHLbNbs/HRUbv0yac2v7pmWxg4ZgvW2dPnRpWVsi0g00hBSnKRPXby5HG7eXNKsjUk0cQZgBdAmV65ckV7AMk81wjLEpaT5A6S9JmQ/dHcosmyu2MHD45LXhJ6N2ao7W2dKtSePXdO43Pj+nXFP8483bNjR49qvfMzzlaK2V7kTOwf9GzRnO/o0JiyL1J0I34JTxb2A4przDmxe6QlXdG/WfNoSQdDh0L29vqK9bZm7eTEuJXXVu3g2AHbrOzYhctXbKlUk5l2H8VWpH5KJRWEnnn6aTEpKqWy2KyO9s3Y2saG3eacm8oAACAASURBVLpz2+bml2xoZETGp8h4wRbBz4LCCkUQztwG0EFGrS26X8aCucO4/tmfvWTnHjinve3G9Zv2q1+9bpWyy1ZxvtOoxf+BtcP9BYOE+FR7nnnRs6e7S8/wwXMP2K9//aZVd6vW3d+rtdrT2SkPjENjByQBtbw4b4OD/XZz6rqdPn3aDh08bP/6b69ZseDmpCp2CziyK3DNBs/K26hCg/IUmYs0WtRgaiF27LNKaVs+FQdGh+SFhEeAEl9Qe0jPlb0RreJBko6UiTaF8tZW6e3TnKDYm2nJ241bU0YdSShSDLwT2nW7tGXFQtYKLbB3izKG7u3K28522R559DH7xS/ftNWNbcvDlsCPbntbDZeJw4dt6tZN62xtk2Ev/h2cxexhfX29duvGDcXKMLVJpgESscc4k5VCtsexrGl+3+flvswZex8yV+Qq7NmBmNVzS81wnUcCGbhP1Fcefdh+9urr9sKLz0kf/fInH9ns7Lx997vfVePvV2+8b9//3gtCvf/il2/bD/7quzY+ftD+4e//3u7ML1qhrUPXw/na2YF3QsmBS3pKLr0BwEOeY/Lm8QYjhTokwOqwAJA6g6Fbc7T5wvySdLS1L+WIDfgvZydOnmj4PElayvaUk2GczN7isWhBwI54zhQdiVtCDm19fVN7I8ULQAfO0vDiDGAx/Bb6+np0NgcjGdY6a4r9U2wVfFC6OhUz0yBBYqWDnI8KoerBeyrEE9cjGclR9uyzTwmsxV46PDikRgDPmNhH8XliJ/En48Q8pDkXzdlguoYkm4rNiWHi8Yc3zHnWMqpOOvmcGcjUKN+iIb256a+hqL3rYCVywTrdOMPEtCami+49yT2y5gT4oOEoeQ68RNrkYaj1uucFMtaPCrkpt4Ktx37FXsq5+vAjD9vXn3/ezp+/YBcvnFeDN3Iz2E48y2rZ/SGIN2HDS1s8yZoKFZuAbZy/NIECra3rqtd1vrmP2Lrnp5Kb8kIya4eYnfdBxnNxYV6ACfJFil9zs7Pyb+SeGK/INyKe9DgGU3gvEvP3oaFBgeucUbaruUXjZ2VtzVnJEbsIMOVxAnOD58J/zGuayZKgTY0K8i79l1hY7IEyZU9G2JG73FXcbIoNmW9ifws0lWSrkqxslHPFmJOUXN0Z8appdAt4AMDhzuysnunTTz9hd+7M2a2paevr6VEjFW9CwIjXb1zTpz70yINWr1Ts808u24/++gUb7W+1xbkZ6yi0WWkTJuK2tXYUrLUtb599+rmNjR600eFx+81bb9ihyYPWPzBs80uLGhsaurdv3rKezi7r6O617t4hO3/xE7SebC+TVcEcj4qWfNFK5YrtkM8ga5ZvsdGhPjt0YNj+5MnHrSPJBM7fmbcb0zN2+ep1267Vbauya8XWTrE5GdAYV5jyLoPkz5j5Ko+gNqQKPR8RsIYzPhkyO7vKJbwawLGUW3pD2T0ggpmjWgM5CR4iifFCnOJSzw4+hfGgWFr+jMIEWEc2I4aqfPJ6esRQpeEA4wzmmcfaiTnOeKQcAz8gpKRQ86AuQjNVc3oXo/KqcvTyDj4XxK3OUNc6TqoDXCdy3IBIpmfmXGpW7B5nH94vpxCgISlg+Dx1pojnRPsNiEaRvZER/e5fYn57Dnp/OGi8Jpo7PnqcMX7+BLO+8e73XHS8a7x/XFfUlJoL7pGLxXv9vjpRFOs9d/I8PL6i8Rigp+Zx+EN1puaxuOsNo+HSlDuoVtbq4CcHaXl9TPO3DOiP87YgyW/JLSVACtekxmzyMoqamEd53jzYfxb+76gx8VkxZnEfwVT3e/Qc996mjoDC0WhNEsjybFQdx4EkyoVD/jaTEfCK32PtUovkecMSF3sX36hiQTEUMTrnIE0MAMwbgFBy+HYVvmxU/IF19+WP/khH4CDGn2YK8qLIWcwXxASgQEbyxyGvzb9clrQBC2l5aVnBCKsUajqBK0EiHWqSTn2lRCSb81I2UlLSem/vEFKdJIozSIFFzs262OzmoW+D9h4dUzEb1AMbC+aKBPszt2eU7HOQIrnABtHX3yu9NjUW8gVR5LvaOxV00FhYXl219dKmHT1BMeGWJGYwXWID4j0HB/od+ZPLu/5pdceWV5cTvdzRIBRN2CTQIJceXnu7ZIXQegcNBK0SxKA05kj+UqGbAmdISLGhMo6MEQe5CqvVqg0MDEhWi8SIjayjC8TejtgZJBG8BtQaGyPURZKUKEbwrNCQ5pq16SaZHad2+kEqJG36e8C2m8DbCRWTWg6heRgQLic/7B/eTQ2Lu5sUfnDzPCnUMD/YTCl2kDAQiICYJ8+TbJKCYtcrjQogQUX8k3vleXL9QnkmrT+CaTZtCjLSAGSDxmgwoT8oBlHU4RpomrHpU8Bjzhw9csQZN0IcZtzQL6FZuSbm4OY2XhPIhLRqzAkI3EeEA9JNY1WAk444TQvXYmf8vUDrzAtnA2GqSrDnKGwOJfeFcPmcuDdPdJO2e0Lrc78qFiedeTUslACAkPTkNwqD9wZHJLZeANmnZVJA1aGbUPDybpEutRtU7dYdsURhiPuEjuuat55s6vOVmBMAuI9MNLcCcbCfaCSwbqDu02Eujdqsy1j5vMwqoRL6KwUm0ZwimQcLI4o/tGKKEkJpO1JRDUhJETjSnaRHxU+KPDsgDvoUvKANrNowEjxJMzWukx+oMLW3ZyT6Koqm+3PJGH8v5hCfG/MxvA/kwZJkjdyA0eW5ouCtZBz0ZZqret6JISK2QmKC8fcI8EKyiKILa4mCAfNMMmWp4K/io5BjHsTzRUGT9SW/hR1vYqac3OdRQrKzz/B8hcpPpvVKqmWwzvp1Twgl86khKJmBhKrXs5ZMiQer7EXsvaw75ioIRenbJ4SiGk4NJoWj79xk2xGMPg88CVCjAl+DJCcQxWqfZ65Xqn2h5g3JZh+W5iNYzCd5ZyCP4FJZ2kOSdBbziL+7HIo3P4I9xLiQcJOE+vrya4s1JjR2kpHgd6Ih7D93nwsCRhqA8sCAjq5EyBtQMkAWPR9EcdKmlzePJ3sY05J8lZN8gSQNxLzw+1DhIiEK+UzmiEup7SqA5V44j8RMSD5MvIc3nn3XD6kr/u5z1enF4ZfiZvIuSRJa4eHx4g1ibyQ4O4y54Q0mnnOgRKMxFvtUJDn86QU/Z5g4u8J9Zvx6nNXCz2NsdY+wA7NZO3JkUmwFzs+DBw/obEH7Hf8Kzk/QRVCr2WdARfp1IwPEGZoXewMUJfJ/aFVTYEN3e6ivx0rLa3by6LgdHB2y7c0tm1tYstvzi7ZW2bFatmD9QyPuWbCx4T4QwwO2tLKi701MHraZmVkhomBwgIo+eOiQYfx89crVhBTkOipiVCAFwnyXTFsydBYAQ4bKyMNs27GjRxSLId3B2sbsFaQYqNliW6vAJC2gGBPr5OSJE7a2guwL7ABvKAXrhrH1a+vWvkl8IXYPhQQlY9HYBt3ubAv2PY+z/KxREwtjynS27dWqVsxlLCc2xQHbXl22wb4Baym22tsffGjbe1lbWMMotigvhnwhp6b+U0981Xo6u62Qzdnt6WmtrV4KuStLGk8MtScmjwjQQSLGnggifWRkVMU3sYyQTNpBhx2kcpKRSEhQ5s7Q8FBik7qpPXOIJRfzkYkHsloSmam4zwqZmJzQ80DCiLPB9Y4z9v3vfs9e+/nPrVzdtuGxYc0bri2zu2dFZElpCEvnAm+APc3Fxx97XEjba9duKMHGIJqYFcmmNcyJKQ5pv3OIKtFQsMzgUuWzGTs6OWn1WsXWV1btxPEjSkiRhpF5uuSf3JOH16vYIjBPkpLSxpeQh1mYdlXJ4tyanrGt8o4YFRX0vRP4g0L1TrUsLXBkMnKZmj375CN2e2pabIyBwVF7/+JHKorV2NfYBzJmB0ZG1Fwol0pq5Hd0derMY68Dmc1+hjQBZ7Kf+QUVXHVm4TWF2XJHu928NW39/b16xjLNMhgyFcsX3BuH9cz8QTKRPZY9zVm2SI32OUhAe3qL/elLL9qH58/L/+748aM2fvCA/c//+WNJvpw7d8b++V/+zY4fOyoTd57xx598KpkcZLv+8cf/bMur6wlM43lBIV8UC6r5vNcepfXqsk6NAocKcWqnJP+QnBpNzIHFxWWNLZU6cg0KqfjucD/cC8Vr9ixiF2JV4s5Dhw6pcAFIiUIMcnW9Pb2SvCOGZb/2saiooA1CeXXNZcX4QjpJjXviWljoCbTBzyh2S/+9rd0Z7sjwipXYovMEaRV08rUXwNgptqoBKm+fclnz8KEHH1RDihhFTAjOs4Z3gZ/D+g+vhuqu5j/rhz2wuoMXFPrd3Lf7LZCLEeNxFiMdxfUrpk0NDAfs1OXDokJrkSZq8tRKprhqMHV2JqYQZznnjoMSYh9T/pHM2ZUtZVoEZCKXcxAUuXCXJAAp2lP4pnnJsPIeNHnxpGH+njxx0p588kkxN9566zc6P9k/quWKAGgur+OMXT6TuJcYl7hEkq+ZjD6b2EneBEmGVSyDTMbGxsbUBCKP5rlEQ0dMwcRk5355Dxq88iXarWkfJPdhfBl3mbUmD65gHkR8o7M4gaWYX5yzXC+NdeJfWMcY0bNdiYWaYhieB3tPo1GBlCPyxKWt+zYqeD3zibiB8wUGD3su9y1WaEhTkYum3IHfafYn5FrFTE9FxQCksH/GfTEe7Ds0yk8cOyFG2sydWRlMw7ZDOm15aUX7EGc25wCN4C+uXdWZdfbsWVtZnLfZqZv21z/8tvV15yyLG0Qmb/NTMyqqM/dy+YwkhTvbuu3g+KRduPCuDQz02YHJSXvt1Z/bgw8+IHblzWvXlFe2tXfZwMi4vfX2+9be3W97LVkxuOYXVqC3SRZQgE2YsbVdGx7sNdspq2FxYHjARg8etKzlbX1ry9585z1b3ti2XWMvJob0WFJFVTBxezUBKLOGfAy+Rt4kZD4IgJBkEllzXidwIE4UkDWekukiF3KmOXtxeO0xB5RjE+OXK2r6AAKgNgLoj9oLv0F+hhR4VU0DGk4Za9kx62wvar+BoZmR9CsA1xbFd2LOA7qQNxd9w2TPraZBzdrx9pKJtks6EfNxpvu9VV0Gqu6xpeTtyAnU/MFfBZAWJsaVJPsW8nv7OdW9Zb3I37w24Y2U6MJFfhDF7Hjt/UqDv69RcW8e3/hd5a+JmUQdRC1jr4vEV3N7xdeMf8X1NF/Xvdfm7ITmYv39rvru94pr3a8B+N567/ebf97Iu+95+7i2ez/V9yNATt5k8BzG997IWUNJg3wNeWPyEOpzzsx2EDM1Ma8x+D1GPhqs+gBZNgMvI/eIhkwA1SLnCtBcPMvmHDE+Q3KFSQafNeMeYh5TN+pDiaHDa0+cOGHXr11PYNGC9nlyOc4EaoZ+fuyIMU59Sx6sezAzaNqXlIt/yai4/9z98rt/xCNwrLNb6Es67E4FremAIeAA1aFgKh1mFIdZFEi/0NiAtk/xEIM/EHlhouc6+17MpBGhwv9OVZqv7a0cJo7OIUBnuyWgA7WG3jSUp9uzswpWhoeG1UQA/UTwSgA2ODRk1764pkYJhw7XyhefCX24q6fHkwNQvTKAG1Kh/IML5y0HlfPMKXX5r1295htWKpRCO+SwvX7jhgKWwxOH7IMPzivI4voIvNFxp2jI74AmAp0JO+Lq1S902IGgQ94K02Y696C4GFt+h849utpsVKC2QIGiiatCeN1RPLyOTQ9pGVBOjPPVq1f1HhzANJDQlQWhIx3rFIiTEBPgUUwm4FcRLQTj0ybtskDRbEgE33TGNQ5bP9bSbI7CoKOIvSDq1Orf6YA3AQIo1Kp7TdDa1a1x4rp0SCTPEhn2qqHhUi8ctiFVwu+Hoa0C8Sa0vpBkyZAN9onM+tKBFUUz0X+RjpFBMfMwIykKNMmhDDOvr127buMHxvReNKyEmMfcOI0P4QzxHsB9giEo76LT5nNK8jo6utQI8ebCngoNHiy3aK4zh4VopjhcrwsxQpDEZ3DosY4IlhSMpwqp6xO7pm/IGnkxz68hGCUqsKag4n4BUTAtFNQntoMK44HaTwgEPpsAE4kEGoAkoMX2vApZjiavqaAmGqxQCRTgHQXuhsd+TQpCEtV6/3r8thyp4EheIbJ5fskwndeS0JLkRYOJ+yU45TPScDgSNMlhaF5lSYbco0IMCBXLU4iWuhBerNmz/oF+FYuQWlHRVBI63nRhPcS8JgETQhyZDZnOOhvDm56OStW8pukGGpRkOTFnuMtIwgmOKTYwf3k/Zzl5kTQYEgpm0nW4vjUoUlBHoWG5/1pJCWGCOdhva+t4qbismlhJSS4l1jR9BcYFFL/vA16YiEDP9dfRzMwq8aa4AQKJ4EampTDGYJ4kZkUg82VimDSAhZoTKyt5PJCtJ/kjAijmC+udvYz9yAnXqfhMs05yRPtNi0axO8lm8bNo7mrsU3NFDZbQy0+FBTX+YDJEB3V/29L3AqWuNRDNRd2jF2V9HbnmdKDG+Az3WKlrnwCxGIidKEA1MzvC3C3uI9BVIIWlmZqeAcjgRmJAUxC5roSm4f3Qxo4GBNJPNAoJTrV/yeTPGRHcC2MvmSx5OkRRH7YOEhtVoQJZF+xPEYxzloaMVQT6UdRqDvhjv+FaKZbzPlyD/KfSc9RaTkglnw+OvhR7Kj2jSCiCAcZcjOeufalhtu1NIjGYmtaTGiHqhjXPczdVpNB96OAhoYbZb0eHh7U2MYKen53TvFNTKJu19vZWNSPwSeLnH126rFiFRt3nV67aoYMHGsbLKrDlMpa3mh0Y7LeJgwesvLklEMJHn96wHcwoMW3u6lFTAgQ72tb9Q/22sLAkFiaFJM705aUlmd0tLa2oUUHccOUKiGPXWWdMKQqCBpa6D/rkrTAQnRUA88rR5Zt27Jh7UVBo4txkjDlbjh07ru8jKxTFNtbXmdOnbK+2p6ImxUtez54gRmNay0oWkxmwQA14f3R2CK3O6+IaGd8wMI3vE8c5K8yb6LvIPmHsvLFqZ45MWGl1RTFeZ0+vvfHbd203V7CVje1903tp8VIkesQ2VtdsZ7tiDz3wgF269LH1DQ7Y3MKcJDpBuRNTUtzT0majq3sRX9T/8IqBFYIPBUVD4tGqM+c4q1nDFKokv2mmMQEVHz5Mu5I7TA1PCXs7BV/Alz6AKxRQXZuej6dR8eqrP7ON0oYdmhz3NUHBraVgk+MTdmdq2mAH79mOWdbZn2PDY3bgwEH76SuvaO8Us2cb2acOW1hedTm8JJ2mhiQa6wImoO2NdF6LHZ2csO6OVltamBPine8XkYMSS8KLfGJEe10qFaGcyUvy7qhxR9vxsDFznjh63F5+5edWrWesjPlpHrAA+wosDnbumrWBSt6p2pFDg3byxHH75OPP7NTps3bz9pytY2DK3JIxO4zgvJ0+ecounr8gRhHxAuuSe6EBgZwKxss0mxhjwE2Sj6xWbHh4xG7emlLTALmjaLAi6RHsUsaGc54mBoAC+TVRDGe/5jPa262joy1df0asgIlD42L3oDv/+q/esr/927+w29N37P33PrC/+sFfiZnz6eVPlQ9856WX7PyFi/bOO+ftb/7mBzpvX371NY0razWklxrS/kkOIgzp1agtunwdkVcUOUBOElvBvpbcotiajmJGzahRVGEfTchhscjUXKiLFUYsxv2wF8CWIdchZvpf7L3nc6XpeeZ34wAHOacG0Gh0nMgJHM6Q1EhMYqY4opbSakmppLVrXa7yfrD/Gle5XF57q+TybpW91K5WK3EZhqREShxqZsjJ0zk30I2c00Fw/a7ruQ9ON2dI+yOrBtKwu4GDc973eZ9whyuQH2W8nsUTrhfmMI1Kmhyrqxs6d6VTb0qE5qUa1ZL0wY8CJLalVHLv56XcC/HTh554PC5euKiGMONPPASCU/Y0xSfhoXNn49y5s1q3xNSW67FePWs2nzWFcszc8eGzL0bxcBJ7LmWpfI08XxeokPCztCESmnxPfm2SzsCwu9la3wVNS6CESa5k28qZZBZvu0ByzBnGj6JOSuOSAzgXsayiYlM8AnYpAG1rfl69erUeD1ZammJzi33VzRvGj9iVvOJTn/yU2PHf++73YmZ6Wk0mxnFubtF64hX28C3lEhT+kw3Nz4ZHhrVGBOgSk9L5IWuGJi2+F/ZRdFPZY+Gzmv84h5AEuX7tqu6H50heyecLHEYjqABUGLtsTNSBNQVBz947MjQsFQDYicSqxM48R/wQOTa09sT8tTQYP0c3nWYXc5iY11I8v8yo4Pnmvid2RGGaJMo7QUv11DIBPgIdHIFD5NXF2bxrdQcDkgwGIsc6PjGm2gYshpMnT8W1q1fUeCOO+PDTT4tNQV0C3wvmETULYoYrly+JtffUU0/E4txsLM5Pxx9//YuxtT4bXW3V6O0fjv1NS9XW9gBmHijv6+7oi+GRsbh4/s3o7O6IsckT8fNXXxOwoHdkNG5fuiTptP6B4ejsGYy//+nLMXZ8KpZWN+LgsCLZp6bmqqSRYFVwnq0uL8ZAb1dUm/aiu70a7S2wCdrizLlHo6d/IP7upy/FndnFiBbkdImT2nVeSQcfv4lDGtG1WF5Aw5790qju/EqWuYrMRSmAgQS9LTPubVhroNbb7PdXfCglKUvza4+aUXu00WhCPlYgvIjhoWGZBvNcYPOsbQIEs3SqvJWQckP2sw2ZVMezFTXI21X7YC/CZ4XPJ/6GYSHDce0FzilhVKiRiSRYJ/6dbTJOZ71Q/9kQMwVfPMBqnk2wrZQPFt9O7U81A5I8/96LT3FU98jGYa5BtW2SWZGg0JL3vl8B/v2aGO/3etUByrjrNSW/vo+MUa/vlOsvEl7KxBtemDG4xqBBgeH9ypi/rqmSOX7j7+fvZL2iMe53OOdrfK/7ve97xU/QMe79EsHaj3bT+8tG1cxJnqPinuK3Kk8kADulNpXKGwnQahwD17eSt+Pr5HqUp5TmHc89c8ijezliZeS9mTEI0NMqMAD5/Bzt/Wfwbq/qppxDnAcor5BDw4AjT4f1Q4xIsxlQAHkhAIaR0VHd66VLV6QCIolwvM9ogn8g/fR+U/mD7/+mjsC5nn4Vq1jkFFAlxdMMhbPPepYEgW2t0sZM9DE6oywk6Nt8wVpg32QBU/CXznxJACXhIKPsPaGBKIKSWBBA5QFDIXSgv1eFfnTmZu7dE6IFFEQG3RQISbilrVlpkXQBrz3YM42QzyQhW9tYj5npuWhvrURne0c88djj2hBu3b4dfRiBd2IiuBzbm9tCw3HNbADnzpwVJRS5BpoBGIjfuXNH104RwQEtxXfQ1yEUICiTUydPxVtvv62fd/f0luANPVeb6sL+4GCjA4rZGsisiYlxmfixkUryoFKJ/t6+GBoeVJAP+gb9TMZ/emZGCQQFZTZMng8UbjY4PjOLQATdMqQS1dJo9fxKFL26xvUD66i74IPhyNg5/83vI7fB7yhZL3T3+xoV5W3c4de27ebOLs0nzwsK77ApCHApHpMgoketILwUPdx5tp699EmFVHZxNQuKkmIRGskICa5DjI3OzlJYRvvcBpp0oq0RPiBGSkenJb7uzd5TEjI2ekxj7do278OBh8wZ14+huU2aFJhJagwkmZP5zq5uIZuMBqKY7cIwa2hq6oSeAUkiga+KzVvbugYGw7S+NgVqWYAViqV4jXCNBE7MNenOliBe/YyCKBB9Xma6KSfhtZcUxQw4WQ+JghZa3pAjox4yWCjsGMad+Iy4hf9UBBHrxWNq6aAjpAnyFHZH8VPnWvxzm4UKWV5Ml5N9wFQC+UnTLotLFMo4kF0UtRmkDnM1cUKol6RI8vYUaix1sCnkn4MHNO67TFkHKVOMI420qGgeGsFAwdQNJY1BQ3FbEjAqYDerOOGfY95J4csIoyMUEhT+spTKMnPQRxBOoRkDvx0hQZF9SFQjYwNK0DzhkLmbE8wjzwcV69XM8PWBIBUTaWVF78cYsqdqvZRAiHXCvyU7UczJuZ40sBRLqQRfzEXen4QXBBPjDAUcKT8+y8Uss0rYq5jLFEwJ9EncaPrypeatAjh78RAYqslKEa7o8Hv/8SB7jWB4yLpysfYIxWNmjQN/S6wxRkZzez/wZxp1mAwHIcVL8F6GtOxADmgzaWVu1tkFmNyXPUQ/b2BH+Dq5fwqBbtDnGs091E2wI9aN7rB4XbgZ6+ZrZ3eX9mkSYjW2inyiTX/Lsil7NLioLLgd7u/H5PFJIaaZr0YBWTchGz0qvpRmC9fLsyCJZA5PTp7Q/F1aWqwXnC3z4GYBz0sySoXhIhZkeeaMEWtQzcjCMOF3WG+pt52FH26BBh9zhHNY+0xZT5mciM3SwEQ5alqm9IOLUaLlqxnqNaZ1toXpsVlo2h8J7pmrbe1CR9OooMk5PnZM5zNNQaHq9+xHQDOBtce5SYGJeAYDZoqOkj6S1BExje+D/3a31mKgpy0GOjtjamIiFmbnpBP9yutvxfZhJQ5b26Otu1fvhRTRnTszOl/mlxbVpBgZHo6792Z17gCaWFxalkcWr8HvymbkVX0+16Gz5sBa3jT3mPNCLkuHfVtnDMW//oHeuHDhojSpOfcp4D791FOaRDRc5McidOuedLhJ7El20LtHOoh75Fnoc7o6YnV5VU1NUO+gfTkbKChQaFPDXo0Ma30zN4iTKO4QA9qfpSWOj48q3mLdLSwsxubaVjz/4Ucln9XSVImh0dF459KVmF/djHWa0e1tda8V5sHo6EisLa3EQ2fPRRfG1PjiIO/TbrDI+tZmDA2NSE5IYBk8NHr6tC8hpcazRyJTMnnsFWVcKXxbTmgnnn/+t+L555/XHn7l0uX44Y/+LqrVNu0/kqGT8ar9UvhKxpkb5XhDtNXlWfj3l77w5fjRj34U88sLMTqOZA6yIvtxuHcY506ek/TTzRvXo72zJVrbK5JZ3N89jM98+tPx+ltvxcWLVxVLU5iDGbcEg88bMRIYxwAAIABJREFUiIo29nUz4hmNcWK9rvZqTB4fl5zQgdDszWpUYLIO0xgJNNDtzAXAMTQMuA8KixTvGYuh4REh7mD7sLbWN/EJaYorN2/H6sZuVFo7Y2kFrfVO+0GhTd4S0UW803QQLYc78elPfTKuXb8ZN25Mx4nTp2MH+Z5qW9y5dzfaOrti9t69GB0ajsH+/lhYXoqtYqbNc2DsTp88qX3w7vSM1jpso+MTE3H50tV4/PFHYmlpRcCo7t7uqESzJVSRdKy2SB5SLLQmI7ZlmExirmKTYyfWAEwi5ktz5VAGtBV8rVqr8ZUvfzH+6j9+O86cOx4f//jH4rXXXldsf+7cw2I7/eVffjvOnp2Mz3zmM/EfvvWf46knPxQPP/pIXL56Lf72299z41B7MY2clB90vEt8Jvm7wkqzZKmDg/o8UrzC+HofVXFic1NxMXlCNp1VnFWsgUcdZu1bir+QiGIvfP63Ph4Dvb0quAvk09Is1DDxNGNMcRlw0CuvviLUO2sL4/eUraVgC4PMhW6K3Gba8B/NPGTjeC3I8JT4Zf+8fOVqPPfcR+KNN96K7k7fC8wSYjPmC9fLdVPsay4FNOTDYDtkFpLAFcWKrp/f/6UmW0WIazevHcsRw4gVUWQuiX0TdME1sj+xp1KoIV7nHOQ1xOjEK443KLgiB4fEsKUWmZfsk+zF7LUAx4jFkM5l/9bnIXO3vRtz8wuWsir7hs5/eScZKCfGO2ewDM9ht7TH7/3eVySV9OL3vy+g3anTp8VmIu7N8WctLi0v6fXswTRbaGgxn8kfiBvTx4J4BI8D4kCKVQkGUAEu/Y1QP+jtE0qcBgmPgnGkoYWMsYA9yYYubEieRBYsjxi1expzfu/GzRs615xT0VzcjgVYFkVSRRJAWpvuJbPnkC8l80XmygUBJmBFkX7Kz3QTpkX7RZ43mdslOAJ0uAqGalS5wE4ekTEfDRcal5K5VefF8RW/MT42IhkzgJAPn3sorl+/VljvEWfPnhVrjueLeoPliQ8FcLhy5bLW1zPPPC2Jwts3rsSf/envxfStS9HadBBTx09FZ++AVQr2tmN65lasLuJN2RHHRvCluBCd3Z0xOXVSPkWTExNa07eQwBseiYGR8diqHcbLr74uZsXW7n5sbJODRGzu7EomSQoRGL5vbsToYF8M9nXGcF9XNB3ux+LcfIyMTETv4HC8efFizK9sxGELa7umPUrSqAIF7AQNeTxcqHkgKU1sAOs583jFZSUP0LOQ9w6FWTPKWSd1PxJiFoFN7OnE3sUcZH4S926sb6hmQExHriZJ654exz2KabZ0bvOsdvcOxRikTiOGPI1N5qyAE51quPEem+ubYvmxFwLu4HVi/xaAJ9di6UaDC/FYApBCTMAcQuUCwAkMLPJ67T1Fvorch7XLz6QqoPj3wc2pfkzXC9cZB5dyewFHFd/JApR7sBnxYLOg8VN+VYOi/jryc8lDmoVtcFOpuxRmR66JB28h37+xqdC4BuuMqvs6H/7k92NaNM6fxntJUKpDG0dX99WMfsX3G39Hfy8M6zxLMz9L9QL2NBoAnKX8HVBE1oX8uQbV8dSpz1Azy2Zo1pl4vX2nzCIyg4Lc1iwTj80RsC3zz2xw5NgdAbA8+pnLcF6lBC7vDaPbMXtV++pubad4lx2onkhMoViou1ufOzs7KzlQapIA0cSkLT6CnAfcI3kKQG41+D9oVLz3Av7gu7+5I3Cmq0eHGoi9NKohuBkeHopbt24rgEJbFkQ6i5gE3DrBq2pUgOKkKEBRyRrylgFhQ2CRcUhKf/vwUIUbkgwST4qH0BqRUZIEDTT67i5R+VmEfC4bEAk9SQ2BCEE4wTj6qzdukMCiZW5kOAgWoVBLMZfDDgOtcxT8YRvA6tjfi/4h9INvxeL8kq6dBLrpsElBuujmUHKhUbe4YMnmAxoBdCyNFZonbL4cyCSDaTJJwtDb169NhSSB42N9bUOSUrzfyMhoKXpCT25Wck+wLHQV2ttt7aLIg8gkwJaGfUe7mg/c4/z8bInBmlQsNLLbrAESIIozbHpCv8qDkWKTizwqGKlQWRDIzo4zRz5Cvpfg86jD7KLaUZJRGBVJPTjqdRQqIsmKN10VEYv2XjZObDpF/G/Gh1BoSGRJVsLFyMYvJ1FHOohCYJV/S7qpBAQ0xxgvkgTmmfUKoaS36vnB/sGQE6QfRRcj+I14J7GBHZDzjUCKgKWlFQS9kWD8jpNJG+pJ31DeIDa3VZIBKmRrWxJedLyVFBT0tv0mnFC42ULyeaTpr+eU9MASYSgBF9XZiCUjLUFDwVJC59rNChU+i0F3MjQScZHIZxdpjZ4SM6YU4Xkf1tXE+IQ0E2v7RnmR+KLR6/qoGwGeB/yugw7JhGhONcpyHek1lhfqGfP5jI8N5lP2xWhCtIEzeLJ0ls1k5ZdDoa25VTRiDmoXbS3ZlcmIpcJcqGdNst9wkCtIATVc0NywlIREpwAn+as6/ESFesmAyYRRZB+hsXiJxr0YgyMtQYHhCGV7ZIqu5BlpL9BFnR1CCpoyzU6QBF0XFLk+Amubuia6vxiJFt8VBYglCTTt2o0DxorPTzaLYu4ipSSW1W7N81Ozr0lJuIzp0nxQRcJR7dUUrGiCSrO4JCg2603kd037D89aSfrhgQJBigJuHtk0k3FjveV6pDDua8jGlgPBXONCP6NRXuZ4BvTatwp6kO8JrViXNzMTQneVKMkGevp9Qb+K6EZyqbFdkH9C6kuGrfhupNdF8RFxI8TPgf2EOUFypQIVrIhytvh6U6rNDSUzMyiaHUoyAObf9Rs33eBtsumnWA2SKpBSvfdV3YsL9pqS+/txcuqkiiUgcPFakhl3xfIQSffWOKmwb4m5bKxQHDHDbk3PP5syaikWSbL80+PpgDrnTCYKJIisXUkOlufpxpJl7pjXQk3Kd8QNU91rCfT5sxGplHMjCyy5n6lYT0Fc7+nEgKRVSXL5d84PznSKMKCOeC71PqNYKm7qch8E+Nb3V3dXkgvMUcaKAndeJ8kwezUSGcgstSELsrcZ1cPDePrxx2Lm9p2oNLfGP/3izdhhDVVaorW7J46Njin+uX79liQnkSoiSQD1RILBWUxxFf+sU6emon/ArFCujZiFPYSCkmKXvX2brBb2g82cm1VM4dlNTU3KX+n8+QtqAiIjiW784489pv3wylWYoYX5Bfr99GmZy0pCA0Qx6LING1jLt6aC1J1RXNkUZiHX9g7i9OkpFcIw1qUJzFpDhgyU721MVXX9AAqa4/jEsVjf3JKpNPdf29qKZ596KrZWlyVRxGcsbWzGvaWVWCvsQhrfzCliLopf/T09cbh3EGsrq2rGEmM2t1WFvmS/Hh8/HteuXhWiVwa6re2lgGLZihaK/sRlNGDUpKoVDyYXXvCnQKqTourK6nJcunhZhUqfzaVYccC6ZgYa3c3vsX6PpDvdiGVOvvCVr8aPf/yTuLd4N1pam7SmQWC3V9rFnDjYQa4GaSCkNlaF0l2cW4tHHjoXU6dOxfdefFEMue0an9+sgpSk0mDBSmaQZnMyeGEcH0RnR2tMHT8mT5Tens6oSP7R8iQ8d9Y7htE+q5piaKBf4Bgk0Xjm83PzWpugUJkHSur38MfYj7au3rh45XbUDpHjoCHZqfuOA3x2IjZWlmJsZDC21hZjdHg4zj30UHz3+/8Yza0V+Y5sA+A4PBBABxYY8lBDA30xdvy4EPMAk8S2bK7E0sJiTB4/bmk5PTNkcbrNKFIxAaaf/aq0H9EAQA6t0mx0OXt6kcphC6UAx1yicCr5OPZgPAswtu9ok7/GQ2dPxj/85J/ihRc+pwQecBGz+iMfeUZs6QsXbsWf/OnX4+WXX42LF6/EH/3R13Xewby5fPV6/MHXvx6v/eIX8fIrr8njQbVdqfXZK0/M3WJmrHhDiG5Lozk+s2SaocKW6NPr4kAAMC7GDWPHNDTOZIou2TUzD1XwQ3JnayvGjo3ExNgx7VmAmdRUokixScxqo2fiTAr4FGVYv2fOnI3Z+bnY3iJuSe8u5rTPrPSEYh4zX5izrEPWE6AF9mXWDnEthfKLFy7obGIPdePVXk5ioArtTvwNEIEmkc8E9m3GxH5GLUXehbPL55e8b/ARau/QmuI5uwFh5itjBYOBWFHAFFj4hVHIIcC6JbZQrHdg9DTFVZgyNDj5Pvkb96emOvkGjODSIHfRtaoiqhgmhWkiRgPxJzlUYULyHFgnNClgd/AePCejvvM6LO/x8Y99TFIeP3/11bh05XL09Q0o36ApwrNB+owvzjJJ2MoUtV1nK9Jd2qKKPwTxCHlOMmYMErHkWCPwAJAd30d+GGljgeSOHdMzA+gnbyHFpAZbiK2d8roCMDkuYZ+Q7NfsrJsSTU1iPuGhxH6vuL5I2TqOc6yMXBT/SD9FRdrvwahIMIM8MQoCX80usaSP8kxfkRtbzEXJC5FXltyOcSDnTKk7xRlNlvnhrJWE9epqDA0MipF0/t13tX543jQq5ucW1PgfGhz0ZwMOamu1x0d7Wzz6yMOxMD8bC3N34s///A/i9rV3o/mwFqOD47G7cxCtnZ0xMDYQq3N3ZSK+tbYTfT39ce3axRgY7o/RYxPxDz95SQC2weHRuPj222Kq9A8di8PmtnjznYvRPzQa65t78da7F2J9Y0sFfLyvtgu4pLOtWVKU7S2H0dFaidGBPj332u5+7OxH3Ji5F1t7h2pUrG8QF9lLihoB++TW9oZyqJ2tHTWSNmFNF1YK84r7tqxMq74vKW6Yn2VdZOHeCPVkN8P2K1LCxJWlgSTgJUbW+0iBKZHSeNLwBJDAF3Ua1iQNB5qdLcTqysEd3xZcjv6ESdhXZM4EGqzti4HOM949OFQziLrO5pbjPRqNnModra1qgMCy2NuH6V5VjIMc3u7efmzvwdhuFsPRkuGOV7Mo/UvFCIULR54cys/qHY3C/i3o+3yfjFuzWP9ejYoHGxQPFvTzOnIVkMPyJXnIsl59phz97/1/u/9O8v0fvKYstt+XR5UmQxbgHxyTX9V4ea/xe69x0LU+wD65b0xKrpUgMDMVnWdk/kg9Mtns6bmSNZVUHOAsYX83cHQrnnrqKcXkzi8tQ575UO5NeQ95rt1fMysNkMIQz5w0c4vMq3QuwkqXnDzNlJqACvKDA7zGudfRLlAy59/Zc2flmcr+qzwfqcSt7ZhbgCHdrv0MphTA5zwDkAIkH11fXQs8gj9oVLzX7Pvge7/RI0CjgsXAZp2sCIJUDLmkT1loxiQQFPRUaGtvF3qJ4IyAhOSZxca/OZDoYGfxReYuCmj24t7MPTUeRLktRSYVPHa2JUlyXInMXty8dVOBMoEZCf2VK1e0yCcmjqsgg14zJnPIKyyv2NCNAoYK4c0YeXZEB1IK+1H8M9rixq2bQdCEvABo9ju378TuNtJBHOhdYoWwCdBokCFZf3/cuXNbCQabCJsC6AACGpnglsI1v3Pz5i2hEdG6ZRynZ6aFiCNxIVggeBTNtzBXMCmjCEVzSIeOdDE7VewgkJZxLaiqtva4dNlITOmvVluip6tXm7L0IWu7QmJKz5yErei1sqH6cDGSWIEo/y4+FQ1ciiP0SUr0FD1UIWIOjHrOilAejIlUvv8Qde+DhIHGCQcJgYIKRgTyFPy7MQs3pVnvlYWtpMLLZKggG8tF6rAvPhaNrAEVnTkA2lrVwOLLyZMLVTxHih8U7AhwCYRI5CjkwJrhg9j4k5mgwk4Vv4sW6Zdy8OvzVFBt0Z8kgzQtQPtxTRx4HCigU0iwaIiA0ONgyUYRAQWJlBHkTnBF1a4hqVK1aXbdONjUPRfij2STFBSVgrbRLEdajfXCX6Fw6pBnDIuevZsrHv80IfdrjGLnmTFXOTwr1VIEPwgVrCjquDlUIiFdln9XBzPoTzXEzKZwsfUo0GwMOBKRYEZAiyTddNBWKMpta71ToFLiVoyvxShh7GQS72I66CkaAQp0lYy7qZBeDSn7Yp+UXgV0vL+8Ccocr1MaypyhEMb+Inpw0fKnUJISZNk4Yf0zFyzFZuSfJKTKQuB1Gfiz79l02GtIc7jAXbhvIcDLnkkyketUmvVKlI1SZO709KKzu+6iu0ycKWw0Fss1+4VSRjqDBjD/VhO00aOEebe3HxPjx1QIYk4g+0Shg3ksT4UimcZ1ixJeJMMc/JKcJGXcRY4j1HxBvlMMzXWdKJ+6Z0dpVEq2xbJBivUzM9GzNJqYz0qzcfY/v6d9HlSoKIyMX4Zm+mFoX+juibmFeaPvuNbicUFB01/MieIdUeax15p9iyikgC4V0pkmQ1m78p0oLLT6+5T74d8UOgcGafTfqjMiQIrKE6k0yLxmvFaz6ZhMk+Pj4yrOsV9JK9iXaj3oMj/F0CiySQS/jBWFKIoSJHKgZy075kaWcWTF86a8T6IZdQYVv6BMZEjiXASgWVgMOAui9CjgMeoox7beUCieLVkAaUReHTWlnGikH0v9PXONCJXsZl35qxJRdNA5T42kPlQhSk2K0sDlfdR4gzlSZP/URCssQwqJnN0qcuJPwPlYjBQxWqUoO9TdEU88fC4WZuejqdIS7165FfPrm1Hp6Ii2zu4YgjW6sqriPTHI4vKSYpXjk5OSd5xfXJDECNr7+GkgI3ThwoXSUKLouK34yt4H9pFKyT7JvzTZjJ79Z2hkMEZGh8XA5P0AR7BukckkPrgmM203cZlMFF/Qfb948ZL2A97jzvS0mBsuuB3G8ePjKuiyVwgNjXEmJuInpySDwbiqeFbFuLBdTQXQ+AA2NG8PI05OTarpCzz67uycdLSfefLJ2ATxu7yivW11cyuWNzZjFQPtdsyvbQRJAUgIdQUMFB0tq8gz2uUzKGBWq4oria04h8SOK3MYRi1sExqm7GMqcLBvqHEAoxLktGeUwRHMmwHth0g/yWOgICtJ+pKVJSaX5tuhCm7o4ktGrwACfu/LX43vfvd7sbK+HN39SA11qiDTWmmN0aGxmJu5K5Q6pKz1zRWhrauVVkm5fOKTn4wLly5JJhQ9cs5/2Hc6m2UmXVVfNwELAAdgSHA/mKhKFehgLzrwNuBeVRg6UMNCSHnkC2vIMJltJf8m7t1CqJaz6+svMpLIVbbF+vZ+zC9txNp2LZqaYWbRrNmT7vfmxnpUkW1tOoxHzk7G0sJCPPLoY7G4tBJvvnMB6lkg3HpQofm/rzkCO4d5xV5XA+WKJ0m1RZ4fa8sUp3ZjYnzcsj1a23tq2qmpt7oqwBPzz1KD+zqXOA8AU/BlCVE/e7WWFCwa0c3cRxud8YBJMdDXE5/77Gfi5Z+9FBsba/aiePTR+F//5/8lnnn22XjskYfi3/27/yeeefZpMbmvXL4qlsVHnn1ObKP/49/+RTz2xIfi05/8VHznO9/TczMT0xrpzIlk6qmJvLvreE7NCINBiEvciHUjRs3b5hKbE8eJ8eEYVICjAhJgbGBRqPBeUPF8Bg2YpsMDm2GXArX9vKzXzp/MJbww1pGTlLwhRt3nlDMx12nIMo7ka8SvyJjyPYBpSNixZ5MP8VxYc8QzXAtxAUzYh849FG+++UYpWAIQadN64uxiz/AaJO/qqyP9Dc4w84HnV20za1PxDQ2f0jDgcTJHmLsqHMFIUnPBEmHMAzFvS1GJMVBzkoZvaTgKmEVzqMQmOjsSJVyYlcYHuASuGP+wrKcKpuOAXByXsm7ICXgurB1AauwRAiN0tselixdienpazQcKT1ns4zlzxnC/+KE8/fSHxSbHaFsMsILSTZai8mgk11qq2qc49zmzJHlaisHkkeTCPHsKvSnVlPE/98MZOEGTcG9P8oNZtBs7NqZ4XkxjAUCMNDei2OyxjCcMaCGHblODmPfhOiSzeOyYnsX84rxCNiPQLdvkOMNNcNWn9zxP9wogTXFOiV1g3PGVbFGunXgzGQ3S/pdpjyV1VKQVw92sYcaL8cgCqnxMWCsFRKVGTJHxI+c8PLBnIuxGipNrqyta4+SCN67fjKXllZg8jkQcz6CifXd2jlpFezz22KOxMH831lfm4o//+Ctx6Z1fyJNpamJKyg3Mz4nJsRgcHYjdja04PKjEyuJSXL9+RXPkzLmH483X34zBgcEYHqVR8W6MHxuL5s6eaG3rip+9/FqMHT8VO3uH8U8v/zz2D9k7D2JPa8Hxe3trc0wcG4qBns5oif1or1q+Fs+g7dphXJ+eiWUaFNUOHV8wKrh/5RTIzuzvycB6f9ceZlmQTR8Q8izJ1haGsvdacgV7eukM5f80rj5PBZgjji+MZj/Lg1gjZoUBtrsfrezLxMpiIBuMSU6WABQaFWusm+L1SANd51eZK6xv4hNYZxiKc552VKvygiJDJ7ZohrGMxyoymjoiYWk0S2KYed3VjgFxRQBbZiC+b/y5CksD37OOTjV9lS8VoGaD8s9RqFt2LDXoABUUlL5zCINtNF9Lvp0AqweL8/nvBxsG+UH5bPK98vs5ZmrEKa8027gBb1dvV+h7DSDSxptobJ7k+kkQUePr7msWlB882ERpBCJpP0+GeKkP3J//u56R99U4Do3v2zherkda4osz6cGx8/5p+bsEnyYor97drEO78EgpwBDA1T09dXCW82zXYXJv1rkrCdoCVGyouThpLcz+hnpMsu9zHJNRIVWM4mNqABfNcM63IgOe+f7hYTzy6KMCVAC6JNchNrLR/ZbOa8AmjMPY2KhyM/6Obx37H+AExecfMCoeWLcf/PM3fgTOdnVrAyH4AamPgTaB1/GJ43Hp0qW60RqxCAgVir+VaksslyYGiRpySCxoguWBvv5Y21gz9ZAAtjAZSE5pVBCMidLUgJ6o1axTD52dwvLMnWkVzk6ePKnxBaXI5stnE6DM3JsVGhD5J5JVFTyLRAaBU5pENe0fxNlTpxXcQqXd3N2OqdOnZKC1sbUheSId+NWqabVLy9KdphAxPjEWl69cKaaTRuUi75AoJ2ngQS0dH5NUwc5OLR56+CEVKdL0jXEBIQWtlSCPpJtDZvLEpGSHCB4pBKho2daqRgWSEssrKzE2Pq4ggWIImydJAggR7oXElzHEYJBCLGMDCp7Ahc0P5AByABgbekt1EKtCckEg2Thdgp6mM4LYRp8UNF3RyiV4NjoKZLipoEk55/mqqFiaCwrO92pCYan+dsC86C1UaBgMUCuhuu0YfVGKUPUudikk1+Vdyr95/mzURk7WVEB0odzzTVIA1RY9pwzwmUvoyzNXKCgNYJK6afNzkKvorhK8Z0MjacqSeirmscx17ldF6WLKxO/TaGPu0pzgetzNr8QhSMgihcY18z6JUqdAqUJ1Mb6V3ETRva7TFeon6/tFGEZiv99XBpKJiGKAKT7xXBg/aXzu7Na15JXYcK8yBMQQGRq9DW75PoWkDGREqX6fL+nmlwREBfmSMAnxUOR8hICqosGIIaWLTsxtzy0jaShOU7CHdSXTtaIhSmFdKD0luWaRsDeQiCfSKg1ECdKZ4hlMctCTQIKkUDGwMHCSps6aZj7QgLXshxMmISpKcZfnLRmrlqoQaTRZhVJPeq9QwvZE4bkmHZq1wBohmKChgy5qVUVIF40IhmH5sPZZ04xFFsNdt2fNGl1NEYpngHEfKMVsEEjqSQwA5leTmqgybcRTqLBw2G/5UhOFZumOUdnsFxQGSYyn79zRmmUvZb0kWoWigpsjxZ/G0aj07GXGu2vJIQdhrdr3pBWsn4FOO2J0qTCgqZ3Gv262ZTE79T9TioBrYL/PvTybr6kP6/PF3gbSFi7F92wu8WxhjoAuTs1iSQ8U9oBR1N77tKenkVxBSoEgZX2zR2ejQlIjZX7Xg/viueIEziwL9gk3uu842C0eDLmyHwy4pS2fYxEhxgB7PLIUTOhkcmTjQZ9TninPXxrj8tmB2j+mOcc6AkWXhQglL4Wlwtw8Slh8DkjuqZifS6ceybJSgKg3nkogr3O9FOVyv+bJUtTKPS+/n2yM3D54r0RDMuaJMk49ce7l6JpdnHCxyf9xpkqPHDYYmulDg54jsOOQcGptk0/UyNCQ5IwoanGvyFYIObVrVhrrAuQ0TR3JdiAlQ0N0pxbH+1rjq599PmbvTMd+c3u8celazG9sqzjb3denMZ6emVUcAsCANcfZPTQ0KFkMiq38HdNcEO8kRZw5Ms0WCyAbC+i4G9Ev1lQxpyXRp2DX2maZSJohgDVWVtYlK8f9Ep/xRXxAIdGHbsSZs2fUiEdSBGnK7q4eNUmyScW8wTtLwJHZWSHPKczAOjg1dSIWlxbEprMHbyUGBpC66o3bt6YlYybARWE7aM00VWRWzD4L+hRNadga2hco+MwvxMraevR0wwKlqA5rr037Oee1CrlIFYk1wT6IwSq69gcqusGc5YsxVCG2SJOyNgUQkNyL2bxGrMHw7ZKB6kefe07xGXEH+9rLL78cq2sbOrG4BpoBzI1s0knvvTBQeQ8nnjDZaKZvxZe+9OX4ux/+KGYX5qPaZmm52s5+VJua4kOPPBZbGxtqnLW1V2NjZ0PxdHNUYmNzPcbHj4l98/IrrwuNvbN7IFaD9qEi6cCZIpPy0oTj2ogLj48NR1dXu62lFZ8B7nFRLYKxI85ZsaY/UnyFgSW2LzrfnActLZZiVMGJz9mPaG6LG3dmY21jO/YPrfMu+QRkyShugdo8OIhHzk7E2LHRuHbtRnzpq1+Nv/n2f421jS0QB7HBdVSrQqYSTzH3uKfVlZX6/g3beerEybh2/ZqKn6xD9P3Zh1ZX1uLcQ+fixo2bNj9vadaZyHiL4aiNzgVl9jr5lhQ/Je6NZ5RAlOGBQZ1F7chF4fnW2x2feP75ePvtN+Ptt9+K3//aC3Hj+m35oXzjG/9cQKyXXvqZ5t6Xv/yVePHFH6mQ+a//h/8+fvwPP403334n/vAPvxZd3T3xrW/9lZkExVOIfcxxUZMaa/aGoxCGdK5/ArwDAAAgAElEQVTl61xIN0BFjCDY2wXWwP3A0GYeZsFBsTTfLx5/yZxVwwlWKsx0/CYKMyNNvbd39jRPMobJs5Bzj2J7f19PjIwMxuLivMaQ4gcNBorJ7Hs0TLe2NyU9O3tvztrxQvj7bOG58lw4k4iXfud3fifGxsfqjF4zfc2qUBGmxMEysz1ArgUZvz2td+LqjW3LRCI/6XULW31PJrh5hqr5WORXHXYUcE4DgEloWeUVBk9wbykxQ5yWMQXPKs/XlEni/pI1oqL/wZ72J84wYhliTDdHLcHKmUODlL1Je3Ycxuuvva5GMeA4fGdYuxS3aayqCCzErJvo/+q/+1fx6i9eFXghtdJhVwnsA/sWPytYJwWARXym6waooFyiKnYYZw0MAdf8jgp/ikcCnzKkwTrE2CfIZK2xB87PL6j5xGdzvzrT6/OTGNJgkDqgqGLAn7wYFRM3yyeF39caZ2/q6PA1FhN3PjtlIsk1BCYqIJzMCxQncNbWZVn8QBm7zFUkY8icKuAJg6osV6mCogp8lvjiZ5znnAWK75ph89KkddMX1h7gQZoUx8ZG1fBfXVmSpNCTTz4V5y9ciPmFpTh96lTx4rQHysyd22pEP/3Uk3Hr5vVYWZ6P/+bP/jDe/MXPorWyr+bmrWvX9OwGhgak6MAaPwY7vbYb65trceP6rTg+fjzeeetdMaH6h4fj/JtvxiRG2O3dsb9XiQsXrkb/4Hhs1vbjjXfOxwZxDFKIuwb8cb9IxML27KhWYqi/J7o72mLu3j3Jm3V098Y7l6/FrXsrks2juWGWliWZyKWUP9P0aqpoLSfghgkjJq3iT8A4BsIISFDybb6ndV0kOLN5LABNyQtZq4wVZ8ZebVvNe8sim1Pd3gaD3Psjzdtu+XEO6LNq+9uKc2kgsB/tHRjAQy4Fi0k5k2eL5uZwb3d0tbZrXSDzLRDbYQgMocaw8l2zbtS42qfZjr9ns86EVMEgr6eRBnCFGHAD6Sj2LhhGiYxJ1nMDq0cZTMlj8u9HALjSAC1ArYx566CiBo+D92MpNKbZDzYGGn/2Xq/z+r0f4NgYd+ff830bWc6Nv5vfFzCwgOMefF/niAoSf+mrnkslGKs0cB584YNNnDzPXcy3eXu+Fw199h55GhWpx3psIz86cnjvy4LUSTnBwLAEAlEP0WeWXEt5Ha8DPClArudaAgc0DyU/a7CKG0OHiumyYWec3f2NqrxPxocxTMaupQOtLgBowIA3f6xY/G1tjt/n5iXpia8N3+d8pj7JHsm1ERew3jhLOZO5b2I2wFJi+X7QqHi/pfLB939TR+B0uzXHaVQkpZYDEAqwGgSloWAd6yYdhiTbqxghCt2yJzYC3XKK8irKFKrT9s5uNGF+1lbV6whwenr7pGEpc0YFfwRNB6YGdtM1jaiWDYrAlgXIl3QTi341hy+BoZFVRl1yWJD4QJ8nUYN2DrYHXUqSaJK1dhBwzU0KXJBngkaqjWr/IM6cPq3fYVOgQNbe2WFTwNxsmw4VJGZTBuQk6HmKFjQd0AGGSULSoWKf6POWj6LJAMKSA5Fgjg2ShMBIz4Iq3d+PY8dGFbzLs2NwUMGWqOCFZs3hzTXyLIxQIrkk2elQMZZquSnfpfh0cHCU+NccCGbRFUQfQThBeSYBGbQgIcAzJBE2ws90bjZW0dQwbtTGzkZuRCPPM9GLkgQqurckkZsbW7pvxgn6MMUcdaxB7Sr5tj55Btv2Q7BEkBI6JCdKcKvAtBi8qqCxC30UIy0XFvgZ14cuOGPRP9AnGjSFPA6zm7duqbg0Pj6hZhcNDZJ7AjgKgZKQUHBmiQ4Q1SAterpAUHYZuSyTW6PYuA/mYVVFASOY83kRWPF8QBby7Eq8VbwEjIbQ6wX/dLEwD+9fPv3fv1ngUL+gcov/hBojhdqdArLclwI4DttS+WsMRpTgZnEyUWcPBF0PXheHvFBP6RtSzO4U6ylZwCTSyFxYU8Q2SlSEmnHa7iJdi9YX61JmZiUhFYIN9KRQd5bQIWEiuZVJZPE4SS17MWIKEi1NrWHBcJibamndXzOGCutIUkQuaOb+lR4M7Bspm8Tz53PFPksN/2IkblNaFwuRsAPhS2PB0k9mfWSwJ6o+SVR/v1hdFP78BIsWb/Es0Roo8gsKyqQry/eMHHZiZpMvsX5Eia8WQ3AjURn7ZPLwC6wX7hFGF8060Na5v/Kn9T6tF5zJi1GA1sRmDPhZMi9ISDHzMqvLchPSaZZPxY6ls0C9ymzOs8coejcYLGFl3406S6LoxSOXRzLB++X9ZcODe7WvhYvO2scLvIhnzX0wvpxheXZJIoRkqdDX83k0IoryewR9vJ49QnugkNalyaLg1QhZPjJ/P/8k0WO/47Pz/RqbE41/NyqJpp6ROwwGDXEkSJxIFZqz5qwbykZ/WVtf+xCNxjbki7YV0LK3Y6ZtzXsb/iZbUojTAiLwdfjz1VhAI7wg82GFcP+5LjKRYSwb0WL5fbHEdilMuaAkz5QGc+18Hc9fKNbisZH+GEKAF7Qe9yhWDa8jEZXMleUlpiYn1DAEEAGr8sTUpOYr18ntUOhBDobCtlg7sA+rmFEvK2nAVBtUKcX4i5evinnpa3KCw25zrKMp/uCLn4rFezOxsdcU52/ejZtzy9HWjREryL7uqB1E3Lw9o2YjZzYNdBC3yKYsLS7L/2VF5qoTmocUSHieLTIm97q1NJ2LQG4GWr6GwjO+MPv7NfmVDI0MqSBGUkKCQhHrkUce0XjcvHmzzD+vLeQtQFG+8855zSPee2b6bl2Gi/V2bBTNciQlLZuEnBCxCsWWnp4uxSE8Iwo2gDDA9UM1B6lJQQjkKXIdFJLYu/ZrtTh5ckosBBVBWqrxxhtv6F4Zd9YlRQL2f85VELGsZ2nDrxJLNCnedLESjwmkc1qib4D1O6vnwufympSDNFCBhqhlP9Jc27FBi4p0n/vs7yrxI7a9evVavPLqq1GrIVXUo+v23njUwOba5dkCs6JIjcAQoAHGnP7cZz8rj4o5tMgxcQB4sIuZeFucPXkqaqWArnOWCgkSFMjkNUfMzd+LRx99WOybq1evRzTRkFEK7eJsk5t2nFWO+SJ6RfPfUQMNs9LRkaHYXF/TWCLlA+uJAnGlGtEqHf6K5iINCq23Cp5mAA6M3KPproJoczW2VWxtjrmFtbg7tyBkKQwPe9RRoNiJYeRQttcDftvvfuZ34p13z6v41NPXGweMf1MlVtbWgp2I861/cFCIP/wqkOigUcg+QBPliSeeULGUBpyaEBubMXViUmv42PgxAWTYPyh05rmc8p3Mc+Y945n7Smd7uzzliC1ZS/Kn2bE3C7E3HhUgt9Gm//BTT8a3v/O9+MgzH5L325tvvql9/amnnpbXxX/+q7+W/wMApb/+62/Hpz7123FiaireeffteOfdC/HMMx+OwcHh+C9/8x0VGJAwU2wOKxY5qh2ATOkFQ4HQcaCa4CoKm23K2nYMbl+c+n5X9nidf3WWWcp+Oqbw/oz8FQCPFkvOHhpckAAbEPesHX7AupanFOCcDlgB1ai2VGJmZiYuX7oS+7VQcwmwgjwIt9YlMTg6Mhw3b9xSvmZAAnHHluIGPo/YDd+cRLQTJ+2U+IXzx1JLLpKq4LNvD0CfBc4/4DOSWyQQQ3uvzHvb9XsugllyTXGz4jKv00SpSi6qSJHyeyqkwgTAl6LIE8q7orVVcyPPmXwPN1UsrypGGoxHad3bR4J1whiQV6kpSjF1y4yOvEakfYm3kF7FNNrXhjynq/DykMNzbtdn08AwjbSQ/xTxMGuF/a6nu1dzRL5hNIUqFE8xQXcjkz/5PnGlwFiFYcRnmPFsticfSxGcL5rwiimbmtREJ/fKs5zrdBwAa8sxmOLowkRgzEEwky/xxeu87pjHfs8sUno+u2iZxXHyJsaQr8a4OouOmddlnMDvZexAHJixigFHTgS4TsueWIIzTcZ1fQcHkjPyPDGzkN/ivTD35pwBOIJiw+VLl2N5eVH7CXsSTClktviZmy94OWyq+c5cP3vmtPba+fnp+Jd//s/jrVdeiu7WSpw+czIun39X8RKyfoyvJbMHoxtpJljTaxvyXXnjtde1l/IcMDlnbNt7B2NvN+L61dvR3TMca4DIJNF7GIel6cR+LFbK7i7CbNFaOVSTYvL4mKSyVzfW4+69hbi7sBKbe0hUI51lXxjiHoAOpHT8Gxkp9gnid41xkw3dM9Hi2WSsafCjAW6s3fTdSS9G7wM2n7dcGusO9mBTtDY7vt7cRF7KZeMdgHoOT+oAL/Ka3p6u6JCk3n6sLOPh0xHLMhWHBeI9gedP/k3soDoB5vAlD889iL0ctLy8MZHKqdHYhVVQYJoi5R7q+gC+9HZ3CaxFnYBza3ZuQcVr9io1xZO7WccM+i/O74+AhNmwyEL1EfjniD2Q64O5nuObMXIZkvf848Emhf79wPUkUK/esExETxbOG8y080MaGw7OPUrOWdZZ5sBqEhfJ17yvxvvL5suvaqY01jLycx+8WTUD6nt+qQE1MDMM4rFEoMFqTiKTzcjeLU8vSc2HcuOsF1DX817ggdMcL0oI7hB4L7MvmKXsxGpXw815B000wDnZGFbjojC85CVJ36OoKtT9qTTRj3wt7cNntgaNRMkKl/ngdccz8P4LA5tck32d85S/w8ZT7U01lKr2MthF1KHIMalnbW9u6PpHhkc+aFT8qoX1wc9+M0fgYcy76nI7loaQ9FAFBM2K0S61mgNT9JOrLdFBsozW3/aOgjmhHEFYgr5BmqAkjwQrnRihYdpWFlxnp9kUw0PDCiAIUCRjUmmKycnj+qzbN29pQT/80FkVmG/p3zUhZGmi3JmZiTvTM9Hd06Xuv0zp2jusQ8o1koBGkyiDA739CiDmF+ajdngQPX09Mve6dfuODmFuHuQ/BlcEZtK539+XFM6Nm7dEyWUzTEQBCOQqWtWgFCgqdCHxgK7tQhw/Mamu55Wr10TRt1wTJtvdon4SBMOWGAcxu7YmOnZ6LRA4Qb9m41JQXYIuEIVGAzmgJsghKOQ1W9vo2hldsLiwrOCejjMat3UPh3AxPw3P0owapA8FBcaGZ5DB4y6oJiHYipRCSZzyUFPwWSRhhL4vHgrJ9uBz2FQJ8kDGgaCT1r4K5wS4NkETqkjv4wJ+FumSfpeHYiKus+gshGw5rBJxAnWbOegmgo2ouSc+Q8VdAv2ebhUsOJgoQlJ85lmTkDM+PcX421IMaB7j37Dtwoholj5EGSchew4PhRxlXdTo5JeinA5nTMykWes9QTT2EjHWD/1EQxVKbSlTv+8mkvfc+IK6lJCK1qVdkUbZhVZv4JU1RDWP8H9h3EsBk7WS9N2kpesaywclGv29LqyR8qpmA6Z+DXJe/E5K1zDeyB70D4CIblMhkuRDgUJpQhD0qriu8aXcZhRNNhfMnDDjo05blmkywc6ekaOlgMx4kYCzDlzQMsIfIQx+lsVS3g9mFr8P2lfMrKIdaW+KosV6cKCCIwX+lIhygOqkgL8ki0FzguSLRm2RluFeqsWPQw1aii5ilDjx4vmnSZYRfv5skm+jzb1GxB4o+sr1xFIBGU3EDt0nhUQ10QoSE6RSXZP6EB3qYRX+KGrfvHHTe9jqiptlpeDvwnJBjqhIYONSnpXNfpHJahKi3ehD++SAJuc+aNKoAVHuJanSkqwoDIOceyrUl0Q3pZ14nfXlN7Ru7XFhLW/LFpj6LP3kgqxz8Eej3CgyJHeQgGPNZjFezdWynjNIbgyi8+8klUeNiiPGhhouBQHvRoXnqO/BjW/OJJrd2ejPJND7uItY+eViidkhKXM0PkajYlmN0iz2J3rWBZvitVIaG9wPBVGeCY1z5ieIHBUj6o2KTOIdsLMPe46YtVCmYPG/8WuSedGY0DQmPI0Nl7zHxgJGNoSy+ZcFDq2pAhKw/ISfv35XQ+o1msi/TIZ49jQDKKbz/NOXQCy/IodQbyAXI12MMVmzFGzlraJEparmMec718TvM2e1x+7VYqTtIH7/c78dm6vLsby1HzfnV+Pi7bvRjNZyT3f09vZLR/rS1etqmjI/YeDQrEDOkaIFjSpABTTbBgYHhBinCE6CzrPkXinME7PIYLTFBRbOTNDzNNlBzk+dnFLT5fKVy/K8Ii7BpPuRhx/WtRMfWJLG2RESNytrNlylCNnR1qFYh7FsqVTVxLDW+ar2APYu4jbkfmju9/b1BF486SHFHIYlkedHc6WqGAZDa+I/sw634kOPP6amP2edvYa2JfU4w+/v7MZAP95mFBGdGLPfak0fUNTY0t4o2byapZhoctBQmJm5q/2F+ULzhr2V905mnVCjkmJMCRybG9NAOHZsRGOkcQcwsbUVGxRQiqcP3+P8z/mZ8gHEGOyJOi2KPw/j94XPfyFefPHFWFxZ1tmivYJiX1TixPi4imIL8ws6ymUMDtBiby96ertifWNVJq1I7V25di1amtvj4JD9AH+XihhMfO3tusmK1KHkCveRtqnFztam5LZYqMyL1dVlxcYUo5CqVOOec/3AjSg1/ItfQV1esuzFnL+YtW5t70VTczXmFpbjsKlZskGGodLnYX21RU9nR+xsrMrvYXB4KF78wU9i5NhQ7CBdhT8CcVZre3T19KjpfebMOTVY+F0KQQbOWLqS8RZTFd+JlWXJn/E1eXLShfiKi2e6f7wZCoOY9+F7bGXyWYC9KMS1i3LEYfKvoPG1tBxdRbZm6vh4/PzV1+Kb/+LrsbS0GLdu34yOjp54+sNPxHf+63diZ+cgXvjaV+KHP/i7WF9bia++8IJYcCsqfO3Fxz7+XPzwhz+Ombv34g/+4AXlHD/72T9pnEDi8ifIfeZ3Xce6BE5u0NsHwXGQC2GcfSUkk6cIz421zx4stmClWc0Io/jxiLBXA2uDmBp0NbEwsS/zIxmT7D1GpTuSBBRlBt5h7NZAD2/ExPhozM3Ox0s//VmQh+1s11QcZD/q7IYpBUsV+Z4+gcrYixKRClrabAmfrdlwqVFtLbKJbJ++P4qLND/tXcRXo8RfE/lgKaLxXjJGlZkpRUsDOvg+MYUYpRRoio8FMb1AbsW/RO+t4jZjaTBWxuqJCicnIMZnH+CZ8DrlqMXfhkIVc0dNFPkumb3Muqmf18VowdiEQxt/l8YI++geeWRvj/ZzsQ0xFkcednNLkma7tR37rpQiceYI2it2amL8KW4sch7MCz07oWh9HezbZo2bkZJzzuewUegCKnB/JRZmfFg7NEG492SP5Z6neKpBB14ssZolgsh1+VxyKL6f+zPvnajjjAdy7yFG5r2JXVjLWYTMGCIbRVkI9X04DnHMgaRaopRdkMwYnNwXcGTmGirgl3XF2DIGZovYL4b5RAGdxiXXxdjguwmzqKurI86de0iNeKSfTpw4ofkOEI+9b3lpUcXAqRPH1fxcXZ6PP/2Tr8Wr//j3MdjTEadPnYiL599VzHf8xIm68TVsATVbmyoxNDEW2yvrsTC/GEuLC2JHvvX2W5Kwbu3A97Aprl25E+0dfbG5u8dEFpOCGj0Fd9h/8l7Z3dae1tvVFtWm0DqGP8Peu7SyHuev3JRHBb8vDxitecvEUvBXbqp9webvaoKVsyGL0cwLNTnZTwWwQnq6teQ6jtc4N2jcZ42C82dtfcPAADEnWqO9tUXgUoq9SCGjNKHCMaAMKQtYOpI4JH+nu8sydDBAMctmP8X/KvcC2CA0WQ1SQFIaVuq+mJPtrVXJ4gpoCLOGxmJRLOCzK1XGwEBWjLvxI1XNp9vAWMblzt05xX8YEsOOy7z9wZz3we+XlNsY/oYfvl9R3vv+EQvqwff/Vf9+sCHQ2ARofM/3+uzG1+Y1KLcsZ5Eix3IzjQ2rPH/rOXUyHYoc3YPX++Dn5M8br/1X3X82jrPmk+eGWV7kBt7ntMbrTVXXkMi5APgQzzl3JTbzfpJsd84wQ0sBcZQGQ2H681h076XyIYnSAr4WWHEfVQVLaPOnakzFKzIlBOvNqPIZ9mCiJmcGtcFc9qTM62prB/hFPYZ4pxoPP3wuzp+/KPDx4EC/9hKAkQBI+JP9j+s/dfqkzihqCCv42NZqYqAi8/gBo+L/z8r64LW/ESPw0RNTJRCwYai0Rrc5LLaF6jTVnqI2i6wmSSGkCECpk6iqidHWrmCIoJxgmsCNLyEzOAzKoQQdFQQZTQ02EiGmRCs0auPxxx8VvXr23qw2l4fOnVOAiRwVZnygnEh+kVeanrmrzYrCAUV3mUsTMHPYHhzKQ4NmxejQsDYVZA529mtx+tzZmF9cVBFJiBc2pNa26O50l/3qtWsqeCPP9Oabb+mgZgMhIOczCGig3S8uLOqeOVyRWQA9OXXqpGSlKIzQfBnsd6BHcE3Qh5kjB+2ZM6fV3KCI5mK7mQroN2ZjhKAMlsC7757XxsZBbHPxDqFlSGq6ujtKsYlkzaa57gQb5cL9sZkSeKk4QpAAym53V7IEoLPZhLlfFQiFZCAJ82bO5s+foDp4PxB5BPRKVEiqhc47KqpyYMiIjsSH91dnmOZVj4IjijdzCwsqAtCoUUJKcFrQ7EpySmAqiZVS1GtE8SqgpUhZjJlJVoX0JmgBpbS5WYoZW0IgkaDyJxs88l9QdplfbPyWf/A4seEneomClhMFJ8EZSPcPOLGWBi4oFRpxdLNpbGBkXA5FnjHrhi8dulLIcDGzjh6wtoaySgcMSdm8v5BZ30Teg1DR2KjIYKMePMmk0g3ARHDogCyJkEylE/WVMkbZBCiIBT2LUrRPpkXjpqb3Lr+TQQXF5xyjRF0osaDJ09oi3VbuVsEGBy0I43IteC8wX3WdMrx2ACWTyHIdrCXGnOIFxcYMEglkXaQ28p91xHqieGvjaj/rlGQ6uo+m6OunWXsYS8uYyJpRn/Jnkk8ojTHmkWRASoEu5bz0Wj3jJs1t1oGRdUa5UbAy+oKioHUlaZJmYZ31mYkpEixqiGHmrrXrBoSS5oKe0zwDTdmKzIdRh+iLI8+Rvjfch/ZuFeNqSiKMcDyMkeFBIWj5HPZk1jTrH1kNI7ltAmrmls3uGTeh+IvHCMk3xVkK8iC8KawjN8TgEZyZ6XTEFGDcsiGe7AkzKor03AOUZeYRhtQ8ZzEqCuPAQSgIUz/nRLo4wCagzcJzq66PPTZZHUp8GhgVuT4fDNh5HY0Kxp+irJso7AdGdbqJ7EKUmEG5Z5WmFHOAwhEyDxk0m6HmRkZjMqHgHOR/8cHgmsSoWFnR3lO/xqKrr9dLI5iiV9HZrjMqdpSMs6cfNSqMZuOVAiHUGzWWB+Be6/J1RU+d+2P+IZcntHpZh1lkyGvK4kRj8SFfz2sy8c0GDZ/N35mXmZTUGxTlPLFxJ825qsa5XrwoSRUSiuNjx1zcrrYITMGXAQ9ox9vAnrMTvwCYPV5Dbh4S7JtFiGzStPZwNf6ly78R7S1NMd7VHJ/9+Idje2MtljZ249bCRly7OyvpJ5qaFFjnl1ZjcQkELECFZZtpDw9r/d1FlqGzS2gsJByZh9euXhPzjsIgE9jyDPtGvBcGGIUBSfpUy/5QjFCRsLt+/VqsrW/G0GC//LCQxaRIYiCDmQHc05kzp4TOstdWu/abu7Pz0Ybs4s6OJKnEQNqvKY6yhIPl6Ggm8HrmOvs0BQOaKSSIzS34PxlJDrqfvQ9UfFdnm5DQ+N6wd3AeM86tbe26TpivktbCc2JoqMjctaqAx1yRwaFkiSzb5QLivhohgFwMXLCBpuK14kdCTJKoa/ZZATkOKOwxt8wTGh4a0PNiLrCWb925HXt7yEM4weNmMp4xWANWGoVKPGoGYg8pKiHfzej4ype/FN///vflpYSRt9bV4WFMjk3EsaFhyaEqfpM5uQE+zHMYEDTSaFZgTD47txjt7V1RqbQWE0+Koi6QEjPxPJEFksdAk+UZ0VVHx4K9u4PkVtIeezZJpbkjD4EeNYhhG/D5krmptIg9wvknySAl2LtRbXWjZLu2HwuLK2K/cd2wGZsxhEbGaHsrxkaGonpIA2M/nnnm2Xj9jTdjbnElWlqb47CpImkRGhU9ff2xsU0Twok5QI2UBCH2nUOObWREcTANZOM5mhTvCwkrVHtzvclH0p1gAuZRGplKTpEmnmQbzBwQQ7u1Gj1IwWoeNUdfd3d88nd+Oy6ef0dec5/4xCfEfvo3/+bfxmc/+xnF23hPPP/88wIIvfPOuzqTn/voR7V2/7f//S/iU5/+uMyQ//2//7/jsceeiE99+hPx1tvvxPe+92I0Nbk456aFiycq2mfhV4ycFp2/NOFoKKGTz3xgTyImBr2NDjxAKfanjEFVhKd5VZiCKr4pHoXZ261i3L279yyts7OrPYfvEeN/7KMf0/6D3JsRmfbCIEZ45qlHhRz/+x/9OKpVcgczPfHA2uMZhwEdGKNPTp6IV199VXMQ5D8FYZ3bMDUUS/n5IZlEnsU5wh7Kz9LHg9cLvFJBMg5Wkr1nOigoaU+wxJLlmKwznuxQo1DNFjBryo04/mNuE5MQ69OQzZhaEoC7xbdMr3UBnC/HT24eNn7x/uwvkuUqYCMVtkp8flR8s2+FgUpVAXJ8zg9Fa3ubcqXmajXefOst5XbyzaAYjA8e8SD5AYWy4m/F9bs4ZvY290HMgGcI+xAxj1oipSFBg46xovmdTAMxDyWp2qbxZe5lE8nPwKwCnimguGQ58H03muw5ls0dFy/t84c8GM0Kgy0c050+fSamZ+6o6cEXn93YiMg8NcFm2dBoBGek9FaCGPI6kuHimMJsUd4v4wTmimPaXZ1ZnBmSY0EqDmCO2OiO/8xAcrOZL2LIU6emYnRkNC5duhhbMDIH+uUpde2aGxV4PhEnM/bkhuSIoyOD8cjD5+L6tSvR2VaJf/bHX4uXf/DdGOhuj1MnJ+PKpQs6z4fGx2N2elpr9MTpUzF3dyZm5+bj6Wc+LIApEnoAACAASURBVG+T5oGBWL1zWzHNz/7pZzF6bCza2gHwNcfF89djeGg8llbX4/rNOyrA41HBvrpbIxYizm+O4YG+6OvuiNbmiPHREd0Xvj7rW7WYWViOantPbEtejXORZ2iwnfyJlFI2KZ4bGRyS5ybxE+BIcuZsKCXgxg2/EHBTMbNnoiVryF+KHCnntf3RLM3MGb+7TUzQFX0DfWoKLC8vKT/IuFcXbsqRGjK8e3eX6wzsgUKvHxy6OCvWvEF+apiKMRFxwOfjDdVckRfR7taOACzsHYAqmEM0VNSYYzpIStNs5dbS8GguSHhAt4vL684jBZjFs8tM6aOvX9dcMHgqGyuNAJ58j8bv5evu24h+3T80ZqmdcETsIK5PJrk+w/D8ukfFg82DzD2yJpD7Y8bwuS6TRWUG5pFpunL5X9OoeK/GxK+/vaMxvq8JA/BL9UUkt3mOPgPsM2bmjJl6zqEEQpOEHj4lVqkwVst1Fclak/cALBP70EA3AcWKdBgBIns2+21r1XUD9h3eA5AMj8HMC9iqxQumgKs8/gYesvdqj8RHKaULJauIFLpZHLwcL1jug/UDMIk9aXUVVZB+xcTs6TCaienZm+7enY0nn3oilpeWY21tVU1Yah3k34rNP5B++nXT7YOf/6aNwCRBdJESQlKBoAdzFhIHOtUEgyxkIz0q0dXjRH1u9p61SKExE3xKMmRXjQPJOJQuOosc6Sc2EBoOlhuqKuDikEyES39/tyjFvJ7iAwEUaHw2LQoIUOLdNGiNDWl32yCU10P/TtM1KPccdJt0+ptb4qEzZ91YWF6KNuR7+npEGSdBBRVDEExQefb0aSHsQUMS4CA7QIIkE+NmCuEg+Yy4BjGgZkqENKhpghBsgsqnWSIjNKHym+oIhOOTx+PWTYKVVm0sbCpGxtj4lTGm0Hj37kysra6LXUK6zfXRpCAA4YvAkfEj4YsmIwgoFNCp5XAnyQRJyRunZh9j5AOnSQV9EgYaCdwAQS8BKXJVMlAE5b3vpMAFwUONB4cACAl+VwG9oZF1pCLXxusIAlWYre1JY48kyjI1LpjzM5J+obP5/GJixO83dtTzsFJxV9fSZC1i9KxBOwpFSuGiWUknwROIGNOISWSrGhuCKH6O94c8Jjo74+qV63FickLjSvEIDwmCODZ+mnBVzPGKbA4BJ+/BZ4GYZC4QBEobvlD1uR8M5jkAWRNJZW4MtDNxcJBimrmKnCmbVOZy4yF/315SkFxqTjR8CQHg/y9f5W+F2mgEeklMitxRNgBUQCxFskTUNH7+EbX0vXc14/VKgOH6vpqEokOWREnfkpY5tFsX4GFdgYaWES4mooWZQBBCgZYkNm+KaSZ/hQ439GiigkzlkOcZkViYlXNUvKWZAZoG2QdJb+0apZVWG/zd0gEeK5qfJL82fO8uBnIUSS0vRMCRbAXuBYTPETLS929/Bq957YltbQrSZQQt7WrT//mSVjiBtrwnzA5xUyc9BcqYgdxrNuWdAKUeRCKJQ/OgaFyajYEkFmb1mMKj0+vgyA1IP5OUyADVKx3x4meRDAP2GK5NyWs4OFOCgZlZR7v2LWTsEnXC+kJPk4KI5GsosFHoLIyF9AqxJ4ALOxkAp++NitEliKyjWtQMqaqoKl3rjY1SYC/MrAZWhKSfYDKUgoSL1Xs2g+zpFW3WJqeYpblZYHPIIxZSNhCcqJv1kI0KmpuJjvUeZS3f3KuOGhVuQPC7nAOgH5HrycBeDK+GRgXvVf88MfaKrnWTfY9AyahYUQpf6b2hREpzvUg/iQ1pjwrmmhsV25It5HeVkJDYJ9OoFP85r2Q8V2QdFOwnrUJz5ahBbZSixyubE1x/o4SEmjalAZnI2EbZh9xXcoyyuJeNE12nkLVHDCnN9+Jpwhmn5LuwfsT6bK7o3KZxD2PSzSyQvJU4ceJ49Pf3xObmevT19qtQx5xv6+jUnGXVgq6kIJVsHprZmAefHGiPz3z0ydje2IiljR0xKm7NLUdLZ4eSG+QLaVTM3J2N/v4+nXEUmSh4co4iccMZBRJzbDyln65rL6KAn+tDHjA7ls80gqtVyCg8DLhX7gc2Rk9Pt5IUkpduocaQWjqpscI3QMWZYgx7+tTJ2NnZVBMGhC/7BAbIaYhJsYQzHq8Linoba+tKBFVUkneGz/aUgxRLUQUDGlrswW72ATp4+OGHJHfEhnfr5o06YlkToRT1QEguraxFPx5b+GGge4y8Eqj+vZrQppLapEABErT4KDFO3Xhj3LGfFHJCxJaNxTbPOc6VFkk2IHvhguauGEbPP//x+OhzH1UMy1r83osvCpwh89AdjEJpHCLf431YjeNi0ix2XNmwbWi7F5//3Ofju9/9bqxL672YI7MX1fbjYx95NtaXl/XeC0uLOsPYZxnT9XUK++gKI9G5HfsHFFpgploKgCI2zQOKmYzL8sJSQdC3ygi6r6c72ttbY311WWwJ9nq8CtRwa3LCnWslkbTcC8WoNB4mnuW8TYlEPCkw1J6+N6smRV//sIAcNMol8bFbE3qfzxnsRM+/LQYGh2J8ciJ+8IO/U8GIAq2AME0VNSoA3SRymwYec4rnxV5KjHn16lVJbiaTmjiWeJvkfHYB8M3ROcu1U2BU0YinDNsA1G4HnmBNsbm6KcYlewDzl3gTdC0+TStLC2pmHh8bi6ee/FC8/tqb8cYbr8f/+D/96/irv/pryZJ85cufl2cc14QB/WOPfSi+9a3/qDnwwgu/F3/zt3+j5/OVr3xBLEEaNKyFL3zxy/HjH/8kbt2eVtxgyQhLTyH7wrqhANjS0irEL/sl65z51NHZoSYccdDc/ILW2daOcwByHmJQ4lPmI540PAvmMutd8/6gEs9+5Ck1N1974y01k9gza7Ac5V0V8Sff/EacP38+fvbyK1oD5HE4VfAZH332yXjmmY/EP/7kH+Pd81diaHCojsTHc6W1jYZBJW7emonHH3tYa/zChfMqPFpK70DjnNreYnlgtk1OULzkGAuuXyagAqHZE4HCkc4DCsfbW24sl2Y/5zVzhfiDBqY8LSS/wfcBmtio2n4Obrrwp6SWiHUorEo+0WxYNSHLVzKgUyaKHMFnVzZRjMDnnoSABdBV2Cw8N/kuYQDe6mYABXNiE+IhclLLTx6oSQdY5JVXX4nrN26ISSffmOJJpiJp8bzIPJLnjeyT9c+9hhlzgG/sg5IDKWc4kk7MP8sEmn2XMYQYwgKZ+Qzmd1iHjGmC22hUNLIs6gNUN4M1UE1ss+I1KV9JSWfas4DzjXwpm/u8R2Pe4OduI3aukfXb+MX9ZUE0gRs6D4rEpJousIdNqagDOuRJAfNGUnYgih176P2ayZFhJhq0lHB45S6Hh4oh8fSgQQdD99Kly2L+4dnCXoTH09LKSpycOukzl7x0bz/u3p3W/vfkE0/E7Vs342BvJ775L16IV/7hR9HbXo3TJ4/HhXffjf6BgRiePBHXLl2M1pZqjI6OxPLKUmysbcTI2DE1JbZru9GLwf32RiwtLgooOTAwGhtrtbh4/mqcOnkuFpbW4vKV65pnaxubxdjZuXJ3Z1uMDPapSdF0UIvuAhQ4jJZoaeuKSzduxjZ4kkoL1CVJVTF3nJ/CviWXCe2PyTziPiUlmo1V5aEASSiuunnF76sZztzM4jDMcJlvW1ZWNZh8H4ACsBuLXxn7Ps8T9p/Pgi17vAlQYCm7SoulOVnPYkkUZQTWGV8rq0tqAG9t21h8jzxOTWBkpw9juL8/NqlLRJMa1YN9A9o7aK4ynxfXVnmxYg0h7GnEqyXrL0Bqa5vrsVsjrhFhUe/1S/n0fTM51175ZmEA5UsS+JRNuFyT+fMc8/ve8oF/NBbrdS0NeX/mkf6VoyxdMXppXLgVVF7R8At5bY2AqcbGSeaYqtUUr5OM5/N3ck/K93rw/v6/NCoa7085cANbI3Mw1Q3kddmiWINagRmDboxzHqjVVWdgqaDimxYqzo1XeYwCaMW/ocgJJkBODQ3VBpx/s9enXw7zmviGWlsyVuXvxV6jNXXEuHPzxqAw3X8B9LGWyNjUQFeOSrzSVs9HyVOlBrG9HVMnJ7VfyzNlfaPOYobdyJpDUQbZJ/YvwGWAA+/dnRWoobujS3sv58cHjYpftbI++Nlv5AiM7KF/2aMgms3dAYRRGhQCSbYTOaEAQZIaA3Hv3l0FrRw8dP0oPFIgQVZkZW1VQSaLTt4QHSzGfSX0FNc62ztUyEn0JQgxvngdC3dxYUEBKgwHmhXoFN+duRsjI8MxdfJk3BB9c0HIUiF8m6vagDiMLBfTFE0Hh9HR2hZ93faH4NqQfoIKiLn1NNrsFPO5f5gSkye0ySgIxgi6r1dGrKBgCGBc9LdZGZ4cjAv0LAqoBJ4g2QhaVtfXhKSleSO0AUWBgQFvIPIssA4v2s1CihcEH8V0NJhBKBldAGX1QIacoG3UkGi39jCFSxUnmnzcsrFvbdpoxwhrG5mrkQS1eJfiboc6tPw+wZALbC7KEdRCyddbNjVpLiD/IIMy2jmViqQECCZsyOg9V11q6d6XINE/qQcvQkoqyLG+HuNOIELTKOXF8rDTgVH0dXXIpuxOKe5xP8xDgl9pSBeztDxQOTSYYyQbjC0NJJJgiiArNKl00LWoA00wxlgzH12IcUE2NWJJKITkkoyFA+NE+KhJUuYayTyHnzSLy51zIDJfSCZVQJB+tgNALrqOLClRhBsV5eBN6uFRlHS0p5RifuMmk02LxrCqMXbJJkKjpJPkJFR8dqOHJIkiJgwLFe5L3JPeAQpe74+M6pdQXAHqSYUDJUdIoscjaVKXYrKzGgE0QShFdV7LM4UZwZjz/DiUsxEAwjPlnjIYImiiEFBH42ouWE81X5No+2yE6jOkI21d47pfSAkqQEeomacGiQMNAgcxA4o2tCinZczWKJzXkRwFcSRkBbJCNP66tK+AviCR4sumz5auUrhC46u/z9R+DKiLnqYL4NbaNMLD5szWOXZB0oiOon1dkEFK8IqZM9dsbx3LrXHPQqkVNDv3S8EHmRL2RQI0CphCFeN902wUrqSwKKC2w/bqidp+rW7+rUYIjAkZjFkrW9dIQal4YTBIyX5wod3yBMlQcMKduaWZK/UGQByqIEzSu06Du5iLq5io5N8mZ5IHgkmm5oMTWEkztTQLZUWBNwsipg2bdZOFd6EKtccY4ZhBeEo/La3QqKA5ceRRwd/rwXpZ2+kvw3OkoMqezzmQ+3MumsakIP+ueymMNq5RjYoVPCqs7Z3XWP9dxpeiRGGcsVe6kF+L0ZERGbrSqNCYSQqRQpn1XYX8LTT/lKhQ0p9m4mWtowmcTDrGL9kXjQ2eTMRyD8/kIxOPZEtkoznHoBGhlfuh3qPQr7NIbmkTr0Ezu0BR+dkyp1lvkxPH1RDE94g1IYp2tSWmpk4oMSdJHpuY0HNX0zAqMTs3p4b0hQsX1dAUExFfEwAVu7U4NdAWX/7UR2NnfT3mVrfixvxKXLkzHxX8Xzo7oq9vIDa3a3Hj9rRMojmTiGdAaXL28J8aGItLMT5xXPsV0k88Z9ZSyttRaCbhZ76mJMgu+07Vuub8iZQXDU3iH6EWSbpre9Ii5+yi0KrUrTw3NG63N9fUAHjksUdja2MzLl2+6oKDGEwRzz33kbg7M63izhzro6Wqoib7CuwedjQTh9gHk1FLEofkSqvul3gCYImKPkODat6hVS9fMphai8Qt6/JCYB+BVeJ5Ypm+nDOck7w+G6rWZTczFp+uO3emNa4g7DlLMT6WHEbZf3K/NmiFcXACSfx17uxpgWqYx/z+rTtGrHIuZ4zh+MueKUI3y2sARk6nPo/nknvUF7/whfjbv/0b6aGn5EiLIHGH8Vs0RNbXxKblvdGsd+HMTb+DQ6THqrG2tqEi9tbmTuzWDIJBzgu5Lkzse7p6ZDAtZFwpBPb3dUeTWCM8wyYxdyhyMqfFSCn+W4wzclmph8zeSbOW3+P8E3BC8kIwAShiVVUUW1ndiI4ue6qIUVF8bDjHDmigHBzEow+dkQTSw488rD+JPCmAESO6l9AUA0NDKuoTdyHzyLdB2LPP4A0D8yjBRoCPkBiCUYEcK+fUakEHsj+QrAMgaeJ95GHkBmZKlBJPwmo2QAFfktbQs6Bg3RQxNDAQtZ3t6OroiN/62HPxl//pv8Tvfua3tS7fPX9ec+yRRx7VXvDzn78eX/z85wT0efHFH8bXvvaCGEU//8WrWgNPPvmk9okf/PCH8cgjj8Vjj+O3segGMM8SDwdJia4qf+G8hkElo+gdwFzEFjt65hMTYzL2ffHFH6iZtaXnUmKypohHHn4ojo2PxUsvvRTbWzWzdkzi0xr5xG8/r0bfSz97RbrtjnUoOtp4GdYPvmqXL182mwMGQJXmQbOAUMxr1jGm4m+/c14NBbEXwt44rAf2T9YLzdCnn35KZz6xFF/sT5zhRpgWI/qmwqItvhTEzexfKVvE2mJfhnHlxpaRrRSLKMjk2V4en1XFC/vO+5pgbyW+Mzs3PSky7pNcXPFxMjrf7HF+rvMPRgiMuE6QuWbA1JsY0vMnfizG9iXOE2tJ0q+WhOJ+sqjOMwA5C5iNuJa9jrmAT6EaBJi+F5YWcjwuslsyzGep0bkUnKQwUOSSYGikvJNjIcuXsNcjHcS5Tl6n+JwxVPHVBTO+xz7L31lXahC1tKhRSMPBfhYZ+zgmRH6VHJeYj7OBMaSRSE3AMaFZBsRa5Khm7xo4lgVJx2Rm6vN38igBCjfMiuJLMVRhk2aMx/eyKJnyuI4TDUA0o9sACgEoO9rdNCd+aWDGCKQoaVfnHwkk4ZmnPx0NC5hcN25cl8fVsdER1ReQkeYZTk2d1DrmXNvd2hbwAbQ+Jtuz9+7G7tZGfOOPvhJvvPpS9HZU49TUZLzz1hs6X8ampmLm9u3ixdcWe7s7sbm+Gf1DQ2q237x9J46fnoq+ITyc7F3XFNWYvjUXN2/MxFD/sVhd3453LlxSXA6oifhuGzZjRPT3dkZnW0sM9HZFZ3s1Dms7Ykm0tnfH8tpWzMwtRktHd2wisyS2Nsy2Jp1FsHxoJKuIuo/3iE3mOcdzHrKHai4V9HmWuFMaNAurYkFIzQBpaTcwdO7vulZDXCCfUnLM4qfTS20Jr6Jmx5OAMNk7XIAIeX11drbF9nbNzKzC3HBhFkY1EpYGqxI37TDfJaNbif3aYQz198by0opVESoVrW/2fICDrJPd/VpsbG+rvoEnqeIZWBXyo6jYS2x9QyyWOhtO3lE+0xxWZULu/cFfDX/PQnkptud6yPg4/8zYOXOHfKfGP+9rUDQ2GMTeVBey/vJ6iyIvqkH2WfHNA3WEXLMPxu0PNhZyTVoa0+C7o7ys3H1hZGl0GkBf73VPjbnP+91rI5Cp8TpT6lZAt0Nfh2KAZMoVBrXBOuSPbkbo3DRC82i8BLD1vpLsCzGE6iDR9JWwHwZ7EnWArCNIFYMcvzB4zaLEo4nmt6WRdRUFEUmeLSCl6pKWpCdt4/fM4AVMi3x4h2pGxLmjx0ZiaWlF7Es+m/OSOlUCdBKkPDE+rniFPZY8Pj0jAV180Kj4VbPwg5/9Ro7A4E5NOuNZkCVwJeHJTZCAh8NeiI1aTQcp6KzF+XnRu/kehXM1A7a2hLqVXEbRFCWwSdSEkRYUb03JVcG3tiujN4Lws+fOxM7utgyveN3ZM2eiraUaN27eVOB16tQpIUan796L+fk5HcJGX7joLhklbToHMtuk6ID+81D/QFy7eSP2MJKc8AJHi1YBEIFsxaZbULBT03x07FhcvEghw3rvJAsUqZEjATnBvUguoRzQC4tLopLSqFBxjAaOEEUV6dhSoCeZAbWPtAfBHPeUGpEczCRRFL5hmzjhdMApTejWNn2WNjcSZYpyVaQBLHUCmieTdw5jNTUqlimi8QA1jJ1bupPb0IjNECEhUfG/tVXITRAzJAIkLRRaaGpIS7sE3VksI4A1mqIYdufm3OoiJ4Evxz2JKkWlNKfGiF1B0oEbPy5OFdqkAPku5gtpXTRLFYBKr9modRcOTEUVGqqg1Wy4bXkl5k+e6eslAbZ+vhttUEPZ/Jm7oNmse2t6sRDLSDcUbdsMLGTKJ1QUiT7avKXoTMFVkjMO4BmbZCIl6tONClO9k8miAL5ImiSqvJGJ0LihZNPhwU3GjYGjVoU1hUtwJVqhhddAh6aef2OAk5JKjeZ0SSV98LOSwcT3uc4iZ11PWNTMKQe27rVIZCn40sOQq5mKQQSUFBdUUNfvQOHe1tpUUaIYRCOfwDwFHSwpo9JUcFHNzYFELWbgnShxPpPAOYtrnrueY/XgDEkzGbGbNs3P8xlYJo2GK4E0TTYXfSjuZFLNdagZU9gNLAMQsMwBPetSZZBGKoiOUtjmvglQQBCyB4l9oEDHBR7el/2V9UohirWtAE06w/bMYf6xHlg/NEz53fQHYs2S3Eu2Sk1Ffz5jRDILSu7uvbt6T8YxG9WgEfVsg+Qbb4gWo33ld2CNbRdW3BDO91bBQKwZszlIKuxv4oRYzaD62jxKWpUkFcmBo4DeDR0Sc84i5NvcbLAptwsb2ag4kpfirGFueT5VikcFhtZO+P2VRaGjBmFKQzlBM13YWs81oRs114pXeiZ19YSiwbBOATbGwV1dOgdpVCTyL1kJeY/eCxLF7cZLJtpjY+PSSZdRYTGRzjGXETxa7RSedV/2yUBehDkM6iYbFUKCCxnF/KRAYTSPEZ2Mk1lGPJtEzmWSwtlCYSkbwVrzKXdVRrKxUMHfGwsRuWe+VwKS+3cWLxLFpWQoTa2Zl0VbuKRG+oNzkL3Zsj9NgZ8HoAESWhfAzf4APekemmWfQLMzVEi10ARC3uXd8xdVRJb0UWkStzUfxmhbU/zRVz4ZmysrcWd+JWbXd+PKzHzs7u9Lp7+7uzdW1rfj1p2Z6Ovt1lkOiCI9UThTOVfYryg8UVS9N3tP5zbobwoIkusQc49zxI1LsxZh/uG3BXvkICbGJ2JwaCDOX7hoP7DeHu2ReFQQH+Czkcwv5i1F0MODmoAYZ8+cjStXrwvJyDPmC7AA8kGc25hm07jv7um1/FJrq+abmnkUSoqMgtg3SLO0GjEPEp1ji0IWcjpTkyeEpKRRZBaQ9XunZ+6pQLC+6c8kluB3tF/La8fJvgAWRVJNjYqSW1Js4Nlm42Dm3l3J0nC/jDFnSF1XXuub+U1TersARTCDNwsHyVLWA4hK5gd7KAOfkjJq2iGXJP1jCh4dOr/kXVIkWr7w+c/L22AN7xg1PI3iZ56emjwRg319koUCJX9AMRbaAdr5tZ3o7e0q0pr7MnI/PGR9wV6AiUuTYEVNIslfbe2I+UpsDfWCuYvcEQ0LvEW4b+aLGKzbOyp4k9im1IqABUXDmeJQxjbyesAgt8gCtrZ1xO4eWujrYsAwF73+D302w2Rsa4vV+bl4+onHtI5ef+vdOHaMRsm2zmjMtGkera9jOu4YFTkNeYM1SGuxxvl9GmuAgCg88VncC7E210QMdFQYOGLP0fiDscTrmZuScmxtK/Fzax1lDbKWxlt3R4cKkWdPn4yf/Pin8d/+y2/G7Tt3YvrOzWjv6Ipnn30mvvUfviWvmc997rPx13/9t0EI941vfjP+8R9+qvnDmnvs8UfiP/3lf4zafkv8/gtfih/+6Edx7fqd+PM//7N4++134t3zl3TOEBtIUmJnJx566HScPn06vvOdF6O5ybrsYnBWLFsCw+PZZ56Jv/g//y95fJCvqJEl6bKIDz/9uPaOl19+WevV8hGtKoIzF2GQWf51wYwXwFN4BLYC8moXeCqbni7gAoKgGMPcqqphOjN9Lz732c/Fqz9/LV57nWJrr7XSmoivdwq4wTJNp05OKR9hPYgpXsA7rB/WnovfjqcE7mBfptG0vqHrzJhNsW7xQ6MoWN/zmytqsktamELrYegM0xkFsEKFMo8DuVGy/10E8n/ZkCDPSjPyPMd4vSXdAB7tas8kZiJOUuMBeTsktHZtBE7MIlm64odlY3AzXpPJYfYfwBXHtUfN9EOdywk025TkGkasgFd6S6PCnkAARGha0HBkrZF3SyareFWRhxmQcWTOTnOahgOFdiGNJedrkIaylkolpqamtEeDtpUc8v5+XQKT6+DfeSYr7sq8IBnqRb6SucQ1O0d37MkXQDoj7Q0MS1BC5j7M3Ywbk1muqKskY41FXL6XbDbeh8/JJoVi9eLfR8GRfYjXElcq9ysGtqwfno89KtzQFNiyFDS1Lmu7cXLqhGIypBL5N+wQgCy370zH/MKSpKGYv+yP2xtbyuExrT41dSKuXbsSlYPd+MY3/llceP0VmWlPTo7HL155OYjVRiYm4sa162KddfX1xcbyctS2tmNkbDxaWqv6jJa2ahw/OSm/zp6Bwdha34nrl2/F9PRCtFW7Y6d2EMvI3ZHLKZ+sxO7evpqtHI07W+sx0NsZfd3tsb+Ll0Z3rG3sxubOfty6OxebmHAX42miUBr2SOmKrXDoZi7emuwZ+UUMIImbAp7Q8y1eQenbxV7IV+YJ7A8AAhSHFwAWz8Om5TvKWSzJ6rnF3oAUX39vr+XJOBN2d7X/y8uqdhDd3R36PRLKOtJfcp3tAq/CTGNu8NkAH5ZWN+Q3weY3Ojwc92bnZJSd8QSfTz5EPYM9CBYja5v7TTCu4lnYeB3tsY48JflMkTJGaeO9vpxHuL6UhXLmZmNDoLEZkTH+gzHwg9JJuTayttK4XuqxMnlyA6ui/gzLX+o9ibLOVEdppGEk0r/hz8bPrb9fYTLlfWSj8cEGSmOz48E8oPHfvG89viuf/X6NjTwT7m/o7Neln5gvxFT2JLKksnJs3af3aA4yzh/tDw2NCjPwmi1VWepy8hMSkx2mF15mbr5z1pr9ddSAV5PiMGKbJmGp26ghXvIz1EY4rzJfAsQtPzpJGLI3FVBxblPlLgAAIABJREFUk2X0c57L/7TFcpyAsmFVvPvOBeVlNOrIEwAXUAOkYcH6JPb6yEc+rH/byJtG3pZiyImx8Q8aFe+5ej/45m/0CEyVgJ9COoEewUC9kFFpEjJPEgLFhZ6/k5DMz83VaYTICCWjAtf5ZZKuYniqwpEakRUVCEBsEViTNHF4UqQzQm4/nvvoh3WAQdPnNZhOsZFQYLYMAoZxO0qsWPYU1dTZb6kq2IOSxSGIpMkWydfBQZw7gyF3W9y8dVNGOmOTx2N5ZVkyRgTINFfYLDDTpggKe4ODCC8KkiqSJ4IXNhyKDkIEN1VienpGzQeQ+xg+UoSA7QFCi6SYz+agdld0VwWVK1euaoMiEF+BxVDQRLwPSfKJE5Nik9y4eSfOnj2l5g9NmuMTE3VDNRoXHNp8BkgE0KQkgIcHJL6WSSGxcfGiouBsdHTYBWvJWFW02VMAtNaou9SW9nKBlECOTVjSVFBG0dUuzWmeGQgrmip5cCvAkal2qLDAZ3LtBBpzs3N6xhwy/X39QgSBlOfwAsUEqkgHW0EDCP1PENxgOpvIXBdGS+G1IPbNFrCxLoE5Y818NKqpQwU/5iwyZiQmBPIzM9MKaJnvMneEwaKg3tIwPGMKMwTcSLAQMHZ3dUiPnMSANWKfAMtrMf9gJFDUZE7ZFPlAyYLQ7GIGIMlltLwRAzaMVaOtjN+DAUrjxpJUzsp7BCv1cXlgJ5KRc0GuqdBcEE35MBO54OszWsCFzyMQSSYM+h01Plzsd1G20BwbPlfNioLkv69Rod/HJNXJmMaj6IGCKONgVhELVkwrAYiTX8aJPYHCpM19rZ1KwuJmoQdEyawKbDTjmLu70hlnfwApmk0rU0FNnzeq15R8viT1xmceEKzYhA30TbJ3SMJIXKU1Ly3mUjBHKqBIGzF/ZLZFslE+lPsTO0lI3S6NAR4/1oovZvIl6WNtEcgoGSzJG7rmy8ur0pUnGDf74ghcw7UyXhSJkJ4hSRHFtTSEE3XI/Of3Bwf6tGcgWZdIGRL/TPjZm1UEK2aILig7mCP5USGrlfs0E8UNhCPCNM9QSJyCtLNGsxuH+VoH5bkWjijouQZ4zhRS2ac4N8xW8Z7mcS8G1Cr2HwWUydLgOSTzL1k92VxJ9kM2STSXZSJumTGujUYFeyJyKG64NEzyhjWY33Yg7xYgewlMLprhyUbM4DsD/CzSc50kUbyOOc55oUY2jIoGqZakFrtpDgoSY3Hmpo0/3bQ4UOK8ub2pfZbCR8rUZZPBBVmzJi3JZ+1xBe1CLTsZA4WL5IYSTpLmwjpLJHwmUI0JTu7TiY7knnPs3y9Iyj1I41OaN5xfXLeQ9ZVKXUc7kyUVTYrfCL5VgCYEosCMGYmtarOLX80kH1tx9uw5U8BbWuS7xRlNUkAcwRphnT333LNx/vw7cWJsOLbv3YzTo/3R390dS5u78cq7V2Jxay9a2vEaQA6kKw6bWmL67pzOYOYnjQrYpMhKgq7l7GM/4XkgR0NT0E1Yo2e5LzN7bMqaSFeaAx2dnJcu0NGsQ/6JmIiCIck3DVWKoawpZEYyOWJ8zpw+HfNzd62928zz39OeQKLGs2QPY18ETIApM+sI6R3OzpyHxG7IFk3fuaPx4X4AQlCQBe2FDBFzhhiNMQYIgEQGRWLiEkpMFOgwjcb4GwNr1iIeT9ba9x7Oe6XWvAp6kn5CHqtDhVPGhnmADxifB7uC5ww7ksKGEO2lWEnxjuaTJOW0DPHiwUOnV+uRe/h/2XuzJzuv68pzZ+bNeZ4TiRkEwBkkJYqWKJqkBlKiRMmSqxzVUY6KinZ0dL10/0ndD91VXdVdLlu2REuWZEuiRVOkOIogARDzkEgAOSHnOW/Hb62zb16mQbui39RBKBQAc7j3u993zj57r73W2leuXRPDXU3hGlvZ1yPCiNa4VQ7YE2oGjK7Bg61feMGNChiaLi43NTOAgniwt7dcKzniTtyevqOcliKTnISZZZz/qG5vTtzSjANSHMDjRr0WzaQmsUQBCO/cua28ad/4vljGi3xpQU2h9dVVMe/yLCTXXVhYUY7HBiJ+AFqzfiBj8Bz5bJOTt6Onh0HwHnrNPRweGRHDD+sT5mxxvYwJNmAAsFyRsnZrhSK8Ek88cSrefPNNxVtUJd29vTE1BUFnXM0p4t3YvjHNIiEP5XzmubHmsJ5hL5hoUlWOmESUrp5uNXf4Oc4eM+JdzJPHsb/4TJ5t45waFaJsagqILDAEEGxtLXq6OmQ19tI3vhG/+cdfy4b1809+TvnF//Wf/yJefvkFNTl+/do78f0/+obi9rvvvCtbhSe/8KSu/c//21/HS998TvnfL1/9bbz87a8p//+rH/4w/uRf/w/x+uu/iXff+0DxINWQxKuj990Xpx59KP7iL3/ohnk2uQWiNsrz/vjx4/GTn/xtVIlJzU16Jn19/co9Oeu5N7wWZCXObvIV5U3E5i3PawFgb21vVYxhLXBO0uAaHBrSPTxz5ozW7TRzATUIuRJPfeFJMU5f/dWvVRedOvW4GqAfnv0oWpqbor2zTWdHKj+Vr3R2xq3JmWhvd74kcLk8H3IryDxNKK0KQcEkEeJDRSpyWxp6ZpvidgKKBSjUuVfO776+Aa1ZGl8ATZDiVJO2mpDEa4rMkfOsNKPElp38bTBzQ7khFrTEOGoszfjYJHfaVvwxmcdNBocKn3ep8Pc8tRbZ3GkdljyU9WaiBsGJneIYZVC2UfMY+czUS2oaYYtVadLcCp5JWys1RlXMcimBtiDBdKhZAUhG3ULeoCaL1CoeWk0MIQ8BXKdBa0tFN4iUdbCOZMNj8kO+Ru0+VatqcCSA6LPYmQufwfmNiRuZ5/DcWXuAYeRi5LvE8BsTVolmHlOf13ANrF32T+YbOasv87r6/CHzAz5jKqWSbCTCQiGh8cFkSap8ZrOWv+d1SFFCs7/Rw+VR9nF/0rZrbW1F1k+cDygq2C+cq55Nc0414EMPP6R7NCSrqMW4Ozejdc5+BeugOWBFxRsxNtAbYyP98eHpD9TkHztwQI0KnCI6+7pjdX5BcztXV9ZkA3p7ejp6+vticHgg3vjtb+OFb70U0dQap9/+MOZml6KreyBW1rZiQ7ZlrRrETYxbXl2XIpRh042xFVtrK9HT1RadbS3R1sacl4jpu4tx9sKVWFrfjkaamW2tUuaJwAgI2twixZsahhFqzqBc49wFP+Hcx4aa5655i2V2HvkC9bkVyFbkpZKJXaOZfwD/K55fyXrR/tGcs51YW2dmBUpe3ttKwNbmRikvbOPVqBjMOdLR2aV9yvmTNWvm1cTPtrZm1d4QZvlMNK65HmqRYebQTc/UZnSpYQf5pBDIIJUODQxGpYHzBOxiVRgFw8tRZYARMLh7jRqmDGbfBeU/KUnIetEzC7PuLLMlS4Kbv8vfGS9rzZe6eXz1+XPuiWwK5F6p5dYFS7pXoyIbJnq9+iTbfZzaXv20/Lv+63sbKvW5fX2jov538tqzyVL/Wfme81wTODMe7f189XGq/vX8+66raDjJIQBFmuy1bW3MPudc10w7FKjURUnV3LHC1q8PWQAlOo0OVLNWC6NKJKdinfPaWcfJCqqo3/hM/I7IPk0NsVXiJRZrRFD2kQbYr7EmyRWdQ9VslLEsJF6rfmXGUbFmh5jSSl5DzgbxqjEOHT6oXGnqzmyM7RsVfgHmhv0pe4zZg6irDx85onm4qEqxuYV0QQxlbX+mqPjvWe2f/czv1R3oWzX7nsODhIfilw2chwmAh2Tw8odfje7eHnUkGRwon/7Nrehob695UwK6wxgkA8qADhuCYAUwjuxd/qAF8DUQQnHG8C4PiuN6OFBIOtoECsNCo/hvDxj5gN53pqcNKAOirG+oEMWWAcagCstqVYnDiWPHVbQDQxGkGpqbBEATDAiBBAKK0v379hdQFLl8t16bZoKAOIFYLpo4zEeHmSVxS8UTSSFHM4MlKSwABWBPEl9d+LfKNgUWM6C8bFw2XViQSHP/bEVTjX1jYwJleX+eBQn/3OxdNVZSScA9BWTh4F5dWy5JQlfMTDPI1gmkfGnlncug8BYl4RnwlpZgp2OfYEA6Gb/5+pZAGyBy0W92hAZfF1sGAibFQP5R00HvQ0Hh4oG5IICyAA8cMPK15Hca3FDhBpGYaMh3sQcikCe46YF2LgxSZeHDjmHsBQium++RTOu0KOGzw4wieIsVuDCvooDrnJyclKUG3wOMYS1SJPvQcxOCNUoXm/fU5yvMLQAVromvcShhJaK1Xho5/DyfnwOIJM6gXQGWC3s8D2YDJrvzO3LexL0CyG5qtPvdWtOCmuseDQzLQ4rqo8yjqP9aDi8XM6qwlDzCuk7sWpdc6bq9yD41xjmt2LWQylTPv0ESaSVEMv35KrYjXvNNsn6i6aOEoVC+bZ1R1XMkQeVZsTZhk6p4LRZWnvXg2Q8AWgBy/LxtnACzU67uTozmhjCsjgK6KDT4269J0wPJfZviHutf1jkU60U6rHVZGgyak6CGWYLDZmgInC8zJbQ3C/OLGwlAQRxQvBLQX+yPxPxFCYWt3JrANtlIaejodm2YuxUuqcqpyl6DGJsxq9YcK00fGjjsKYFnG5sqUHgNAXxlpoUaQYUJSdRLyyaZqkvFZRajPGvLjAPHGsd03ltAAT65pIyac4NMfPf+Z79RyXzOuylKBxJODdGsYv00rLheX9jXPNaLQiCVEtlw4TVJLInNAHoUnznDQg2Kun3qpey9mYoJv07szqi463u0uyP8w7XEvWyF+qYLAAuABXGmnjEoAKI0YMVQK4ApZwCxnv1Bc+LggQMCCDjXxOQB5Cprwr7MtmtI5hf3kJ/ie6OjY2qkYb8ocE9DFa2oAhivNQhlnefzXoA26kPZibnZgkUB972e5VQPMuRZk4GgFtNKc6G+4PgkQOLfyEKOfycrM0EjWZ/JM9zABPuHdYitihrqRTkkO4x9+3Sd7GHiAj97d46GMTGlK27cuBFHjh7xfJbWVgE+xHWAchqYLhTWpTi8ceNatDY2xOG+tnj68QdidWEhVrYb48zVWzExuySvY8+YGhAD8sr1iejr5cz3MG0ICBQPPDspS+fuxpGjR1Vgf3Tmo/IsYdi7qcLz4WyAfWXLA2TisCCZD7KqcxiABSYiKgad/d2dys8gL7AXGbzne+3YxoyK1tamOP/xx7LvgKlLw7yzw4Op/X+a6zlAcEdND+IbMSAl8bzm2XPnSw7QKMa8nR7dEGtpaxGw/9ipRzXbiv9zpnrwblP0DQyImHHz5q3Y2kGZ0FrAN8C5NudrrW3KUcgHerp7df2AKICTAinbeUYGqWlEDPQPSDmTTWz2Ic9bFqOypLHlJTMAiE8vfP1rIibw+ufPn4+333knKs0MkXYTXHYsGwZQM26w7m1xSRyy5YoZgU3xwte+Fj/60Y9ivdg5cg+G+vtjeWFJeSrrDjusZYAyxT0Do8RbwDJYntzXxQUa785jzQBmjpJtV0kF+RnWshUfW2LqonHDNmpwsMcgVMkxJibvaH1gk4flD18fHGJo+aYUG1j+kCsCbvNezhtXpY5jTdA8m7u7IBXE8jKDz8lFYbwD3jabJYwFzPpqnDh5v4hCrEU34t2MZ00B2HFfAWTJe9o63DSkuPfslnntc1jhttorHs/KT6qxtrGm7/O65OecnTy3JEoo/0EB3WaGOo2KklLo2rE4Iy9GxdzW6hkCB/fti/uOHYkzH52NmZmp+P73vxt/8Rd/FT29/fHiC8/Hj175Gz3rBx98UH71P/zhD7WGn3nmy/G//e//MQ4eHIuvfe3ZeO21X8fa6kY8/PAjas5Agnj77Xfj6vVJzYYgflrF0hj7x0djbN++uHj+guxFDey3OL8strQiJrEuelAwr+qe8nMeoOz4Swwh1pHjUAvxPHmP+44e0ffYW+xjZl6orils8m9/6yX58J8593FR7KFcMhniqSdPxQMn748f/+RnMT83Hw89/Gg89tjj8e7778aZs2eUb0QjOY2BJZ4ruT77nFqM65IdH17eqENr6k9bfOqsg/TSAADoXJucOxup/B7rBWKPUkQNizeYxf7i+bKH87OSR7CGmNPBPYLEQaxnr0vpUGZVJAs/rTJNdPJnoH7hnKuZuRSiShKEnOta9cT1JijPM+Pfabdb3xT1HAvyHchynlvB+cQ9IveEGMeJDDhFDUlzj7qUwcvsZ88CYobDsmsLnQO2RKVZBnDl5gtNvQbPBtrBv7/Hysu6+VA+R0teW3Ifqe5LcyYbuSgEsrmQ56+afGL77v7Jn8GWjbh6Z+qOrksKvLFR1baZE+TZndfDcybvYf/zh5+r5bt7zny+z3Pn+lJ9blICDTHn+8prpLK0Xz6f1bM7csCznrxUz7J8xlBJdjXr2g/kkiatrSovQsk1ceOGauyR0SHlyxcvXdYaY1A4jdb9+8fj5o0bUjEQt0+euC8uXjgf/b2d8cJXvhxvvf5q7B8ZiPGRwbh08YLwiLHxA7JaI+ZoLtH6WrS38qy3o621PW6QJwz0xvDIUNy6c1vWToOj47EwvxqXL01EV/dQLK9vqKFRaW7V91HjyF5vcyMefOBkPPbog3F3bjqmJq7F9iYDfWGOt8bC8npM3J6JrYbmWN/cFvAvkoIGaTNXqj2YR0QcqW5DFuwV2GmrWDe4PL/NamSdjZw7su722ae8scxPYr2wPzWwuA6EZo1KkZSz08rgYsW/YitLlsJ5yrPEiovnlPNaTMQqlqpldqYbpiZYQI4gb2AtUq+oIbm6KpKZcmXY9mIapbLEJECqqs6WVpEqyCkFYletqtKZyAyNpaVYL/PZ0hrI9nMlOuzKFUpubJJYgu/1zYL6fLiW19apiXLPZL2SezFz5PpcOWsMERo/sUs/sWNrzhSOg8rMreS/xy9lQ+FeL/f/pVFR38DIHCrPjmxUZEyprwnyc+d15Hsn0SzjHPbmxEea4Xw2nr/s5IulpM6FNccb1pmcBmTIoUWkW5DvK3cX1fpWL2sdF1eXbMLVnAL0inYsSVIZN1T5sWpmamjbuJO/q1FSDeU5kGPTXlCqwk0s1K22b9CEFNfE7CtyN2bC8vuQKwaHBuR4IjLaBrjmovar7Oi7u0VaAlfjHvO9a9dv+HE32JYegt1njYpP3SyffeP39Q6MhWce0NEmyfpEo6KpUX65JKWSvrKx2lr1/6UFigknBBSWSlAADGRnYA9fJIyyBmK47dq6fp7NT5BJWap8EGG6bG3H4cMHyjC365LHnzx5XIEEVj4sh+HREc84mLsrJiHyeOIyr724uBJj4wwSXdfvDPT3RVuFAi/UxT/78ccawv3IE6d0sN2+dbvmp4hNEb6/JDUM/Ka43Ld/PC5euKhCTnYoTZapAkC0KGjSENjWNZBwcujhe01HF3BEZwSfvbVVjRC8EImd2CkhY+ewVrOEw16MvUYxiPlFqyIqMdA/qAJbbIbCAOc+Z8FD0sC1EXCXFv07npGwWZNA86w4mOV1WoZPakAxQ8jWYdGWwC3WtJkTOXBTtgHypYbx7oRBB1OdJyLJDcCLB9lte7gjRUtzi/xsCaq8JtYEgNCDQ8OBhYPZy/glmxVH4kTSnx7V+Xm5T/WHOOuQ98zDx0kWgZ7Cwp7+NCgAgTk0uNew4mB6kghlUszX6T6LnbTDweMiQu9VDngXRAaReV2pJfDi1+9Yvi4WL0z/IqEWU0WSRF+H7W6cgJkRUIaGS+q/K8N2UmNW0D2TiMKYqP+u/n0PdncWu7VEpzy3+iHCCQroswG2lyK6JmktyZXvaV3RUECePdBt7ZITCHZRa/abS28rKqwqcQKB5Rr3hPiRTRAKOzXEMknEY1+Mbw/Els8w81skIXbxLqZbmQVhKyh7sbK2SCbUWFtdra0ZXXvNVzOthPCTJkFwYsJ+dhOJ9WlrEv4NWIoPMcxcckEPZDWrXSy3bTO5+DdMYhiz7A8erteRmR38HKARn4P3rYHY5X4Ti2Hisq4pNthbrEeKfOIbe9RyVKsn+DnJtmnklZigYrGAFAILiiqFRUiDJAeEcX/4AGL3i7VqP38lfhpMfDCmpu7oc2ITCBiVlnKAsb5Hu8Phuf/EDrPczBxPC6OcP5Agfc7JyQQ+rWEALpi3wHqQsqsMjfbQbjeR8p65ybYbJ+RRXxiAn2xUsO6KzVzayeUA6bKR7OO/o7jBPsfaxOvFRYsf9O4O/eRu9fc106O3V42KBEF5LT2jYr2Q/+aVKGa57+kTjJKQGUz2lbdPM+vSAAGWayhbNqPSaHUSe4Chszwf5luwPgHkBfSnCiWtFErxT0zi+2IS6QzyMzKCxOc1MSHjRMaSWgGxR02VZ0NaXGWRdq8mRX0xpxBWzhMVzrIdsxeyio/WlmhvbdMeJkZhVSTbn3bAm50YGR6qeWGzpilmaZaTJ3CeQ3BQY3N7S2xdchKKA74GEO8hkWWfE7sjYqy9Mb7/zadjYWYmFtZ34v2Pr8b8ZsQGjYKe7ujtHYjZu4txZ3pOw63v3p3VYFqKBNQaaZdJPoQagP+fO3tWAD7rF2sumgh8bNZZW4uHllJ0YdHV2magiYoLYJfcYfLmpNjRHe0ouRplCcUfChU+T4L3qDKXlxdU1LAvYHkRMxXbsvmLvL2lWZZqrLn9+1F9DBZyBMoeWzgx0Fe5XW9/zM7MxZ2paQF/AD6APzT/eT8GPF+7ekUsVVhp/OE9aUZcvnrNTQnljW0CZmkqEV/zzCYOkR+w8Jz7mHnN/qdxwdc5t2X/lzY7io1Y8jFweEuszFyD5DEUj0ePHlIupyGylYqGmLLO2T85A0u2dEVlxOdGlZeD7QGJyFM1O6ehIb710ktqVCyV2NbT2y2L0aWFBSl/Z6dnYnz/uIgL2xBVVjdkC8Xn3dp2UUuTqbOzO+bnFtV46O3rFmN0c8szLVgfzEMAJDOxh3gH2O2ch3Osvx/WtSmTnIvcHzd8PfCce8Xe4NpVFKsJbVXnxhZDu8vA+irkmw0Ri/g+cytEFi2xDmCVYrml0qBGDN97+KGH4pbsZzgfPXiYZ8r+ZE1fuXJF61gFeLGIgaQDYE1M4zVQaTDIHjXyFArkrg7VGKid2jvwou/QnAvOPdvBJDvVKg/WMfdblkvEMdS/KyvR291tH+jNDVmNQaZ68OTxOHjgUPzwlb9Rc4L9++Ybb0oBdfz4yTj38cdx9sy5+O53vyOg8tev/Sb+/b//Uymb33rrjThwYDweevhhDc/+zetvxTe/+aIISdevTeiedXf3ar8QF8kD1XjEx1/Wj8whWKkNdgWAQHFCQ+Wtt99Rg2F9kz0Pa9L55COPPKzP99Zbb+trNJilJtQabIxnn/miGo/vvf9hwL3IYdrkUuynl7/z7Xj7rbfjOjUIeZEs3bBta45HHjwplTrX/sEHH8b84nI8/Mgj8cRjj8fHF87FrTs31SAUu7rdSiD+nYOreR7EYg0ILfMPdL4nWaPk5dwDgE7tI2wKyww71rNsJCvNulfEaxqbnuO2O89MihFU3dQeLS2xsrLkHOwTaord+XzOq71GrOozwMn9VOOyNCI1y0RWUFbgC8Sn+Zw2Z8U6ivrUeZSVtvVnmMkpO1HlfFxfVVyluQwhi5qVWMPnYQ9DJmArQTRDbUGNKyBb8y5sLSs75IZKrcYChJU6hhk3mr3m+o66k/hHTeGczva0zidsKctzIFej7pEtCEqcSpOa6FgB1gOJahYWlZ3yh5ITu641eY8cyrMuTAyj8TYzR15ikto/eT1UQF1YRxMbnHvvBV6zbst8IlWQ+ZrEDRPiCmGqSJKs4mm0kq7kuwJ7mZtS7iX7zUos1KaQOyqq+9iDNCAB6bE+Q6myb9+o4gxxCCtXbKZFxOzujluTk1pzYyMj8dBDD8T7770TwwN98e3vvBAT58/E5vJ8jI8OxfnzHxsc3DceZ86clYUfTgNiaHMdzKvr7IpFQPhqNQ4eOhC3bk3G6sZGDO0/FBMTUzE1dTcGBvfFxK07cfbji9p/KPhls1qpqNk8OjoQX33+6Th6+GCsLs7G7Zs3NESXeL20thW3Z+Zl/dTUAgFguVabigxKo2bDawNLSJ4rOZTsPqmlGZxNLVp1XZ3PlLVhm1E3j/U8y2wJzYbjf0VJnTniztZW9HR3iqR4F1Vpq0l/vJbmDZZB2uxPmiDYULnZsamcjtfFpskpuZtv2RAgJ087bc4T7UuUWswDIV5sbSpeFplTzcrJOu8GvU9nW6sGbrMnkgwFMUizmWhWllzZpMC9jYrdmSwuAHa/v9eWeW/dnbVNDTBXHp+frygy6lRN9flwLf78M+RA59OlEsli+9M7G/8EXshrqf9G1sd78/f6xsTe3D1jMH9ng1LqgRJDk6SVeVrej/rXya+5fvAUTNSGxP+NDWzkja0oV9NztOIgZ5SmvbLUjAXAT7KXmm/gPBBRCmlPda8sl1NJjgrI61tq80Kwy6Yet3mjKMCoJ5RvyfHBVlOofe7OzQoryuuUopZaSxiC70fWgYJ7Gjkj16366uyIK1euqi7ApSaJPGBYeZbx9wiKf6wLN9k7S8JeyQ1PHD/xWaPin6zwz77we38HHh4YKkmNh8wyp4FDIxUVGhZWA2oYeG31xcL8ghIAQBYOEL4Gc46DXl1OpL5I/AqwTcIFMH/yxAM6EClQ5AlJJ35jTfLXBxn+uLoS165fF0vi/vtPaPPTOZybnY3x/ftVDKHymJi8aZ97bFuME8oHUjZI1R3Jo2JrO0aHhqVUeO93v9MQzvFDB1X80vzg4OQPIPnI0IgCCb7iJIXMorhw8YIOeHsJN8h6CgCKId03JycV0JCM/u6DD8SyGhsfE8glD/kGmOIUpk44YaNcu8rn2hD4gEWE/V7t/8k1c50kvxQiABF4BmswYUOj7EB4HYKSBhB2d0VHpwtJ3s8zIFZV6PuWO+HE35H/BhzhJsEGnZ6a1n3kWsyqt5znAAAgAElEQVRkMjPRRbqTfQFk5cby3yTIYlUUhiGsIQ3+BkAsLFr57TU3qRAjSQRc4Vnjbc0fEh+KS1hDklZjbSPWjb1O+SO7Gdl5OWmiUFUjR3JrD2yjKCDxEfjL8G88iUdHtO44WCg8sLUhsed1aXJxCADqYAfBAce6hgFCYi37naoLCkm3GRpX2KeAQ7KAaGwQmMM6l28uDbKisGEuSYVZHmWwUg4f4/pVuIjxxmu4oLJKxEPy8utidn+KUMEg/ydJ3fqSMqrC9y5o6ifyk2w2lEFhKtzKNWTzgWsCtOHeqhmZMy7qZPG8V7Ij6pOKBCM/keDUFXaAjgbHiuwTpqa84K1aEKsnbCVAUcj9Y9CcDn0VmBX5pLPOeaa8VtrUkHRwz1SEFtshijuz94oPerEsYg0R03KuQ42Ra36MVBNmuC3po/C+YvXlvSpNJKw3eEbLays11YgGG3r0hq6NZwpIaAsCGKUG7hLATZk7z44mJ58JpqB/xsP/WF80e9kjTiKRJdvOxgmOlSMkZ9ngyqKcr8lOzZ2T2nMT46jsMRq3xAzPJdktCimi+YAACiT/MEOJy91d3XHr9mRhkWBHsC2VB03ckeER3Ter5wyccP36WvFRFtBX2FFSpdRZoNUrKlQeFF9bFdgoRJBpr+TAzWKVU0B7NV7K/UiWbq5PniFWBTAJrdhyTHQjrSh2xK7ytUk1p+u16oHf5XOyt3cbFWWl72lUpBoj9wExkjOE8y7BE/mqt7bqtQW0lWam44GBLjeK7J9MfErQ1kWDWTjumHiYNvuG382mOK+hZ7a6WgbaNkqdJGAyL73ETQFYNQsl2wHKO7XGagNscaMi94HUHGVP1McB/p0FiW0pfIM8MwgrwcJ+3pMtZcGSxbHufxk4D0DOWQtwwe/rHG3AQmTNfv19vbG4tBJPfu6JuHb9aty4MRk93Qydx96sMb73vW+L+X3l8hVdz8wMFhbbApKZvUGxe3PyVqAwxAIJ2xMsYtqbG9So+OazT0V1YyOuTs7EhcmZuDGzGETrjs7OGB4ejdm7SzF5ZzoG+nuKgqJXigrOa1SQaozv2GpJzM2LF3U+kZ+wpilwOLMpLIhtFy5edMNli3zAzQyKMBpPnGOQH6yoYCbGopoi3PPr19NezHZe4/tQCjapCcEeR1HhM4jmLexSwCM3UxcX53WuAUI/+ugjen9iMOchhIIzH36kQmh8/IAaFFhc3rp1Jx5/4nEpdqambkdfT6+YYNevX1PBduLkCVm3TEzccnNILOhibQapYcOqVK4p2Wu2gysznKSqbFJjY3hkOG5O3FReSuOKdcCaBdQmngMoGsxZEsjB7gaEsn+5vf8BDNky2s/b27GyArOZe8+g9fkyA8DnRX2eKws/AWFVNTuIxd94kWHafyOrCO4bxBTyG+x4KHU3aJrsVGNkdCTmlxdjoG9Aags+M6pWfpb8mlxxdpaGGxZ7qJFpbG8qv1xcXo2+3n49c+WpU3e0pmma8BkA5AFXsREiB3ND3Uoonh0AFHuWvccz59+eXWCLMp1PPaxZPOzbxdqlQaAhxyhsIZhAdmG4fLtzR2ynUA4RDwG6sCcBrOeZzM1jb8mg1FXltdhfihG+saHP6iH2nmPH+pqenlGej3Uq/81nWl5d1kBtrlXK3KK4SJKIyQZdtTNUJIho1P3BXoXYZjLCSkzdvqNh2qjSRoYG4sPTZ+Pf/ds/iavXrsa5cx/F5z//eeX2/+W//CCOHz8YX3jyyfjzP/+rGBzsjW9+86X427/9W+0xao/Oztb4r//1lRgd7YkXv/HN+L//nx/G9uZKfPvll+P99z/QUHE1JpgbtbUda+tbcey+I1I7vfHGm6obpGYruS/373Of+1wcOXI4XvnRK7FVNVFF+aIGb29obxFj3377Ha0xwECaFLwO6o0nHntMtRP7fnR0WM9eSnPsJ1ta48DBg7W9btux7ejt64mF+VnVAjRp+vsGYmenMd57/30pwT/3xBPx0CMPxvbOps6XjOHsFysqHcO5fshHPA9iGTUBz12xqtjA6HwLe27LbqYJlQHAvwllMNBpZrpOslWTFccG7NIOKWe5ycZWUi7n0Hme1jcl7EnOecb/W6QWUx3Q0mJiXYvtWNOOis9Ty11lLwS71jmLBqOXOUap2nCzk0HaqBw8M2J9a0P1LmuR50ukqDRiAVLoDFUP6OZ9pJQRcY+94DoHZZxm/zQ2SuFHHsnzYx2nkkjEFAFl5oZRA87MTCs3TcDQuYQVwIDNQ0NDZfYgzR03NKiNOJdcT0FmcT6qukvqmWJfVdSbrEUasKw/iCJ8BpHtZJdI3U8TvRCukgQlFTpzFm39RHylbv9EbVCaSZkPp9LW+ZlnnCi/gKhQ7HVERKJGQLkCxrAJac+NE35fipuiCCfrwOpHJJZyX6wU3FCDrrOzI86d+1jzlI4cPay4CLEArAH1LecU5CFm3SwszovgyIyKK5cvaj7Q9//1d6JxZT7WFu9Ge1drnH7nbdUO+w4eio9On9a97+7rVoMURQprpq25Le7cvBU9ygMG4+qVyzE4PBydgyMxMTkVd6apHTvi7sJyfPThOTW0UFTwLAXua65EJUaG+qWqOHrscDS3NsXM9RtSTV2buB1Lq9uxsrkTOw2VWFxa1T1QPUCN1dqhodycY40NxCqfc8rRFO/Z36h2PIePpgHxiL0pq5qSD/NcZM+4s107u2XPBqO81Mo0aIYH+9UQygHAYBLs/yRMca95ffAh7OawsTI3ryE6u+xIAZmAc5QzxHUP8dF5pex4UcG3tOh+8yHIO/h9mg4oUVQzlUYAc4FsWetGRwuz63o7pc5kXd+dX4i5+YVorDTHquq1it67Phf4p9KETxbqvpX3Lt655vx/Pcif/66RrYpqqL6mrv/5f47wk3tsbxNh797bm7PXx5D8Xn1OviddL/dkF2HIa69vPGTTPvOpbDzkz+Rr1tcR2ShJpVbeLxctVvyzz4mPKBI0O1LuHA62nIusYxO63KCU/XJR7PFjEBSEk7VgC72mxoFJiVb0cTYplmI/LWzBNU3GzLxuZqvyh1ybvKxWr4D1ra/F7NRMzMzMRiezwLg8SH8QYAs5RiqNUrOxYjw3kjNwSyRA6hqap8ycwFGA96dWoTbH/pXmCGt//4H9yo2xU/VabRDZiYbsZ4qKe63cz772e30HTnT1qNDTkMelRRcOkoxbxotXdnYTxVTubPdAzpKkytu8FAokpxSBHuK2EZUWWxloUGNRVYCVcYjh28wfWAwkgGOjIypMSaIo5EkwOAgFnCDhqzaoay5AftUsOrzsYW+ogOrqkh0U4BmdRRWFHV1x5NAhFQBYYHR0d8YSSVZDg3wnQRhJQinYsHMikNEk2GX3m2FPYU0H9s7tOwpkzLNg4Dd+w8xd4BBuaW1T4kpyQjIHuM6hngkBHVISofT+BEAT45HDuABXJEuaabG+Lm9L1Aj8DgEQBQiBXMN1Ojs9a0JJB8OqWsXmQV6cTH8xU3YAKjrVgKCIJcFurniYJ2AqCSCsb8ltxVYy2Mr7GPQnUBvIUzMFT9gtg055yCXbylZVXgsAJfqZaoOeNQCr1A3yLl5R4BbLvIwYss1OYdDKk9f/nYezvMpLMmuPUuyfzIgy05hGDUlyvwplCmQPTG2PmdlZAZ4kM9zb4yeOx0cfflTssyiOAUG2lKQtLixo/dNsSesozxYw05F7D2PXjQc30GjMLS4vyxuUZyVcvgDnYhbx2TiofOaq6OLeCRwtzAoSb98w2xvc80/aLu3tV6Q1UzKhxfTYZX8kCJgNiVSocG9rSRL3XgOSPXg7n69B3bTJcAPLcn03XQQKlueW15xpTKop9PWC5KqB1rA7gB0wUkCoPNo9MI+iF9UAYJqYmXis7mxpn4rdJ5aZfZthBqWtVl6zrEDaWsXMwc6F34HRq2L3XjIQrI46O1SsUajmvRO7vPy81nppLPB5SWizqce1y1aqzB6p2YiUYc/peQ6ow8sQv1CEyKKpPGtLxCkU3LDYZPglDUTJ2jfEauZ+UCBaWWAWnRItyf49FBl2OVYpbp7YdxlWFxfH/vAg5TVb6Ghonu11uDYKFK5dtmUMLN7e0r6lcOe5ExP5Gp+VdQ1gS1zV2laCWNj4AHswBgvwZdmsAe4kBe0O4947o8LMQKkjgpkbAzofzLbykNcUdGWTSnYpmini2TJmOpVh2n19AnUMgnod6+dqA3t3rbPcqDBgyt/EAdaaLEtqe6Is5foNmhs7NzAAfZv9nGlU8J7cY9mgFGYn98JgnJlB2KzQ0OK6WYN4uRNbaNDkjJvdeKHs1w0IEulScFLe8/kBsHlmgI8k77B/1Jyss50TeFkYP5qRQONIDSQPonQMg229VvOX3QVMdguy+uKpvhirV5HsLVBqcaJOseUQ4SYFaw/WU6qssL/I5hyfR973q8uyiwMwffGFr8ebb74RV69OREsLyhDWOoqDfSp6TaJojcnbt2Vtwj6jWB4bG5akWoqKotrrJLavLcVIW8QXHj4RlWo1phfX4sbsUlyYmI5tWZq0x759B2JmbjGuTzDcuTvuzs8pD8BfHiAWlREgFWcKljzEIWZkaV8WSwQBKBrW3Cp2uJqTzI3QWrVfMmA0zxNg+ezZc9pXsPhRiQBa8UxoHuyurxZ5bFtVyMDuttqAQDVvafhXXJixxmn4EFvbWlvi5MkTAh0Ac1gfZ8+eFTuT2Hnq0cdiYWFJ4DLr5eixY2LmUxjBkn/0kYfF2AYMI4YdPHhIz4whl6hfAbsAujgraQ5wdnM9tm6xbVySJjzM07YF5HTM4CL/kp0ouUUB4j2zpoAPrbaG4vOyZwS6rK7GE4+fEmDNnqb4w4t/bdVgrPe61XN63dI4dNPeqjdbDbqA5Rqee/ZZzahYgknX3hb9gwPaH51t7bIemp2aimpjo7yFBWIyxLQ0hohfvEdnOwrc1Vhdsf88+VVPL8q6zRgZG4mFJeKdWebEUJTBzABhT6P6JVcGSJeV5+Zm9Pb2x41r19XU436Q/2Crwefi2QEakU8TxzijaNQRE1lLx+47JgXx1PSMVW+A0mU4ryziYaF2YlXKvBia070iw3A/xAQvDQXWJ+/H17BQotgmjvFMiedStBTgmPVBTgjIxLrgXDl89EhNhc3aYy8Qn5grRr7N36orCqgqALf4TvMsWRO8x9zMrID0hp1tzXj70lNPxW/f+I3u12OPnYqbNyekVHjppZfi0qUL8d7vzsZ3X/6mmkGoKh499aiA/t+9935cunQ5vvdHL8UHpz+I9393Ib798lcFGv71D38ef/Znfxq/+MWrcfqjC8XOwecvLGEaddQ2v/rVP2i2Ag1g2/vgS82w7MdjbGw0fvazn2udVmWRy2doVB6i2TOVivJ9e8RDvLGXPDl9t57HphqefE/3Qs1j/r0qoPjGjQmdmZrnt8D8AxoKS/Hlp78Y167diGvXJuL5Z5+X0vitd9/Vczt5//GoNDdqbRucMVufdYHnv5/ljuq5rAfZJyIoFBuUBJ5TiUDOpvwMJrUagVbrAdqI+ELdITKLCS35mUyUcrOS10c9BytHM7Sw9pI1XFuN7apYWXJTE4qtevDsQwZlu6kCOAr4qsY3zTRstdZsFcy+qgFlwGHFplHNvnLk8TXVRMTPJnJlz4kSYQgGOgBUmReVQ075bDQuW7jeVsD2VjUh33vvfe1pKeyoZ1FeFbUH10odWRJxqQz57IDt5BSp/DbYZ4s55TYtzR7avWH3gmxSkougqBArXjNiymDzJDHkrDUp3P3sAdr5eduRkXPbBQEAP/PUzEny/OZMIxYQazhLPANx94/rHqOL/DubLLsWeB7SrSeodUV8ZpHZ1kXvQ15bAETlFo3EIqvRlKcKZLcSiKxHzY3tTZ0DnA8XLpxX3j00PKimhKxTojEOHjqoGUtq4s7M6Awm3sL6hyRJo+Lb33w2FufuxMhwf+ysL8eFj89Jybr/yNF457dv6TWp4antK20tVvlt7MTdqRnFBGLehXNnoqunNwbH9sfZC1ejqbUrtqtNcXduKa5cvR69YABYAhZVIef4zs5GDPZ2x+hwn5Qc+/eNqobYrEa888778d6H56Kh0hHRyJlqaza5E2gOBXhMlLW/EatrK1JLZfNf66HMI2KfW53txmLuZ9ViyhVco7vmMemAXIrf78CebHMzOtvdaFZTfW1NTbgVzlzpYU3QI9+xcr8azcx0a7PNWm9fvwlYVTCgJdUXNGw0t0KOEFj/2Zp6bY35pk2y+qPy4P1y3hWfifpGA5IZtE7NSIOUnGcddXtDNDfyO31ltuRCNMmNAntb11P3+mPyV6qrd3/iU358FyMpZJ+sUfk762bXRyZJZU2QpM1PNCrufUm19/C3d68kre7q3zNfIvP2/55Gxd78fW+zJYlMvHb+OxuP9Z+jvmFT/1FqGA9Ktbr7ZHzCVktSU0MeGxgslmQd+qhuQLG2XN9SmzqnKzMwyx1JW2w3vryW1GhAiaEmuOsPN0JtyWSyIoRUEyaz8OQO8zO4lPA5RaagSUwu39ys2ZOQoghbPE/OAfnIJRF020qNtDSTa4M2VVWkP1RZ5FgTE5NSnoI/3Z2bV94PkZn7T3w5ohkVt6xeg+DY3aU9AIb7WaPiUzbLZ1/+/b0D9yNdZ3GX9qRZwUViVTUbXd5w2FZIJu9DEDA9u5AkifbWtN+vAMzCTgVw5jDhD8mhN3SrQDSYLhTjbGiSbBgMHEq3b0/qUOK/Gf4EO37qzrTk2hSHJNh8zZJjZI1mjaV8VCyjtlYNtGLzA/jPzM7E3MJ8jB/YrwE0U9NTlr4WFheDMEnEVpaWFbhIWHgPkq2dqpm8BE0NheztVQLX1oI0q0ns46UVZPx9OhCRVXfi91rASwItbAruK0AGhRyzOiicMlADqpPAEvj4LCT5sNauXb2mxgcJGl1hgbQk5Ur6zFrlNaamZorHpO1nUkLL81IRuboidhNAKT8vFYQAYgNeObxMbLXCajVA65PZw2b9PfnvVczkqh1+GqJlhQMFwtoq8wNQLuCVjsepQXrAMApoMWIKE8Z+sS5iJN3VACEASxoGHq69O7sCBpqZStzrtKdJ4FKJl6TQtnmiG69BX6Xw4nppUjHcXGCA/Hfx5nRBSYIIeMNr5+C6LLJylgsFC3shG09qApXPz2uxZ7KxImuqUtzVH/oAXirKCxCS9z+BcicENR50LQ3Zq+jMRli5fTXGdf5Cvl5aSunZCvD1K7EOxF5L1jYgrpJRf1/pZFFcqHEoALyiZ0MimgzxXAe66hwkVq6/PjFCpcPvECdQUzkhsbSYvwG7PLsjGzk53NugPIUve5NET8Np09O2zGFIpp2Zo1Y2oNIACPZ1GJzy0nbBTPKb4LXmdggLRr1h4DZBrPw7B32a4e4ZEbIUoaCjsbLtgot9CLifzEjvOxQMthBFFg4YRWJi2zZbqInFy4yKEtMAWvJZZWNzF5C3FZKGzg6hjrur2CeWU2HT5nXwHEngPQj8k81AnlvaGsiHszQa3IDwMEw+t6XivE76q2+VGRDEUifgBrCSCVo/BFt31utqzzDtki3aq182TjsCf2kwA3pJdVCafAJMBLbbQ9cNWMeTtIDiGecQYw2d1udj3bnhkom85hwVRmF9847Gsjym5+cFrGQczCI6m3z+RMV/tDS0aFTw+4ADykGLvZ3susp7KSnW7I5dtQOfiWbU4cNH5HPK55ZFX/F6B/wUEFOaikqC6b8V+xri1P4DB9XA0wDy0oRSfOU8phlCQ6OAIsl+JU77s/vZeqigmbP1ipu0HBRYDOMPeyaBCbsDoeV7nc3YArBkvFGxAqBQm9Xh4oT/xvIANZHPq4pURjwbg1bFDmp7U00K5xA02Kqxb9+IfnZqajYGBmCBhoAfqRobG6VywHKFYdaAWwB6PAcAUhXeADz4rRP/draiur4SJ/YPxrHx4VhdXIi1rWpcQlExvRSb2FZ2MW9qWPts9i6sdOwiYZz3ic3EwGeAYVhQU1PTcWD/AQGQ2MrIekrs97Q28ABLzjfuTcZSrAz1I4225QQsIS4C6NgyzBYbrMVUvwJu8fl8Nrk5lSoe7fVNzjY/3wS1WPdcO8sD9hZAtJlwDXH16vX40hf/IN56+z3lOygwJ25gH9IoRdnBw9gqbcTly5fi2JEjUlXcnLypNUscwpaM2Ib6lfuByjJVlCIGwDYVU9K5Fc9UjbXih0/spbFBDgZYjo+01ZMdymVkHbq1pdyLfb607L1i+zvDlX/4zDOyF2JPXb16NT786EyNMFA790osypxHhW4539sY6r7le87/n3/++fjRX/9Q184ep6jk/qu5VK06J2wDVG2QsgkCELlMWtEAABEjmxoB31dK87JJw9N3thlOjR1YU9y8xSBtFB9LMTw8YPullpaYnb0bgwN9iu/8N3kUZ7CGqx85HDcmUHAxMLVX1kxLy6uxf3xM64afY80TM8RsB/Ats0L4PACjFPLYEdmijNlbnpUB0Mc1YPmVbOq0mwH8Y83QUONZsw4d2wwgANZzfrFfOBuHBof1XPMZanZYa7ttOddWJT8AvCd+qXG6sSULLa5Js07aWzQPhbgHAMEa45zc3uS8tJ3I6vJyjI4Mx77h4bj/5Il4843fwtGO57/ybPzgBz/Ss3nqC0/Eq7/8lfI9ZlQQ0376s5/Hqcce0738P/7P/xSff+KxOHXq4fjRKz+OgYHeOPXYqVhaWJZi6LXXfhOXLhfbNVQR2AZVGuPo0cO6Fwzntk1rWt16b1I/sHZR7/b29vnMkmWS1bcJ2kPG4kzPwaECBKs7cfDAfqmzsLrd3NqIzQ1bX6AGI378qz/+4/jlq68qDlmp5DynUmmI5577w8Cl/e9+8aqsxZ78/JO6r6+99ppqHGqyZAbzmikl1EwG5nCUmXHKY8Sidk0gpnWx6eAMUQ6ForzNTc9UPEilX1TZmSMS33kG2QCQUrvEBM0jXNuQQoL1RH7EPRGIz7DpotgiVxH5ifWrNUyDgv/7nuTe1uuW3DbzYqlrFY4BCv05sybiZxIUlw1Ima0IqImdluuhhmipMJeCWRUeKp7/57wlxlLHKcg2Ngp44s/r//h6sZSz4ki2N8Twwszl+n2OOkeHWEYTKodie//t2vHq80Q1Dhw4KNUFtU9eP7kIoJZIKeXeEpOc8xrc1EzA4mvP6xLzyfeo3zgn1YRgBuPCfK1myTwuzy5+hrXN3iW+ECv0mnUqVv4zraZSBUOjgT+Ah/pemRvG15Rz16xXsUx1oyxzOM3r2nSuu5u/JSmIcx5S5bIssagDsWviNSCvjYwO65yjCY7KiXOqr68nJm/ejM11kydpFE9P3YkD+0fjmS8+Fu+++Xqceuhk9PV0RlNbS9yZmIyeoeH41d/9Uvdn37hVL5AiGipN0dzYHDubW1LvH9g3phkZbe0dMTx+ID46eym2ojl2ohKr61jH7YigyDwJqxFX5b/fjOKzGbV1azRWt6Knoz0OHToY/SNjMTF5O37xD/8YbV39sblDk6FdtTd7knMBBjhYDOdBpRGbLNtI89rJds8zn/XtJrS/x0w7GnlsGvYue2d1Fdsvmoft2oOcGdQTfH8Zm1RmBFYaFfNZy8RmSDdqEipnNBDMn00RdNwMJ29Azcfreh6m61LfAxMAeb6oHRLEzj1H/sezBRcA6+G1OBuJNRBToQlSwmreQI4+1CxDrrs15qkvmNNWcgftCbP00uSptD+zyt2jsagjBu7+xK7iqL7uz/2WP5exKdduPXBf3xTw9dRx7QoQ8EmcIF/V81pqNXmp5euvbW8DIvfy3t/h55LMkd/LBkR9Xa/6qhDvsgmZdVo2Lu51PfUxLGul3Qt30xmCK2cKOTY5FiSmXMeq6SAl9/Z4pg8Yk/AEmuN2kOC8IAcXBlRwIymGNLvWROisp4kBECOIF67HmG/pRoWcPko9XG/xrZl5ZV4mlvjsOztHOCZLASfikWdz8cxFGlLscm7HGr/vvqPlHMBSCvVIg9xTIOHQYGM9Q3oix0R9yzqXgwruHpt2Gjl69MhnjYr6hf7Zv///cQeOIzWU16sHBpIYkDBrgE2jWVIaOlOGHpvpZy9zgoUb41Un5WKsWnpJEqJuY5OHgZGYs5k1GIzGQnurwHgN3mtzsXP/yfuVfOOvymyMRx55UMnZ6dMfqtDBBgHGEbZLsPsUGAubB8mk7FQ6O2W5JI9YBbFmFQcTN29qwx+77z4lUsizEiROWx9/3mUdksi3+R0srmA40wzBT3jf6JgKT2Z6wJYCnIAhhm8vBQogHQVbdkpVUO9sq2HCwC3u9YGDB8QkxMNc0rFiG0Mzg3tI04ZDnsHlsP9J5PFrdkKLrcOcDnP8sf3snLxJeQJDtjCilKSXBos80H0aWR5dElVuIECNBg0VtqKT+F2pdR6m6mIXayiCNkl32nqIGSxQ3vI6/hBo/ewXynDRudi//4BAAzG3sUIpqopk26gYEsDldZbzKBJsJPDDCGGdpIem2R8UMSRBZlG1NJOoMXxyUGtPAww3N+PW5O0YHxuNzvYOMfo0Y4PkjXsg6ypks1tSVZAAAUQIXAcgxwO5FCNimwHmlhSGJIv3tvWWCxwOLLPUDZolQ0WgoRgAuzMBeP1y0/xX3QyF+sR9b9TZm/jsJjd1AwRLoqLUpf7fBZzOxExNv0w2amBymeFQAEU+twtr5P1FXVMuSp+7eEiTYugKMkkqQ9qS7cZrkFiyStIyiQNb0l/uP/7XJNTypLWigefA12nyiDFWGnKyKJANjln36bsvaxwKT4GABiW5HoGjZWA2a4V9IwYe6hrkzgBnO9uKe2qqlEYWQCrXz+A3/zEjX3u9WKCxHjraaOBVleR4Fo+L7FwXuV+JmXw910w2cHgNYlcO8tYQRXnpW7Vg30yc7az4UuG2taW9Rlxyk4zGgRuSunN1hZzA8vEZ9z8AACAASURBVFqTalfhk1Qi7f8y0FoDDcv7Mk+7jI03C19NBYPcnkPRpIYN5whgQcZmNbfEotodXJ3Fhp9HkVpjo1AaNawvgBzWGGAWXweoqgcdZG9C0VPYSCgA0m+e+AmAOXlrUqApfzb1+ygPzIYRgCvmla0PtGYLu3BgYFBxAJudlL/XmnvFAqk+Ma9vcvAciDuA01Yw1StHHJ+JwUqaiQ+lGcYPArITIyl2WRcUU3wuFHtmvzVEY6VBTRu1jAXyWv1CvMLiDpY0lh6sfTd3rFYQEACzu2l3eDx7NG3gUmXBvVpanveckaI0MYBmBm3eB+5lekLn+kJplOyhXWYaIJBtzAxg0vj2TAxiKkBODm23QtJ2FN47NJyXtU+WVpaCmoEzHc9h1gTzEQBPsDRcwLqvF0soWyvlzBburxqIOwyJ3DQ7u/jna84Tszw21qOztTmattZioLs1Hj55LBqqW3F3fjGu3ZqOq7fmYj2ao62rN/r6B8T0R03Q3tEp1iBsSQY3w8SmuAZwmJmekTqGs5qzPpUMtq+D9clnxBO+UeoGN9KsarIVowfhqhGleSJNKvhz3XM/ZXlUYoDAhZaWWF21+oB7kMOnKe7yzPdg8nYpCHW2NAJAsF5skcbrM+z5qS88GRcuXorJm7e8JqdntX9m7s7F0MioiBOXLlyIvp7uePDB+8UmY61SWKIK4HOI7IHVFcPNe2wfpBwTKy8Vt7t7jmtW/JV6sU2gxczcnM559hE2QwzpBbzl+aHSoDhjvQDsSw8oBSBWNVsaPMjfFK/sNxWQyk9adJ2sA6vUzKZTdCN3LcpQ3f9CXuC+fuWrX4kf/OUPys83i3VMXsr6Yj7CHCqm0jAdGhgUmBkNBkdZkwC3lSbyBOYSOffFjgc1RTU2o7unI7q7+wVGpnWCbLJoLJBTiV1uEMds8x2pi/kDqUfzP7BlRanQiuVNixoHIhaUpruJQ1iymTmKShn7E+75CgNXYYSLCcj+qmiGAg0NnhnXK4vNoqSzoq9RwBYNDfJIFMmA6j7fK7G2viLbKNb4wt3F6OzqEVEJ4AyVAbM7VhdWorOtKzarW7GytRodPZ2yg2qKpqhuYqnj5txWbMfmzmZUWppiB79qWf5w5gDUY9/Sq9xwdWkx9u/bJ8DxqSc/r3vxd7/4ZfybP/me4jls9n1jo3H/Aw/EO+++H0sL8/Gtb38r/v7vfxnXrl2L//Af/qd4551346MzZ+JLX/yiwMrf/e49+cv/8ff/lXKUq9duRGsbfufYC3WUOXYMtjaYMT/vZqVsFAtoLKvbci8vXDwvJR3NJ+KSrEliOx566CE1wk5/8KGs6gSmcI4D6jVX4qtf+cM4e+asrO5aWiFS2LrRyoNWNSp+9vOfx50702rcyFJqgz0V8QdPfUFN8HfefTcunL8ocOf5557Vuv3ow9OxKJIWr2Uyg+1/nYc5ZtumiqaygMvCDM1B06kI4Jxhz3KeJMFLnvACw0Pr1EoF59Wcc1jJ7WyZAIEyXGxq5Ww5lDntYZ0rpO99KqA8lLv4vYscUE/0MUhJvEzVd+bROhfZH4WRq2YD9mM0ZpoAa1v1OdgDxHHPTjB4l/WWlCXF/oa1SP1G7keMk1oDEGljS4OOU9ksILXB95bmuVWz1M+tItGJxb6JutgxiEYx+SJnTo1cpefuGW4igkU1jh+/TzaB9Y0KauhUltbPW3P+em8+OO/nHNbuBQaCsY+7W2L0Lsktz34+C/EqLatyqLZh3ZwpQj5ZapNCTOPaybVNiKRZ4eYGIJ4IKtSm5TklsSHXElfv2Tq7jf4sOaQQVPxcVZ0OpkGjormxSf/N58FmmliF0ozYANkBhdXy4oJmcmCleO3y5Th0cF88+/Rj8dqv/j4ewN7twLhnMHZ2ax7CRx+dk0IGYtzs9LTmPrW0t6p+RLnBM+OMuHjurFRnQ8NjcebcpVjZqEZre0/MLa/F7DxNISvKwEY4k5lf09pciZGBvujt6ogWCS5ZD13Ri31RU3O89sZb0dDSHsvrKKBC8/O4mcrr8EnifAdTaGnVPiB+QxrlLOGZWWXTUPIK1880CdlDiglVW9RQr+ncLv8tILrMsiAOCw8SY9znOtfd09WpWR+QS8njOHdL5aSYB2c97c5EoCFutLVEF7beLbaw4j23t2yTzYu7MeV4iLLWakuTzmTtzEzVMj9jhvMIyzop8quq05Iwwz5HlQsJAhInP2fQOpXbu24C9bn+3hpcn2fPjInMkfVe95g/ca/X4Gu7tciua0X+/t5GwN5GQf17fqLJsefNskmb113/7fprVZwtVrX1r7e3ubD397O5wd/ar6VGrL/evfeH10jMoxaTiuU2+B3PGmLfMnFTyi83jq2+t4qdtdLKzNWikshmgpW7xSa6BId0Bqm0mgCn/GILu8t2NdayRqDuEq4lwiGGk7b523VycP2a9t6zs3N2E+CcEF6GWhpCp/NaXWOx5bRF9a7FNPUD6r/bt1Bq92lfkIsR/4nfUrHS3NjaikcfeUSNCs09W1+PaQieO9siZnymqPi03fXZ139v7wCNCg4YHQLyzuyWPxpJJ1+X7UaNiYmUsEXJNptR4HeZE8AwRHc7nZxyEJIE0smkeDl5/0m93uVLlxVoSOZSaqXhZWVoK+cEbKDOLoo2g8sUjppFUQ4EFYRNFSWP7tpWNXyXoYYp+b07yzDR5jh86JCCz9Xr1/TzJG00KrA1SLYM18XAMV4LJissDFgoJIwkDARBD8OuxvLSopoONEoATHg9hvqq2QJ7AQBbg6ucmPNeBMqjR45qkBcsb3kRLyxpYB+fLe02BocGJTMliHI/+fx8bgCFBDr4LNxP3hfWBjYQ+PcStLIQEiCFXVNTRQlKHgpip5TCx4eCmRJ8ncJAxWxa+RQlhRgudYPN0vaHa+D9MrHPw0/AWxlgSQAF3CX5IrEChGNtZFNLQCsMdw1rN5hcG/Qo2bkBCdLaZJiktzX3qBBTtVYoJuWxLuCDoZPYDeDb2yyfeVtTzMXBcQ8hpfOtRloBKbGy4T3EzIkdASIkith4SGVRwEDJ8cvAVx9QBrdbNGtlXZ9dXXRZPlj+lyymVIaYDYbth4eyW/5JQmPQ+JPJQv0Qr3umSLVio75JoYO/rlGwt0lRz3RyowIA116K/KzufWlOULDxuSxnLyoLWc7sgpaZaORANseFMqOiNoDbqht95jL8kVfL9ZpKhJS2U9yRtPJ9/U4FFRZqAJi1VlClFRJJS64NElU+BdLk/JwUXE6YdmqAL3t0a8tNU37eoI8HCxKHSI6SFcLXrSAyQ4K9z2eRDLT8UdFZAEL2DEoox5jdhC/VUPXANr8uMID3LGx19iGJDYmMm3hmwNUniUqCJZV2Q9K/4yZZ3mOrU+qaVqWYh5mUDRODzf4ctj6CB+rEUewnGgGSWKNaQDpt1r3YVKWYoHAAGKMvon0hgBuPW4OfBkndNNlN7A1+1xJYqV0Y7u59gLUeSRmgsK6r/G7ei0yAbX3hM0fqiB2G3HvGAeopsedLIyobi973fi4GhJORZwUItlOsQwBG789dS7b65FtJc2lu5N4lEU1FhZUX/swGOhwTAC/4w/POQEZCTNygYc2ZRHwVqIsNX5lfIYs+hq+VeTOaM7FTFZjC+gccUyHKALfyGdX4477K4ouBcpZOE281sJaYVVROaSOxvrGiwjKbNzlgOAuvZFnJ87oAQyZk0vgoTE9aKVr7u4VcxluK3p7urtpZQHEgL/YyiDnViBShNN809LjF7Nux0SGfbaurKv41k6VqUEUKDJiMsiq0RR/zbrgumvr8mxxF6jkx4a3owBpwZKA3qutL0RKb8Qefeyw2N1Y0k+HclesxObMem43N0dLZFT19/WqeoY7E/51mKg0XzmuUD/YBNzAGkMEZC/hhVjJezJ060zUEeM2MLSkji3KNaybP4ro4g3RGq7lhT3fmgvncrsT01EwZLG+LtQMH9ut1YPNzT4iFrCten/cGEOM9YR5ji8h7yCe3ipWQWdLENJpH/G0W83bQuOMeaj3SoG7i2hiGuyQbHoaOCnRcWtIMANRu5FIAHQlKa61qeHybSCNS8JQmY/0987wm7JY6Y3XDYB/rBoUQxRqxHyKKGhrNqBMWxWY3zd4xjPMfUF3Kut4efYtiLlVAVv16nWYsTqAzB7dyBqTSg/v95S9/OX70o1e0pthPo2NjmpEAcUT+7QuLBcD1swcMx/cfuw3iOAB9S0tbNDU0x9xde71j5VNpwXMZQgSElrGivJ1SzIFFyPXJ7gfgF0uqtjbdW85FPIqJLuRj/CGW8bNq/jUzMH2ugFPMyaiouYL6QOC4vJirsVzASNQ+EHLIpcnHs2kmRWAdyxmVCqAfnwkgntjLvcN6E4UN57ZIGY2h4diA5KyfuVly4apmcPDZsExjPge2pe0t7YH5+PzKQs1Hmhw3thpiZ5O40BitHW2x00SuUo2+rp64euWKng8AN6pIbPB4NuSZx48ekZoFJfb/+Gf/Lt74DQz27bj//vu1h37845/H17/+nACJV175WXzhyVMiQf31D38STzzxiGbHfHz+43jzjbfiueeeicHB/virH/xNHDu6P575w2fjwvlL0Vhp0TwajsjF5cVYXVuK0bERrb93331P81DUTBTgYlHeE088JuunV/7mJ7G17SZxe2k4cPFPP/0lrd23337bQHghH/E67OEnHn8szp47FzOztrXj3tII4vzqbG/XDIyJGxPK+1mTHe2dijc0cPh9hp1zjjK758bEpK7lmWee9pqbmtJesW+951KwRlknrH/UTDT8lNOI6MBsDj9r/pB/iMBWGlmA8QIaUd+vr+u1+D+vT8xmrXmWDHYcyaHxTLPMJ90EcL6Rf6xsrZrhWhQZxLE8i3XPS2OXn83/szd253lYJaWmCox17KXqclvXb46fNEOp4xTv2CtlZhI1rD5vmaPn/eTn7JOwziYG5W1hrOf7tFQMrjU2uAnN5/Qw7RU16vgcqFxEQoG41tOtfU6MznzK9r+lZmhsMJHv5qQAYX6ffco8MexCMp9ULK2RM3ZrinpLEkh3Gna+sqwYQQMC4IxcLPPGjMtJwOL9hB/A3pdLwlqxuHGtKTsm1nOTCQ4JpkPaM8u+2NaiHK2vgwouIYVMGZCeMZurX1nbqOWGuzUQlkI4NrBWq1JW8j183iHhHDpwQDHyytWrWh/Yc1FjDw8PqubbWF+VjSIEwetXLsUDJ4/Fl77waLz1+q9jZLA3Do6Pxptv/jae/fqLUixtrG3Gx+cvRP/ISHz4/nvR190RQyPDwgasMrkb9x09ElcvXVIecOjoffHBB+diu6E5Gpra48btqThz4ZruEetxC0tELG3Eou6Q9dNgX7cGVG+seQbIFhZJS2vxwblr0dzRGi2tHbG8wpwFKyGkZGpuFNGSHJK1xXxNclqxzIuPPnuR50IuqMZ/IT6C3aheI48qecLqMoPC07aN9ZVEPOdXkBebqUHKcGH2BEQGGvLUaJqDtbnlfUTuzXzASsWEIPPR9HdbC3Z37Z5DVVSiayvkAh5Ez/Nn/xLTIEKKHEMDpalBBAYIhyLNFGWn3lduC65BRfhSDtUiRYXn5pjkoDy2CBL2NglqcWl329RyiKzTMqeobwhkPrhb++wqHupe6hNuFnvB/L2Nifrf29uYqIH99T+059+f9jP1r5XNhvrrz8+QL7f353fzKRPAstlR/9n3frZ7vRYLgZjJ/iG/5gwjT98ueUvGURQ51DQ03pg/k8S1zJvYK4lhGJ9zPCV2ot5E3QmxiHjGa2AbzRnG77FniKXEXM4C8l2puQuxVIp4He7kOh1x5fJV7YN60m8qAvN6kjRCPlJPNCKvYs0TP7HcF8ahGrsluiArbm/F3OycsD4IDczbkQK9UpGSbmNzXU2WzxoV/8yi/+xbv5934HgXnmgrNbCI5JZGhTY3zKCFBUupJKtnFkOrOusACFgZsNFs/dQrRicb3R6WDUqszFiz5zdspWTqmOHphFhqjUZ70UkCLcAXJleZh7G6qsOIgKTBt5WKBlMbvHDXnSKWwgTgTpJGmNWNSBC79d6A1WafoPTYUtFqpsuGfD3p1sJ84ABXp76tvUhozViDwc9BBkMDNgbDupEZikGyvi4wBRCba7546aLuEyw3pFsA8wQxAw+rNe9oCgMCkQrSvh4VelTUNB74Oe4l6hIPq+XrnQqmfCYD4LszNLC2AuRHsitwAeZgkWzToAFAmF8AdDOgSZFJ4cHzFvBXLGEEhBaP13sdhAr0WwxaXRfLU40WyegMmoqx04AE1Q0Q2Gc0AQATYLvC8BMbfwM5XqdADA+Zo8ljJp4ANaNblu8V5pwY2iUp59lpGCSSdQ3eHdLzJOElCQZA4JAhsUaZwmvBzOjv69cgdYAfBsYB1vC6WfAAEGEvYssVN+NkLVCsKRIAS4BayX2pSGyP48MZgAbvb9hxCbopkSkZe8oNnSw4caoxwgrLyYe5WwOfQnwq36tvGJQiT0VSsTFyl6ImBhU72hPM9MwycQMo0XOkCC2M43qQXAVOAZxdJJtVVSsaKCrll2sgR5ZOOUi71qzwc80mEtegQ10KHoO5rN9smlGY2JLIhcxuouh7LBC+3CeB+vLq55oiehmmXjVjD/ZazRcVC5RMShnG1UqRinUH8cxJh1QWBZzmb8AhrpO3Qv7Me8oWp3wWJdOliNq1tinrFc/5Yl+TTT9+L38+VQCpTtKzKfeNvSSGU0tzjUmXyV9eZ7LOKHTZd/x8gvoZ87hvsrorqgEgnVQWJKvKoIqHf9GMY18lmOXZDoVNWJguDF3FXxbAgoaPZbFeE6wx9qaaIHXzUCz7NwM09wPfL24tto4rzMscgAtrWaqW0qiQcqOAI7Zt8L6SxVp5bsw2wWIP4Dj9+Y0fZKvN4Fs2HTLx9JrORsWmzjmpxUrxlvc+mxeZcPM6CZRY7dYlFoxs77IhoqYVViA0+je01tP+jvsEQMq5xfkjIEcDKgGoPQwRaxTA9Z0GBpEyJ6Ui9Y6Ktgo2NWbaCRjCXxVQQLMJrD7jHhEfExQX87zYymChk1ZUatBVt2SZoMJRe8z3xfM+srm067dKUZh2IJLYV2g4+edoqMPO9l734E9mXXG/aHylzB8gNyXW5B0AdgZIC8tNtjack706z4jl3C/OSq4N4JgEn9egEOaaUiWQqiuKcQFOKytiTGqYO+codkrtzWpUdLU0xsP3H4vFu3Pyiz5/9UZcv70YW5XWaGxp9/wYWFhSYLmB6v1tC420UCM3sF1TqwAf4gzDnrkWnjU/hyUS94TPm4CPbDXXyTdQdu7Tz5A78TUIE/N3F+LkyeO6nyg4RBJZWdb7jIx4wCSLDkBCftTFIpP1wh/OXtYJCgidVRBMOmBLbug8pzEhL3oYxS1ten3OSfaRlCkadkozG2saz+IaHx8TUMoeBACamLypeIoaQAMx26w4ZM3nsFXOAFnZ6cx0HOf1BIqg+mjviJm5Wa1X7lFTS7MKNf7wXuk5z0DvhYW78vn1TCiv8Wef/UMpQbjPsNABjx1fit1UsUzj9RxP3FDkZ7xOC1BcmrdPP/10/OynP6v9HMMPAdAzFqHSVS4Lu5Th1319agADFsnOQjGSJgqMVkgYkBWICZwjsEXNPhwcYJbXcszPMderX/t5bWVVzU81qtoYntwkNiiWLsRLgDjivuxLevu0ZyH0aOj84pLyL84QCDm3bhGX7Gev196wVz+DRwWCMk+OQciVZuXwgGysZcddk3JsYdCg1yZOU+xzjpF/0oyRUnUTW6oFEW/IadkrzAgBmOT+bPOZYyfG943r/Ghua46tBt8vHsX6ynq0NbbF9O3pGBsZiwZA2yA33IqtNYNVBnh9DuMxTx6OvcexI4fjmaf/IN767Zuyg3riiSfi/IULcfbMx/Gtb30jXv/NG3Hn9lR8/3vflc/7nTuT8aUvP639e+7cOakQvvrV5+Lnf/fLmLw1FX/6b/8oPvjd7+LShUvx3e99P/7u57+IS1cmo6UFxjvM5abYiU0x2rnHr776ei2nq+UGlQYN8+bev/aPb9TUN1prNDEbGuPxxx/VOrly9ZoAEayz0noMUA1LK9YGTficR2erFDOPWQc0KnjWrDUrNmyRxj34zRu/0XnEdZ45c1YzK2B/M1CbdazJC9tbAlg1xF1kIZM7WBM0F8h9AedlTSWijkktUrYQS9WYL7laI3t6l0DhWooGQ1HjFUI/a8kNfc4s4rbryoyr3ANAyzxjrWy2UkjWUfydNlKlSZGOjfVMZJ1RfCaasFsMCPc+RJVHHHNtxD2wqo37pliv3MLe4mLPFjtF5eUi99j2NvNTKcE194/cxOoL4qkb0E2Kv9SPIsC0dehzoZ5nT7P27y7cVR2sWlYDZanVuhWzraTVKazvp10V18FAe5Q/6RbAXuW9pqenrbDUnBdfJ/cir3cvcEiskRoEdj8K9Rbyqb6Ynp6q5UKZW2Yuy88QCzQPp8TUtPnJRoVBYCPSWSOYqOe8wsSHJLPoSyITUJuzrsgXrOJ1XsLfzIzLPHD3c1h1JvS6Wo3RsVHVuxcvXtDZduwoNitNMXnrlu4Vlk38Taxg/5AT7B8f1dypyxfOx8MPnIxTDx6Oc6ffj/ERlBajsu86cOhI9A4MqUnA5ye3QI3V2tKgepdGKNdEjN03MhzTt2+pUXzioUfirbfej9b23ljbDDUqLly9rtjAPdvUbE/HwfHR4WhtalDzY3tzLbo724UFbGxXY2r2bly+MREtnT2xtlmNxUVmTjqWqMlHM75RGXc0YXtZHDNYN6q1i0KovvEj4qKGlKPiLtayML/JAZW72NovcyruL3mhrHiVqmVuj+bX6wxiCYRCnhnrkYaGlHmlNkCBlk1LKcCLLRQ4Cs9RZNYGGvobsa7c2Lm+MAbsybOKLnUTzWHwGDW7yXNlDUcT1TNpiGNqYLa2aR6G9P8aSO975X23S6L6l5oE2dBwXWhSU/2e+ueA/rLKa79T/173AvTztbIhUv9e9ddc/7r57/rmRH0jZe81/EvvW/8+e5sk+b1siCZGcK/3qG/q5Pfz3itPK8SekcFhnfE0KlgDObcJ/GhgoD+amfEoe3OvV/4Y6zOWkOo9KcrLTCvyQggOiytL0YFNoYgru+o7WXwWkhurQrNWF+6aqFIIaibYmuzCbN+c4VXYZybiSU3mXCVzRfaXsRWfg1wnTWYraG17y3olHqaVHnvepG4rqe/cvq283ApocrtBEzYqY0/dWyd3rxXx2dc+uwO/B3fgPkDkpaWaDzsAfW42FbOzswK4EjiUT38rPrHLKhTV0AiGTLYJJHQxbImwhmkVVggHBgkAXcm0dalZuogNuRb3o7pYX5efNEkMSQ/vB9iEzzwAvRURC0owNFBKXunNZtSVIEMQq5D4NHggIok8QD7JAkUEm//OHZoEHrImaVmlIknm9evXFTROnjgR58+f14GtpkEnMwVgZgwLHDKbcFUMRvlVz82JlUHw4zUALygm8hCROmTbDC9YTBRtSHRzUDR+kFwH7w1rhqCET96HH32kewLIATOG58AhT8IsGwB8HFeQnHbofqPYyAF1Ur6sr8srW4mjWNMM7jODh0BJIlVvPyKQs6DiBnEMROfnsCLDjGc1mkpEZE2k3JIGlg4IAcI+sC399uBMArGCNgkMLOw6ibGY6rKSKbY25fdtRbDLOicPc2ccKboTGRUhxee9u6tXsyIo2FDEcE8BbWg0XblyVfZP6dUswLbC8EnbvGAt5MJrU2DP1iYAgtlCkrNLbsyQ1+J1XxgmvD9AmZo3pQigwMmBuHmAat5GKczqLbgy8c7mxW6jQkf/PaNJFiz+ZhZK/rfSxKKQKA/Q7Ypil/aJpKYM8t7YtmwxGy5uQJlRwx9ZlRWAgIahkr5kvFJAIJMstmEwbaXCqDUrdudhkFCo6SMZsRsVPF/WFENulezKy9GyboOO9gUmRrHuUUW1lMHtJPaKP81ueiYoBoCZMyo8C8PsM69/g0ySYpahn1IjqCDCEsYMYD5jqrfMgHNRlYlNJuNuuLoJxx7J62Sv5n6z5YGZn9lMyGIu1Sjeq2aVEU/TCovrMMuyvH+xT+DnVDxrTyLB9vBOniHFgKyiytDF/BmYrZpTU9h13AcDzJaasnY0q6D4ybpB53VIQS9bBg0M87UAZhSzr1JE8p4GmTVroFyzbYFQhrg5kclyFq8GLPx7GnYnEGGh2NPt2lTpXhS7u1qzrCh4soDG+ok4L7sn+VMnW/OTe8nFhb+WTEUKde1nGMN1TavcM/WNilTmZeOde8W5RZOas0eAvOY+uTDkvDIz3kOAadEpHrLWsR3cP24AUYNSbZkFMERSLuC9gYGgJOtI5D1orplGBYPXS+wSS64wON0QczM6bToApVOBwGvkmc/zlIqtqSow33G/xPBP+EAbqGTvAMYjzU+mue5RqijE4s8mnxvYflE36vI12Av4rfMZ+dzZ0Ks1arW6qmJWHb/viAtWFFWS8FQFjpMncO+5B9wvexyv6LlDZEjGJvsPRj4NgE7u1/aWmIYwFdsatmOwuz1GB3tieXFeHvOnz1+KuyvbsbrTFJV27N/MENUAeg1whuXfrmuAjUle5OId/+UuWZhNTNzQXoTkQUHPHAEGnh89dkR7HEKCbM84X2nuYOO2shIjzOXq75MSlVwHP3++riHRTU1iQVN0sx8gcrBuxcKF0NDVKUIGr+tGK7M/VrXGaHhgTSawqiFibdPX7BjbEGsrZuCzr8fH92l9sEM2sWSR6sWzeFaWFnXPiTfcT3yq2Uq8LveDvEj2MWXIoecXpN1anlmAfI4jAO38jIDxxopyFll34YG9tqqYilqEi2H9Q2ihqUr+h4JLoJkaEC1x+PBh7Tf2hYYLr29ofkvuU84X7ls2IT2DyTN2NEARMKPFICjL7Nlnn4l/MGshNQAAIABJREFUePVVrS1ZQlWalZdxbemLnSovnj3PmtwEMJ5/G4QjT0WhaDsKOaU1EjvJZezH7kZEJSYmmM9hJTFtMBj4fb2dVlTMzwu4vHVnWjEY9ZlY3yurAqsBs1H6HNi/Tw19njs5Gs0JwGteI/OQGVQBOwA52BsUUpJys1Zdh4hJ2AxAeFlejp7uHj1DNy18FvPsc34Fqg3qA2Ibignu4fT0nJTEba0MVadBgm0K+3RNQBT3a3VtOaKpGqvrqwK2nvrcF6JxpxK/+sWrssqigcLtMyFlqzxb8kyvRYIOViDkl0MDfXHk0IE4efxYvPHGbxXDv/Hii/Ef/9N/Fkj/wP0n46c//XkcOLAvTp48KSAXhvRXnn9en+cvf/CTeP4rT8eRQ+Px3/7iB3Hq0Qfj8OFDMXlzMvYfPBi//MU/xLXrd0S/LVi18thHH3lA9+S99z7QGuLf7Cv2MNfAmiSVogFObGCvsOfY76z9rBkM4DjXJodUQ3sbBVyrrCGoAZhh0hA0EQysUw98+ekvxa9+9auYm5vX7xgMBuDbipdf/pasbt5//3Q8+MCJ2Dc+HhcvXIgr127EYH+vwFGOafYD+yIBN82iKMA4IH7OHMp5O9WGotoUKF8IKiUHy7OR5yvbJeUbVpJYzWXFA7HMVlONUr25KcregzWNgqKwumsWZs69da2FOOW8y6ow/l2v5khlqBsNnhsntWxNGVzS63yYtWy6KEsLCcUDW7F0c2NCjNayZ4hXzFwk9qD85Wd1HrWjmrLPuZRtTY1qUhD3rQzZVnx6/fXXBdBmXiMiXZmzwV7HnxyVf+Z7SRxQg1cWddSw+2Qdl42KetKErUd21X71KtG9wOTQ0LBcDzSjAGsV/P87O6UkTEJNEm2yHjQDmea8m88mQJb7Wux0NBS9VDNaD4D4a1YBsA9E9qojk2Q+Qi3LaxFzqAXydW2VZAveejCY55z2dxA1BgeHdP1XLl/W9d1/4oTieDoecEajQuJcZnYk5+foyFAMDw7G1UsX44lTD8cDx/fFlfNnY6ivN/p7u+PSpUvR3TsY7V3d8c67Z+OLX/p89A8NxfzcbHz4wbuajzQ1PaOV1NXdGQN9fbE4N6P1eeLkg/Ha629HV89grO80xOT0bEzcvuP8e9v4CXt3k1g22B/VzY3Yv2842lua4+YNmpjN0dnTF/NLK3H24pVohCFexRYGCznnOpvbVu3CGid3IJaT54hdXur8fAZpPZxnZw77pQ5Rvl4wIPCEbMbzEHKuA3UxbHM/Ots+ra9DeCpWu2WANjGQHEUDsoVdOMckv0DlzXyLVAwZAHZODimRNdDSxBlpmx7t9yqzCpn9lRa14AJedFJ5tzZHD4z7dhrtqOw3dDZBNlMTBovmou7KWK6x33WNir2A/l5gPmvlbFY4ZzbxYu8eq28U5M7Y+3c9eF//Xvf6+r2aIvXXca/3uNf373XtWet82nXm1+/VqMjryvjvZuSuiqS+2aL8puAKWZvztZyDSF6Lson5san+Zn9kvkgzkXOWNatRQNStm67r8w+5SQ7l5ppYByKgsbYLyZY1xNqzitBNWjBQzZFcRiVG3eYmghRDZfC6FaWs25zn4dchSXXN7qZqqtA9s8x2UbZz8pp/4IEHVDNi7weumPefnA63gGxygGMlMQWbebAtyEXDI4Oqjz5rVPxLK/az7//e3QEUFWwEAjbArVQQGojnA+3O7TsKApLrFr/b9Ijn0CIpI/wQBGQFhES4gDRY7cC0a2hqiNu3p6Ors92+wcVqimKJpIQiCunf/Q/cr+SVoh4gBq9jmPJ46MLOgzFJog5ASRDhjSk+YR2R8FOk2OJhLbB+Igg88MD9sh96/4PfaaMfP35cRQLsNz4HwYbXgp0Jc/D0hx8q4X/owQfj9OnTBUzxgEp8qLleBnGd/uC07guAAcU4A/YAaElaW9s95JWijoBEMiQPzHnshkiaBuVhC7CSDHKC2n3Hj8X01HRMTt6KEyeO69oUrJsonJsl3yVgacaHgAcXlWRpBGVACyRs/EmWGcW8BqsWBj0AO38yaPK6u555tiRJoNrASRmSBCgJy6nMJ8hDJxk/PAw9k9jROvEQoY1gSDmNJewgbly/HgcPHlKxhDyTe7QGc6POB12FSxmiLWm2bGksu0vAj8Ojp6dLSau71AatNLxN/sDzMTgwHFPT09Hb3SNZPsAMn+falasxNjoqGwWaV6hYAC8AsmAOUjx2dFliyGuRrCdTnXsuML3YK9SaOkVpQNJGQV/rKRTbLB2IKgLxksWews0CvW4rwI2Hv+XBZwVFqiQMin1agrNXabGbC5hlXksN6v9NIlUSsTwM9Ty1nwD/aCgVRon8kxkobbmj5j+UzyUWIQ2d0pQRy6B4gIpF74ytMAdSum+2vZhg8tY1syWTO74uoE/gd5FGFhs1S3MBerH0crOUuMV/w3wwOGkAw/6mHuxrFpEZ5kqAygD1XLP2DaYxYlaN9p0SeTcYeD6y6SrqE4HO6VGclgMwQCnQxJKAVWs2N4Cqge5d9lo+W77P5+W99O8mLMss2RcoU+x5HAesVOLzeLhl7k0X3IA1vC7/zplCTgB9PTmzwmoN2zOJhZRKl9I8cZHMnJjdRNuNAH7WDBBAR16D4oHiDvCC/WhLmlYxvmkuEJ+ysck5kden+FRUEzW2fGHZZaOC6yAm87mx0GLf4f+dayUTTViKtmDzjKVc76zXgX4Pkcyiw43UXSs1/Xxt7oItG1jDrOfBQTcqmD9gYKDMAaqzJMhkPBnfvE+qbzSbR7OKbEuV7EXWIWCrwNqyxzaIA+Uc5SykwBUrsTTxtC7W12NpxXaFqB0AaNWo6OzUPW5raVMST/xC4SXLKnmgsh92tObX11Y0UwHgkMaGij0UhKU5lcxMeUNXHPvqm9Tak7Ks87yJBLP4N0sCH2n+ZDzgc2qOQEn0URUKIJVMn3lANMzdxLk7N1eT9LMuBZgXO0CtY83WaLAKoigm2WsoZ/isfE1WQazH0uQjFlR3ALmxenIzGpY+IIRs4ra2NPdKVmEMcd1Yidhci/HB3hju74qmhmosrazGRxcux/TCeixsRPQNjUZnN4qOhbh585aIAawRCAxHDh+RtQQgogH1ZVmIkVPdugV4xKyRFu0NPgfrg8HTAFC2JbLlEs3ubHbCFqP4ACDiWfi8bhMgBHtcKsutbV2H87MmsdvdmIfIYVsWYimFHsxUNQ+38VK3XzQgNXZOIlMIFHWs4f0AqqT0zMGZzC6jYCtzl7gPiqdNjXHq1CmtS85721ZyxnoWGAC8rcQcV7xmyKvSDs47lzyPsx4gTwNxAViQvnd1x5zYbGZRYvNpdRKzJ1A9gfgD+mET4zhOzOC9yQ+JTcQgkRHKvCieRT0gy/tr1gVACw0V9oHUnMjrm2WRgyUPZ7x+Twq2VtmbyvaiWI+Rd7pwRZnVK0k++0AxoIpdRpssg2gkcDa1tQHEbmjw9c0b1/Vs942N1ZrIANOZJ3K+0qji2ZJz3p6aVnOB39E5AhilofG+T8xJocEgti9g0NZWdGiweav2XKWFobe2r8ECyhZ5bhSjDrYNl20QucdcB7EpiSSy59NAaw+4pDHIfcbWjQHnO0EBPRxLC4CW2J716FmynolHnV1tAvY6xBSsxuzcdJw8eV888sijMTYyHlcuXo+Pz11Qrv32u++IdIKVycb6tmZV2D7MzYvuLqxRsPxoiNHhobh+7Wp88anPaZ399Gevxv/6v/zPcebMGRGQHnv8cV3zu+99oJ9/4YWvxV/91Ss6s773ve/GL375K+3X5577cly9ejnOnT0jK7HnnnsuLl68HO+//0Gsrm5EQ1NzjI7tV367suLZOAAaWOcQi/Fmh5nZ29st+zf2Beof29URp5djemba9rvrG/Hwww9rNh6NDtkhiRlqsA7w+3NPPK7rv3FzSk0ueAI7O9i2WHX0vT/6Tvz4xz8ue6JJzV88/CF0vPjii6qJ3vztb2NhaSW+/MWn9IzPnj1bwDvHzhwCLTVdUd8aPLY/fOZgUjnJitD2cWm35GGmjboXxHHOx1Tos8ewlzIj3jkg60sq7WI/zOfWf2OrtLGuaybGq54qcwkBovi+FJ/FLkZNECk2CzO/5NSKNaVBQm6keQdFzZ95Jx0wq3+dm0pF2NioM1aKwPI51ExpaNCe955wbcZnpabIJgwXQTyXLRR/b21Iqc1aQN3Eel2aXxJZzs0fk0bYG5zXnPfce1SU7C/iNg1CakDmytRY62oC+xmwWADkmW+VRA7OB2KDrZ9MzMn7sbemqAdkIQRyPiRZgWfovW+LuawfrRg1QJfK4FSXEmu5P/5T7CCLoiLVFOQsNZJRWhaLAOdBzYqjqvP8LKyoyNekebsdG6zJ8i75F3GLnJ2zcmtjXaotYsfly1dkp0QdyvUxQ4n4CCmQXJEZB4CFjbEjC07O3isXz8XnTz0cxw6MxuTElRjp79X8F+a89A+NRndvf5z+6KyeFU3PA/vHo6u/JxZnZuONN970MPK2tjhy6KBiHvY0hw8fj7feOR0t7d2xxlwJlI6oaYsCl3VI/FxZXIz5ubk4evhAdLW1KO84cd+RuHblWoDH0+C4cWsutkm91OhhpkWbznD+iCzY4HkfKPyop6lDmV3lAfbMrHDzwXbfrFc370XWU22KDaPnFDFomL1LvGHN7ip3bC3Z290pW0Ia8TTtNB9HA+HLkylqbOLOQF9/bG2uKd9hT62ucd46zhjkZ3g2zVqXzMyv6GDuiAZuM6dyU7kOc0RZ/1wvzYkq+7usMzUid6rR2c76Jf/kullbVraurWPNuO7fU14qzXmtVnQN5Vyofr/sBeezFsifzT1W36jgteqbDXuWrP4za4i9effe363fq/Wvc6/f+7Tv52e4VxzY2yC517Vm7Nx7L7K+zTjAurGqd9c+N3PA/Fx535JkxmtYydWsHBdgfmHubi1OptNGqmZoLpkM56Y58YC6RkrRUmvxN2szm1+cwarr2AOaz4X6u0NNU3I51hM5gvZRUcOrNpKKEhWh1Vql1211l+zNaUi36bzW59gysTiffaqU8r7zOdlH2FJCjCM3YjbeffcdUU1LHOK8uzExoesnhzh27JhmaB05ckTvQ55NvYYV6GeNik9brZ99/ff2Dhxtt9SIwwEQnG43SgEVaJWKNgAJQtoBAU5x+LGxSBw5QWDfolTgvymgCAAcsiRILkbtdUyiIHmwGMoUjnj/eygxgQgAhSLLHpdOdtmUJPAkAVwjCROHJ7YasDw4ZPhD8YKclyKS92ihuGxqiqPHkHjaax5Qi6SOIn6WIYh1MwpIVLgWNjuNDa6NREbXDfOV4X5KmrbFrPr47Dl57aKCMLt7iVNGHdiPL5w3ACZQEVZVm4o12DK2N6IzuykWlySWW1vR3d2lRgifm2CXcm8N0VldUZGpz769JWUA7wP4yYFLUQ+LhkSS+0dwhq1LoknDArAigySHfw4HxpIqrXUI2LYEMSMxDyEK/70SYQJxsiLN+HKx4OTVsyZgWGiAF6Dcpgf98n9ba8GeMYiATySAVTK2dKDB3hAQbBawWTZORGiO2XLDa4puNYcZgE4ypnVQBuvHoA3PtLevT023oYEBfU6KhRy2TNHAH+xCVHR0cA/N6tUsDNnKGLwhqU3GfioN0i5Jr7GyouvjZylKrBIw2J02BRxUFBWSxBYwUeBw6bT7WaVP5j/fqPBB7/BT36RQ0lPXnHAjonjA7pktkckC18RaoXjwH0vxBZCV+SUqTClYKXiyoMsET3ZdeySv5cKKO5YL06LMcEJqT3HWE8wJvqZmiaT03m/cr2RtpaKjxqgvjUYx/n21koIDOCV7DtUQMcTgfsl6i8WVwX9bttB4qSpxcfOAe0YMTJBan03AvwHZGkCexW3aFhW4nH1gwMjKkyzo1CIoDR01R8oguEzmZN9UCg2DYVboaHBYYQRqjVOgSmIPK6TIUUuzJT3Fa9deZ7ujQWLl57LgFKBe96xkv8YgvwQZBFyWz95AAWPf+Lm7c4qX3AvtH2y8FOe2bYlWmm6AV2aYlHkJtaHMxe5BDQC0BUXxE3ie98X6JizoRd1H3YMCMDj5dLyxSqMoNIoShHVCo4O4KOBB6hkKXt/DTFa5jzmLJfcc1w44y88BQmfxkMk1v5NAJH8Td/M+OrkGWMWzHjA1Wye+dzDH+L4GtMHMqTSr4FRcb2tXwsw5QHwj1lGwci6iBuR3Zamk87TEljLwF+snzpv+/kG9Lkwb9hrgj5szDD7cloIO6XyqctgxAqE0RJfGIcUy9j/YDxnIzs+Q+yHXcu4DhworG2gopIqRz5YxkX+zNvhd8gf2BHEXyw2xXQvNMpuhri+t0XGzJ7Q3Bwd79TWKbg2OL40jWf6VBp/irOJHNdbWYeHjteyBnbyRbVEqAqIPHzoo4ICGR2ulISrVjehpb46eNhqTGzEzczeu3Z6y9VNTS3T0D0Zra4dsse7cuW2bRpiY/f0BC/XmzZvaB5pjVK3G8PCIFHbkRlrHmiFjsAA2IQAnIAZNdfIw/OR5BpxbnKGca22A5hqqTePUhBHyJ+4Jqgyxx7Dj2d6W8jMH0CfjVXulAPxS7ey42SRAjwbWFo2pigFq3XcUOsQc2/FRdElRK8uWim3FGlgr+M+vie3PL/JMsNRg7ZGX8TqdXd0+LzbW5J3u/ARFpc987XlZFHqfpLKL9ULROL+4qN9h3SDvJ18iHooMwf0oTUAADggxahYUxeKDDz6k4cHch+vXb8SHp00u0RosayTzGMdzlF9uVPOenPm5/mkEM4yYRgXPMskFYn6rIN1RTokSQDODOCOqoeeh69+iIQgY1BZ35xYEvuAIYHYrqoLmePLzj8flSxddTO+gZBmP/ePjGv6cDX0aKDx41jhgJtdFEpTsQN7TMwDcdCDHoZhH9ctnbutoj9t3IMiwtgYU32zBQZ7nAazEaudERVUn72Y/A8AeWRCUYd7kpzTXuG/yCxdIZcu6lbUVNYkAdTs7ugPlBvTepUUrLdbX+bs9tsmtd3ZiqL9XYNWBA6PxtW+8GEh35uYW48zZ83H/Aw/Ff/vBX2owpXOnaqyvb5YBqM7LyFG4T7ByR0eHIrY3Y2l+Pl5++aV44423dc0QlXh+//DqrzUcnef/k5/+ffzRd74ZDY2VeOWVv41vvfT1aG9vjY8/PqcG4zde+rru34/++qfx1a99KQb6B2NqZjbaGKbd0i42PI077d9O1tf/y957ftt5nmd+9+m94VT0ShQSJNibaJKSKMm0NZZlT7I8M0k+Zc1/laxMPsXOrIwUjT2SKZtFEklRolhEovcD4ACn916yftf13HtvQOA48y3K4vGSCRzs8r7P+5S7XGVT821tFUlUo38ptsKYeOnlF2NxYT4+/t2nMlVnP8/YlzPqxZdeUOHt08+/cPNXOutIaoIQb41X/+RlsawBfrW3t4gp0dYGo4T11x2vvPJK/PKXv9TccyOhUUwW5vIjjzwiRP69u/fUUF1d34ynn3xCwKmz585qvxKzQUa6BtcQq1hiCSlgm2qnfAbzhOt3DOPYiLWsxl5BKwO8SDYIc1LNLPLNOkvQ8Syy4SCGg9iszjlc2HJwa0BWAfCUwqEipyLB5OZCVVw+z2PWMnsd85PfCale4rdsenK/Lc2c4fa043MEwCuSsMpTZRzsa+J5EkNlDpLoW85uNVdSXqaYsFracDPqm4y6VRzIc5e8DcbjZlKRZ4uNUPJVBolzgAuRVFRHh3LGBNCkR55AMOU+9+zZK+kng8YspcqapXlhZpiLhbUF0ywslqDfBbsiX+lnYiar2ZAGw5gN7T/nZ2ZOlw1wF+2yyOtn6QaQ437nAUb/s5+auaNgvGrUXppP2vdyj1bc59hSzWzG9IFWhcGT7YqRMb0+fPiQPhMzbT5r3959ymFo4BB7UfBTo2KwP0Zvjuqz9+0ZkXzs7RtX4o3XX46O5oa4d/tm7BkajO7OThlod3T3RGfvrjiLXnxzSxw6dDBuj96Kx0+fUvw6Mzerz0OqcmhwVyzNWxbr9Okz8Zvf/T7WNuuisbU9pgFfEt82WS6YGgpnM/OinSZkXcSBvbtjcx1fyAaBDnp39ce5i1diemExliXVSIxFfcQybNRHxHwrTSJ55dBAI3/e3NL5yr7AXCbmkCqCfL3sM8Y6WJHvGzFTs/ZWckMba5NTYRJs4JjX51YM9tN8wFduIdpam2JpEdAiz95zXzLP1AuYT3gmtbcpF886Csh1rbXSnVBuWOTYFN9JgqdFjTuujzPQHmw+D/km71vkssQH2j71Q0MaRQXmhWLEndCZzd5tbyZyQfud1iTTlfj3wYJ+rpdcT7X5Qe2aqn3fv9RIcIPmfhWL/Pza73uwOVC7djNmqW1E1P45r+2rmhHZZPF6q8pY1TZH8jrznms/K5sNWTeSSkENIC7zp4c1W3hvbS5Fs4t9b2R4dyzg9ypp6aIEUJrouhadXa7viU1XWEDJ5pefUon7sumgeVO8HdM8mz0oQRfyZZRcu33k5GlJfQAPGWJhGHPkb4U9YcN2N8GdI+HHhmQZuXp5QikP6Idkf8QtmN8rYlvyX2Lq23fG4tjRI/LQYd6TE9KEYGIDdKJeip+tVUAaxFJlnanM87X0U+1S+frP/38YgaPtnaJom4ZqLcjFRZthSYZFptRGs7P4aFSQNPN3DhhWRgdGbRQD8R1oJXBfFBIm9Q+hvWZx1xtRveQQUvqJYJbDj6SdoFg6mNtb2qBAxY5PjMsIubevJ/bu3Rvj45OSLeBgxZSajYODCUaF2CEN9dHfu0uFcWm5htEZs3Ozph3W1Uv+JynOHNj9fbskrUSixUHL+2A8mI2AD8G2CgdcExrAbCYEmhS0uD5YEFCpMcQmsWwSsqvBrILBAbEwkCHB3BDpp+7u3rh8+bLRSdJWZbPp0mZrhktDDA8Nx/kL5/UZBA/8ezJXhNxtc8eWsQVxxPUl0k1JvA55I2pdgHCQ7EDTz1SBcdnoXQgtps5Fdse6pn7eeXBlwTUDUxeA/bkcLDpYMU3s7RUaurOzW0U76HtK5tWddgEcU1jpYpfCJ+8VCr2gmN05Tx1WEIk+PAn0fU0UKHcUyMtMewsZkE4ZN3KILK0si8WjA2B1Nfbu2Ru3bt6Uh0gasVIMFXtDJn1pWOxDiTkO4geEOUUkIcNqfDJyfKCrZ2dcjZ6KLr3pzSmhkyiDDASrxb5sIlRRB1m8SUZFtXmRO08WQV3srfy2/JGgNJsTtQFFbeCUAYaKMuWZUOhS06RoLz6YBFS/x80PzRlHU0VuyolQmiJXi+D+PeveBtn2VMiEy0mQ5xE/RlkUNkl+R35PSVb0vYnUKMVuzYlScMogLxFrphM70MkErBpFJGXXyVUtkyUNQ/Pz8r2692ICbONomzxm4ux7sDRLFnozuVOwXAJy+VoUU2wV+YuXhFGCSRV1A5HxI3Fw0GYzbRJrvoN5QOHTxvJV/5Ccd1wryQfz301YS5JUGBel6C9/lVUK2qbRuphCIcBJhMannkSzKv8D2tL35AIzetdaxzSBhHBOBHW1QJnPQvOzJNDJHCF5oeCJ1AvrjnmZyJsMxhknPt8NJQdqlp+ol146iT2fbZ1w/3s+QxX3ClOiTKsKwwKEOv+ugn95Thng1z57PttGxf7OTOLZqzk78rpyzcgIEP+kwsgxetmlXopSSDKBoGG/UlMfE14KtPIdsvQXXjLS88V3pYbNxP1RGOc7KIqRcFFMUQOidDMZZUkWSWqBxpz1hXUOicXjM4KglzMu7zUbM5mguHlQTapAu0mGr9Vof/YP7kWIRzVcaEyvFnN19n3rmXtftAxIZS8piO5sZObYNYLY6+nSd9BYEKNTNO61aKUZQTOmFCxoRphN5OfCHIc1h0Y8zfcvvvi9kHwkAzD4GMfGuu2o31yJ9qa66O9uj/WVpZhbWIyrt8bizsRybDQ2RXf/sNYaBTaAHaCZWH+cP7kHa/0WlClFbJ4HzXLOfoE8iJPa29XUht3H/Ll77151vZazj7GHqUGjYnJ6WvOBcaVhdejgQRWxQMzLV2kJtky7YhgaJ8QxvJbxoRDNs861zHgieaW/A87YoDFcTc7zmeeJQnE9WTRcsxpIsBVWV4VwpAgnTfa6EGClUmSQL5Abw/wfcV3GMma3uQGlM76cBzl26XNAg47YkrMZ8Av7MJ/BM2MeiJKvvZNmraUFUwbgpZdeFpuF+BIkLfJa8tMqTc1ahl41eTaAwM07719CTTc3x0svvhA/++nPyvrg+tl3bOxL4Z+4OWn8zEUltxFiElu+htiC/QlGXHMsL8Ke2h3LK4uxsrKghLijjQbaZvR02Zwb3WJipll5dVhSphKLI8WysKjCphpgDY2aE8SnoILnF5bi0MH9eg3x89DQLt3L5PSs5ityTYyppHNA9RWDcpCCxJEtMCoAogCuaYC1AYNuVfuqzwAjCIlJ2aOJ6bPJxX5Nc4brYSyGRnbHzPS85KWmJyelsx47FHvX48TB/bE2PRfHDu+P3buH48KF89FCY2QrYmO7IUbHxqVlvu/gfj17/OZY7zB3iDgwTuVZ4mO3tDCvc+Twof3x/NNn4vNPP42e3s44cfykzCfHJ6bjjW9/M95++12Ny1/+4M/jw1//JlZXluLFF1+MycmpuHz5kgoBpx9/LH78o59ES2tbvPnm6/HLX34YC/Mz8e033oj3P/go7tyZiu26nVhZdeOLa3vqySe0XX388Wcq9jJOmq9NxIdb8d3vflsM3g8//EjbhZDwO/ZtopHyxBOPa05fuHBJHm48c2J1Gk7sE2JwT08ZBFakJiss58BYu1fNiCrz0NrysHAeOXYsfvvb32rdkKPRTGEBPvbYo2Lw6Awsi17F+MJo4pcuBiVLwN5+eE+ooV58d6Rbn0W/EsdljmXfMMslEX84/veOqXMEICRzAAAgAElEQVRI355uumVfKDKb3L/9Sh1XZBNEHhYg+ZFqgyUoAJS9ZeRhUaSFeA6OM4z6d1DpGETIcfnaWQ5ETHh884K5bZkP4jmdYwWFLZDBlveRPC/lS6Qir+NWwXlKbCyJ0DoDALSfwAhmzqoR7MY55zFrEuYV65lnRPH0tx9/rHFjjbEH8+z5sXyJY8qMlWkOkoOmpJ9iDKHh23X2PFhIrSQMNVI1mceRJ/M+nm9qsDN2aSBeyd8Uc1bBDIx1NknsT5lscMf9yvkrTQqzTdNX0IwdM5kTfaWiaTaOS0HQFm7O/VTEVqMiGemO71NWTHOlvk4MJ54tzXLeScOSgh+sei6HcRsbuxN7kM66e1dAkP379gh4eev6pfjWay9Gd1tzzE2OR09np0ytb966E+0dvdHW1R2ffP577ZcoOHz6yafR190Zx48/EoND/t7Z2akYHxuL5aUFNWpf/sYr8bvPvoyG5o7Y2GmIm7fvxOTMnOY5+y9yWPLiwHtraDBieyNGBvqjA7YcsdnqagwOjsS5S1diDN8SirYNgLVgQzcoRiAekyJDM80PwBj4uDQqdqF2ksx5eXxhmI5nGmexWMWbOvPkk1IAW4w1Y5fFZP23sJJ5TqwPxoXYIhuDxAsAX8WSogGZzIQS77chiVb0/6k98f32v4HpsGrBzwTu8Tc1WnaipRGfF7N1iY/ZI8jjydWpnxh0ty32DP5jxfZP529He4s9QxsbY2Z2XqwNWGfK5cumVMvQebC5kEX32vXz3/rnh+XguY4r+VUBFjrFLT6HZfxq4++HfXdtYyI/Nz8nX5+vefC/GbvyOuZuvv/Bz8yGROZTtf+euVLt3vDguOUeUjsW+Vm+xsIgbm52k5TcvTTSJGFXJLeJX1KCmPXCj0C3pfGejTfLj5tVzwRxXGPwFPtE1s6I7/O8SiWACqCvgEmZXzpr8GDCT6bIWBscVGXRCzjBvi+mkKWS5XckWWzXtThfkLI/eeJEyTcB9mzobGPfhmUPcER+cb14gDVVfMzI0YnvVf9k3QHY+bpR8d+6HL9+/f/XR+A4MgbI3BS9diUdaC6TgO6EzAs58Aj8oO6TEEl7cWLcOm8Kumx0xqIxSwKaP6bJVTmZSqJckMKwAEhuQIImBR8ne7r0t2/fERISlAPBG4EXFE2aB6CC0F/FB4LFvkxy19GmABtDHAI9BZnLGNssqTFBAjV2d0zdx4OHDun6btwc1fVSUGJDQ36BgxkEFe8/dvSoNCils4mM0cZWjIwMyhgbOuiVy1fEbKhogq5vqOvJwY4EFKgN4Qy3t1WwIlDiHhgfAgKkN0ictXkpUN+R3AiIHFAeFOlIstmwGDuZ7KybxUJxgnFJVFvKcdCsSFktIVeEADeyLyVjSKz5DDWkFpZF6VSxb8vXzDOV3EKRaoEvk5s2H8Q84FlL3oBAGF8AkLuYRhcd0izIktAisyWUdQnkRWeGdVA0d5vb2szKEYPHBbOUDyIIURcbo+1igElS4iIrGrRIHVAgaxadnCAszX9JCoXQkWySze9o5KChDfKJggrPGcS1TE2LQbnQemJEOGim6KPiOTIOvegMu3DLM7PhZGOsF3S3KN7Fn8BMBBvvpTGgkPJKAI2088HuIqpRRu7UP7wh8SC5udqYuD/h8N+qoBCjl1LSyMGKWQOmj7ux5AO2aDdS1KWJlDJhNUi12u/y2FabFApohMbxtVJAqpWY0nXBgBESz5r8ZpEYMSeGlhIOTNscOKbJaiZQWXTO71CQk0Oj66kW84W0L1IWqSesgmVplKQhHKgusTb0WvsnqNCSzYVSVCYgUUGfdVC8A4RSQ8u8ppmrpgaBe2HqVOY1iVqNDJCK2IV9k+OgQnQpZGfzR0FNCcpsJGhZsGQ8yKB2eUXa4yk5xbB4jdnjIwtxyY6j2Sw5rIqUkcGLSZulAOm5bHaE566Lyl7nNkxW46AGCSlPhWKKSQPRBW4H2dn8Yu7n77IhVIHUl7nDZ9DQhR1Gg1mNmMJuyuC3MgdKodtyY5Zp4nrZ02k2UyyWSTh7RkXGysidvI5kv+Ta27WrX0EtjJFk1eTcv69JVaTIKtdU0Ibs3xQLszjAWCc7MBsD3DsFORIstWlKc499RvIya+s2aU298tKEoUCKBIKKqbAYVFT1fbOv8V3zi4uWVSqmt7q/UhRyIdbrLiUYmMMqGEkSjKISvhhOlvk9+xZ7oIpjRYKMsWRvx8CNtU6xNpGWzB0aFdw/Z4CQSEVKRGbppfAkFDTnj4L3ep0vNCCqjdeariummEMD0d3Zrc/iuRDEs4+AklOxojQmZPC6AzOmW2joo0ePxfkLFyXxwD1MT1pqCYkakn/O3Ka6rVhfmIuh3o7YO9Ivz4qNje24PTkVN+4uxtJWRN/gcDS3tKkhjy8D6PG852QkUEAi+ffe4AIVTRrYqfyZAilzG2QzCEyKUphi2+fJmrkCAayuCvjQizn1nTsaJyVUG1tqSLDWYGIQsyHJQCOdeUfxGYCJ9KbVsOR99UJlS0IR0EN3VzG6rpf8ImPnprnlJjOpM6rYoBUX7Rs0xxhfCsXsBcvM1fXNOHRgrwoHJIugPbkGoZiLZOK98XuVIlbBYJs1Kdk2I9aSzcm9dXR0CZVPwZbvp5gun45Wy5yp6LJAgX9ZsVADxeBSbGRuy6y+JIXMK/YAilPsgTqfCjOY8WctmkVp1pbi1TL1+Duvefa55+KnP/3ZfUzD3EP4fiSUMv4VS6to7bMPInGkoh/J8iZFaXxhVgMfHSSDFpeQ4ojo39UXTz7xeLzzzi8L68CIVjFUV5ZjaGhY967mEGba9ya0RxAbz87Oq7h65PBB+bwtLa3Kg2F6alrPl/0QEAfm0BTALVm1qviFWGZhyd5hQkIW/zIVTBVrmbXDemM8KPTQ9AGAQnxN8kxzFEmzwcFh/Z5rZA0SQxGn4xu2ugwDhzhhO7q7YB8sx7/69jejbWMrlubwM9nRvL83ORXXR2/Hvdm1qG+uj6b29hjZs0eAHDwwRnbviQ8/otjfEI3NMI1hIa2qgSt9+cFdceqRI3Fw/9549+13Y9/+A3Hg4P74u7/7T/H6N1/T7//vn/xEfhXItQBcunDxavzZm9+J69evxQcffhxvfu9bMTM7Fb96/9P4qx9+R/vc+7/6IF76xjfiZz97O26NTUVra/G+kUn6Wjz11GkdkR//7vfR3tYidicbbVeHDZOff+FZFR/GxsaUb3CuwUghpyD2AzVJM4ozCyCS2KXlXE42lCRjW1vVhDcbgUboqmKQJx5/It5+5x01hBSvaK91Uebf/bt/G++++57ykWeffTbu3bsbZ89d0B4Ic4c9ntyFNUahVMhUzVkX4bOon9J+yjEkteSYwLElzAMzc4jdZPpe2K45/20ybS8LAQvEZGiuAAJgtshHr9FnD3Mr/R5g5dOIVOGq+NGwPyXTVvIvQok7FjdClTEyk1tI9SITm/GNSmIiBCaSuTBpOfOKrofkQYu0b1Xjv/iCFfmnbAxkQ4az0WyNFnlU8D9GSfLIbUjYGNnNXsfr+HtzKywZs07u3B6Ls+cvFMQtprG7FBcQs7gJakaGATVmtPCMBNrC96SoEzDWsP8qMVZFevN+499KY2V7W2ua++X7ahslSD99VSGV/ZYYJ5kzblhUwVRmT8OoKDKbkr4kz7J3j5u+lsGqMGn0YgOanANYqiVjFWLgjU0zKhL0ZZYefj49WmvINJF/U5Ng/+I6hgaHNM8593km+w8ciFu3RrV/wUgBmMbeSa575+a1+MbzT8VgX3vMIxfc2aW46OKlK9HZ0x9dfbvi3KXLei7Hjh+Lq1cux97hYe23axubsf/APjEjx27fiomx26pnPPPMC/HJ519GV+9AbNc3x8Wr12L01t3o7et2QV/sBcYlYqC/V5JK9RQ9G+riwD7qLxPR1t4dF69djfnllVgTm7VJBfeWJoyF2Q+azJyGebC+Gq3I4dIISC+zGkCF43ObrcsHgFHh7E8Gc/oQlsaY8y4a9JYc5AeWqQ2xDV5V062uXl6RAA6SLaVnXBpQGIbTjGC/amlpkHRZJsA0dIllswGYUjubNPvD8lN8F2uBGCHZmcRalmeEhV4ASgXgJVZHYW279kF8uiJWs2Krsl8moimL6A/+92F1vSzUaz9JYFBV5uC+t3xVo6K2eJ+5Q+6r1fldnetfVV/U+siaS/ECYhyTDf1gcyKvuTbPTlBY/pd/yziQ9yeAtfY9/L52f8i8KD9fIJaaxmbtWOXva8eGGA1ABQ3SjlYUWlB+WVONiLlpkJ7ZXTTjAEqrvlL8hwwS8L8n4Iz7sXqIz0byAWpybkb4THPjYks1Mc4SYm6uRWyx0k/n0SZrkbhTjXEZvAO+JFeGmdsWK8uL+jPXJGDm1lYBcJjRzHlKjnv69GnJtwPuUF212Wbwd27ftlF9YaaQ6wDYllKMPmtFeS6y78z3rxsVX7Uqvv79H+0IwKigkGBpDCSIuhQkpbEtkkZa5ARq6L4h29Bsajmv48Bm0ZP8ERASHKiLvgzNF6RjVS/RHhYgLkHhmZYObTo76rv37JYBJAUeAhCuxQ2TnWI+16EGBMhIDmKaBiTlLHSK19AhCURmZ2e0kXFdR48c1QIn0afjyOJn0SOZUEHq72zH8OCQAmcaGiSP6IES5HBPbR3tShpIDAhGDh86GBfOX1CHk42EQoHoYej472yLQppGn9r86iIeOfaIk2RQCqvWVpUOecrg1O0oOGTMLD3Sq+ItgQVBCQdvHmJuUpBcg1a0dwSak+g7Z0FQ0g1FszjNgSXrJDkX0/hV7KEwJEkMFw+NArP8kjZtJexVhJPRiEY52LjO8iWMpQpHqzSooH874QWZhqEYgRra9RRSGFeeHY0jAhaKG1UPik0VgXXgFbZJoqhIlPkhiaHQQl1FhdBtkHlGmXCI8SyQ+yBZHhwa0iFAIsD9UqCCBSMEO5v88rKTJEkbmULKC230ZZ3CbMKlIakYKKWozVgyn0gsScrVKElRzRKsEAwJUV6aG6wz08kpfBcfAZkyVtkE//UNxcF/UWypFuprGKvCsKZ3cEFmZICW11cJphLJXu+Dj3Wexr0qJJb7uO+aBDhVSfM+0nV9aRpks4r3VhHG1jJOtF8F2VoQnG58FjPsUtShANGM7IC8CEoSUwr39zUpNCAl4yw0SzNCjPxMzWGej+ZQk+/VZpZGXzto8rOXnIeCHb/fY2kUIAgtrofr5XWWznOSbpNwKNcO3pmfMmatCc64bsYgC+BCx5TGkTSQU8Yg0XlFU5n9LBH7iWbh9RTTr129Ie1ioyVpPFev100KN8VkOl8YSRR2Kk2U9GEoKSKme2nGaSo/H1iks2BKyKvCWs45P2hkNNanBBfrek33wrhZNiDUeDDq2OwL3uv3V6WfVFTd3hHKE8k/zgPGWZJVZRyFBheboFh4FwktPpNCN8UMDEwxN5YHQ2nMiPVQ9q7aJkrV8NvXg7cO+4EYhcyVZJHUmAPmted+qM/etokjchrs2xncsycZlW5Daa8LI/9gFyhxEOK0Pvr7+qRTynOk2AAClezeeyISZdZtNk6dXNSRM88V5h7IaM50xpEipHOlIjlRmhG8M6+NRp3nk31P3DDF96cq/aRGJ4WQGj8diqfah1Pyb2uz6PRzjy2OKba2XDQXcyX9bWh4WFM7ExcvPsuppXdHwnvz+rmukeEhNdlhQ3R1dFYarYyBi9yWCPMablRxFYRkF2aZK5bmSFYia5SiFZrSfPbYjavRUrcTewe74+knTsXa8kIsLa/GzbuTMTq+FMvbEb2Dw9HV3aNz7t69MSGylPi3tUn6iTN+YmJSEgN8F7+j8XRnbEzPBKbO5PSUixhrazoHKTLDqJBBM346ZT/hz8RDxEn8O/I7yN2QoPM+frIZkHuzzEw3N+Q/QMGDQqFigqJPLibHEgXvQc0vFSZ0ljnGE0JMKGNLq2kvKqwhxVnNzQKQEKcsgEidmpAMBkUKYj8KiWq0FiZHR1eCLRqFGuOec5917GMkGwwNMw4cXxC/UHyYnZ9zTMKe2QKLBkNyCjFuULEXg5hkrVLTUnOtFEdhFzFfiQ05r2G0ulhGUXlFkpMJNsiiAIUWyx81STYim5LsJ08/83S89dbPK8hus95sCMw14UeQgBzLAbiIsrm1rqI1Y6O4SiSTxujs6Io7Y3fUkFhaXowWDMmJNQFULC3qXmVQvrwsXW7ibQpp8hHRXlin5gDjpOvHC6n4l4llVmIZxZxra3ru8g0ohsBOuuv0+STjSI5wHooZKJ1/M+60p26s6+zIBN4Spm7o8PxoHhB3M7YUiATEqA8V94eGh2JifCr6enqF+O/r7o7lpbnYWMVUviOO7dsdG9MzUb9tmRNkG2mw3hy7F3en5+P2+HQcf+zRWN3YiIlxG86efPSx+OLLCzGK8S2I6rp6MR94DhTkers7YvLuvXj91ZflB/fhh7+Of//v/+f43e8+ibv3xiWzxfzBr+HAgQPx6qt/Ev/L//ofYt++ffHaa6/Ef/jf/vc4fuJkPPvMmfjgg19pL9y3f5+Q2ICZPvzo45hfRI61NaLe49DS1KC9xAbEBhfZVNkxj5s97P32JqOQz3OxlOm25HlgkLOH0MSEeQXYKgEwfM4zTz8ln42xu1PR1EhTEdSwAz2Kgz/84V/E3/7t32kfz38TaGF7K/7N3/xNfPbZ53Hu/PnY1dcnxDdn1OWr1+XHI8ZE8YAwu61CPrD3Vg3CN/EhOlr0e9ayi0esXa5VeQZM6TrLIzI/KYLaGxCJQDOlzCZkrwYF689T86F4ODEPASWx/xiIhcm0Udf8XU2JNRtPs2+JxaL31AAkCrjDeU0pVpZNMwtxFF1dYAKMZJAAZxChE3uIYvhGF9TFwG4EQGIZQ/1d0js0dX2OOvazT0Jdg+Udcw+A8aYcqkjdkseSD7EvOVZBQrI15uYXSuOB4ppzPqHYS4zowiGgFLx5XJTlh3wxfdF4Dc+5tjjJd2dRsTY29d6MZCGeK8tm3Bd5S/5tZma6EtM51/T6T/aKYyqz0lP+xMNcZVQYX5EG7MnYtZea5H1K3pvNB5rHYrLrrEABoOpvx3evab8pnJySm/LMVIx0YC42EXnarVu3BGqAyUjeOz0zresd3j0SC3Pz0d3TFbdujmp8jx4+oELljSsX4hsvPB0DvW2xMDMdA319UbdTF59+/vvo7huKgZE9cX30lubcoSOH4sK5szyQePLMGUm3UD8YGRqMfXtHYmVpISbGJ6K7uy++OHcpGls7Y32rLsbujcf10TF5vSF/V2GD1tXFrt4eST8hHbW1vhZrnLW9vTE4tDu+PH8+Lt+4E80dLdoD5R+F10O9G/MqsrK/bG9FpxDXVRNgmnc6n2Qs72eWsSnDpny4+IVkjM98dXxIE9TgNvY11jdnUSaDpGAYf+MxyhhSfKXuIakmGokl5oBpyGenfC3M3C787sTU3AokaDmfzMrFTwvfCse8rjtV5VRZezR9W4rUJvswdSjmgPzp2CfLPOEz2gDY4OEpCVE3TCz9lP6QZeY+4E/xsPXy4O8yHvuq/+b6e9i/1zY5cs3m6/PfMq96aG5+H7vI9/Lg59R+b22DxcvlfrknP2/Lhz/4vbV7SDZSHnx/7XfVXm9tUyZfk7+rjGed/W+pA/LsiGk2AakIOE3cYkaN/STMsKVBxvdUZYutQJDxSkomO58y+1lzEgBIqXWyjzJXib+c+8JOLqCx5P8VMKvio3XX9PhhP7E3kdnzdYWtDmBKPnXUigogCYAXspX8/dFHH1OuOzs3o/mfOSSy5QAZ2Ltg19Kcw8/i/LnzAo0T/4nlvbwoBZCvGxX/0ur7+t//6EbgcKtNsH1gbWrSi04P3RaNTIq1JYEWAoZgVGaFTpIUhDc0xsjISICYa6xv1AZCYAFCmqQaJgA/0vJubIqF+TkheNQAAZ0FQg4zR/SM60MFZlAUFBlI+JHfoNhNgQJEGYfaJflAIIfUrWC+jWYBSP0NmzZ2d3RVdD0JjEnyZKxIsai+Pm7dvqNCfqJvCczs2UCABZIUc+U5BY9svCsba0Isknzs6u2NlSUK3G7QsClBIe3u6ZGOMkwMAqV1zBJbWlSooOnCOHPtJHztHZ16XfpREJgMDPYrsVHwtbYeg0MDcfPGzdLgIPAAndiiayOIYNwI5oy0gnlg4zZRNEtRyWyNgpgvMjI2LwsjtlZJTo1A4fOE5EAPWoGhymAVqqf1RlP6xQgEMxqsHU0DgsOE3yUFGkNNDjCKLT4QLdOlA2drS1rbFOryEFE3XBIt7kDTtOAZcb9s+gQt8nzgdxvoYGOc3KiAiGfsAjnFHoI9S0+AwkN+iyS3q6NLyCTGimJOBvyMo5A9QusYKU4AZmSgizhiwkir07JA6bchPE+h71cYFTXIExfMHVxJZ1+0b5uVGZ3uYpBB1X5tBvd/uKFUmxSVV1X8LNRa8q+Fvi5JpE/9+/6Nf3IDwUV8v8SFYyeGWy4Qaez/0KxOqUcaRJULUUBUGBEKONJouyAxJPnV4AJ3FoP0OeV1zGPWnlgmpVjt6yvBdTGzzsRS9P2KaEAZPyGuipxAaTo44bbubWoa2/+kSJoxr1VcM/rYDRDLR6l4V5Bf1cacDSCZWxj4cs0E1JJjYryEeEWGZ7AUhcyIMGLDz5jxycJ2yqqkXnqlaFYYGBQsLJmSs8JyUw52tu2ls76tAiXTSCgStDMrpsJOCrkmJwAMahp/uQmZQWZ2ZZCboZGBxEoyqpKGbckn7sdorSzigwCj6ZPBrhJSsStAENvglYK9kluSoGJ+puJ0hUlipCVzUGt6bU3ycTSruL+8ztogtxKIp3cE+rttlv2bmpqu+BhoLkkT3ImRmh2S6TI6yIgVN6owQWbuTxdGRW2CwP3ms8uAmt8lYod7JZGkYe1CgmUTpfWvRLEU7GW05memz6TgsLEVQ4MDaqQjycieDOJd7CIx37akdc3nSeIq11zZV5HXW15Zs8F0aRYzf0kq8xr5QhlSFlkG/mzmV9m3aR5TxC+MIDc5NHON9KWYKN+Cqhk8gXqubc4OnimF8JTDswyhm1Net5bJ0H5XGqx5PpRqVVkrubl4U6TQDwJYgAX203WbQKtoVRrzkhtCcgck1hqvo9CKbFaD4hvWPYUifijyJUJ/c3Uhmra3Y1dHQ7z+ynMqCIC2uzE2HlduzcQayXFnr85uYgzimLa2Dq0/zhTYDxTDsyCMdA+JBAkTIAefL8xBm/HpzG1v03WCeicxktxG+TePo6UY8lkQL2XjXoUgPxYX72GIdndr3hC7qKlZmBBq1pX9HoRyykJyLtPAAUmYzXSvZzPTUjecNYJ5MwAO6OcUjHhOqytIO1jqk0YFcz+LVaLGw3KkkNXcIqZsmm8mEEJzVPdr6btsDNjTBK+eDT0zMVRAhGqeMu/NeGAe+CyDKm8DeDEZmhrj1Vdfi+HhEa3xzz77LC5ecMxY2X/K+lDBsBT2tcer2WiWUCbdNCqefOrJePvtt71/l8Yy64LnRJwHcjS9Xyw14/0ERkVTU31093QqJkRDnB6rTE/FsETeCkPeZsWvPFdiGsUExRgYPe80P5UfTZHvtAGo5YUyLuQ5Gv23LhkOGmRq3ra16hmnGS2x+OIyzSpMRde0b6QpKftWxRtK8YHjFOJP4qDcD1TILBJE/C4ZAN71KX5vicVBXDs/O6dzq62pMVob62JpcSGef/bRePr0ydjGAH78bmwhUyYW1krgrHLj7mTcvDsVB44c8p5d0Izd/f10VOL9Dz6OpdVNGR7DrICpvb21ESODA7G0sCj5tje+9Zo8ITA2HxoZkvTK739/Nt544/UYn5iKDz74dfzbf/Pfxa1bd2R++9d//Zc6Ny6iO9/UGM88+3RcvnI5vvj92fjen35b8iF3xyeio6s3GpijRRN9ZXFemvase0xt5f8iM+s1+evQuEfeAV8eZKh0rhOzU+Aosd+LL74Q01MzaiaoOcDZJBmlHRUxn3vmKTUbpmbmQ2hknTsUkiL27B6O5559Jt7/4APtNZZ3bRKinH3n6aeeFpPj8pWrQm4C4nn89GMxems0Rkdvu7DCmVLYzRlvWOLCYArmjpp47P2sQdipTTAf/G9iLpUzjrmbfhU+Pz2HaKDaa84sDUkuATQqmveMp/KYZB/Ln8c5QO5hNcGQ5hnzih9fZzZZzDxwkbyhXDtSG86P5FdR5G6Z01not5QjBuVtKrLyXQZaeEQsYZla6Y7p1PDFM0Wsza3Y2XQexbOnIK5mlNgq+JW40agCYPEuq8jraK9M/weevY2QAbGlrJKkRCufk0AEx3e7+ndVABKMNd6H/HDeZdycscuDxc/aYiaAMp5L5gNmgSDrZPBJxkAJNsn35vM0G8dFwGRymD2TnnvOh8yogwWTkrduiLEPV0FcPCvveYwpcUfKFGvv26gy8RSP8b96+wyx31FLgFHBeykEsmYk/TQ3H3fH72lfpNEKgr+3tydmJqdifX01Duzfq/z+5rVL8a0/eS662ptiYXo6hgcGlBf/7tPPS6Nid1y+dj3WtzbjxMnjcf7s2djV3S2Q3vjEhMYfZuee4UGxN4lXbo/di08/OxvdfQOxGQ0yz+XM7u7pc5zUiMzWmuY9oJRmMSI3Ys/IYGxvbKgxB394am5OhtpEAsTeSCkjPGZCRJG3xRdiayM629vdUCxI7Mw/BQIqhdXMUTSny1koGcCS26QUs9aZZERdnGWPp1GvNZ8sq21ULqiRgIrvkhSgzdMxD16PdVQc2trMmpDsreWh6CcAykApgTmXfm1iSPH+LTNEWadc1/QMZtxmWcAE51rIf4h5kANkTGiSSB6yyL+yXVB74L9LYgnaF1A1Djld3P/zYEOgtrhf21j4gzeWXzzYDPiqRsWDhfrav9d+dq7lr2pUZEOB97BuMq562Oc92DB48LNrmxF5H68A54oAACAASURBVLn+FX7W5LP5fXmtldys/OJhjYraz6i9RxQbaOyzhsUuQMZ9a1uNCMc/BlHIU68At5SXlpoR95EMEgOZqnUl4kmeP+sc3xQ34avy5r4mg7aoZxKzsfcx59KHlO+G5aq9q85sE/Y85hr7GvNX8wmpMiQcYb+VXJN4iO8HlMS101h+8smnxHLkumGH8HnMeeQoqT0CLuB6+A5qo0jVqS6gfZ64vNsska+ln75qGX79+z/WETjW2S1TSskbra9HT3dPSfibVHyTTmBBmLHJr28SvGyrEEN3T2Y3be3aBED3cRCTeLPwOGg5NIT+qrPRsBAmzRjMWAKGg48FiXQJQTPG23QO52ZnYs/evUI+wIZAqmn37hFJN1EMAHGkohsyIvJraBMaBeoXgQw0MRY7i1hNlHv3hM5Dg5IEAYSjDi1QL3TiOzoUQKBhySZ48MABvccJ/1Zs1u0IsbV7ZEj6cNev3agYa5OYwMSg87mrv19azJyAQlc3F8RlK0yFHRUsGLvWtva4eeNGoTiT0CItNaLCOPeHJASFtitXrhR0kpFZbFIEW/guCDFXdARl7iY0kVE6SctTM6G8jiSZf8e0B8QeAdG98QndE3OAIgjPGi1iNlUCOcksUUgoGzdBM4G3C7hGQbrw5gOLZ0Ahi2slEbp167bYFBMTUzE8NKR5wQ8bvpoSBJX4cqzYLF0HXSloJevDyCjLH0Bzc/GvHAxCQG3rO5hPNNZI0pG1YvyQ28LInGdP4nj08BEddhQ0YKBIwknJtiWpZIjeAZ3VBwDXy8HhAqOpfJadaKisDQ4RUMzcv5KuErx5TzCbwqhjEOXW/a/0ImqKdPp9Sbh0UJZXPUhoSDapUNE1n1RpUlQ+s/whRzbfqIJuQbPLR8AHdAa20n6nUaWD2IWgpMLet89Zcaby41aIixr8CPlVjViK5NL9uo6J+jKy0IwJBU6lgQHy1AVVq8+L3VOK2n9w74VRoWJgaVJlYMoYuhnmsdd3kAXi07JmpD6FuDSapXjA9yTaKIMWoXq01oziSs3JRLAKdVLmCUVKXqemUZFJYF2qEVQkCpKayvUoqOL3xVRaa7h4hajI3Ii0iZtIvN6JpIvvzU1GZfC5MrrWnDO1Pv9uqSg3NxlUmbHWMGbSk4TPZg3kOif59rQsyEmZiFkf2g1JN12gVSvg39gwu0syag6S06RSn1kQKLkvyZBP5nY1zx9Ww8CACjk207ZuLtebxcNcL0ZzurmhRiMFNRnudcbU5KQbXVy+shkXMTLQFpq77F05Vfl39g7mgph3NR4PmaRnwJiBeG2jgmIzTW8aFZLsW7OhdRY7ktnkZpfRbEpGhRJaib2794gxsLC06IZuKTgzL9I0jkIUNF8nFeB3vdL6Bwb1XDlHtD+L8mz2j9CYRa7PCEi/V99RfHj0lOWB0iT0pJe+i7sUSzhzeRPPNfc61gAFTMYJmReCb8ltIF1Q49sh2bVsyBY9bxeVXIjL5l02Kh5s2GpdqyBmXXKaV8lCQfpPTKZSzNI8KbGBWCyg6iWHRlHEa3BtdSU21lkDmFMuykS7Hk+p7ub49msvxvLifCwsLMW5qzfj9sRa1LU1x2Y0Rl//gM5PJBhpnNA8p7AD8otidZ6l3CtNDTUvS9GtUGB0FlGAF3sCBkFpXtuzxwW2RLRzj8wRGqEgprgHpMkYN1gNkoqQx5C1tkmoxicnLOFQoM8kSjBQ8Lqg+Qiim6YDTUAMeSvbtJ6X44d89sQDnJGc+SDM7C2yIWcVUNudHS5GEENJPrJIQaipKDN42IZ1igWcxBn5rxMHeTI1C+2po98zbqUYzquYi7oWeVBZnoXx03pBVmwDgA3xFRKRjhXY/9h/+VzmKc+Fgi+ofzP6LJ2nc6pGTk+FocL2NVOpGMS3tseZJx+Pd959r9LUqMzbAsQg3qXB4uSYZ2itY4YB9DUSpdwjEkGNDS0yPmU8b98ZlXkzY453A8+XWATWC2bXiuc2t8SmIC5hDxc7uakpFpaWzcTo6orJqUkzUdrbhRRGTuPo0SNx7964isApF4aXBmNOzJRsFuawdMSl1+0YBpAJz1ko+SY3rJkDnUifwJ5dW5VJLEkyf6ZJYIYKTe4VGWmDJGcYafyOj92NHc7Dzc3o7+2IjbXlePrMCbEW1lfmowXfu6nJmJ6YEgNjp6Ep5tc2Y/TuZLR1dFsGrbtbslMtXZ3SdP/ot59EXQNFpu1YXnFxlBt57NTxOHrwQHz+u0/i0KF9ceTo0fjwww81Jq++9kr85D//Q/R0d8Zrr70W//iPP1dz+MyTZ+LKlatx8+YNIRZ3j+yO//Tjv49TJw7HqVOn4u//4a3o62uPZ557Pj76zccxt7Acq+tG4IuRvLEZJ08c07O7dPla2ZtcIOGHgtmb3/tu3LlzK748e17mrvwLDJQMsfBBISanmcC/V5sFDWoQPnrypPIj1hVnHAU99h32uATTiOEFe1wSFJZrpQgLW+Pz33+ufRZ/ipmZ+RgZHohHjj9SjJqnBLRyfE2x2A08x04+7zNOzCIz85ymrWROt2k6UEQ1mlTG0hQWC/ClgrQXgttnmeM9x2Ri67E3lPO5WlTz+KlBWVgWBkA49hD7XwxVs3HZd+RdUXwqWKd5brE2KHIncENI4QKAyTxXLJkSw3LtrGvWIOcq98T+yDp0M8V7pQrraQBMMan8vlKmT4a4GMVuNmvPLlJQij+RU9sEnQ4IAEBdQ4zeuq39i/XDNQuUIulYYiYzRQWqKQjzoeHhuIEBa2Gykmvyepmu1jQYElxSAf2Uc57rYByStU++w3zOGIB9pNpAMmCDH+0XRb6LP2eek/NHhrKl8ZaT2rFAYYNKXqyYpdfkPY4t8zwAROVzSE2eckZhCp/F0owp+VjOI3Lz3p4uMU3tA+W1hscTex5rqbO7S3sYQLuuro5YpTC5sR57d48obh27fS1ee/mZaG2qi4WZmRjaNSATcNZwXXN77Dt0NK6PjsbcwnwcO340bl6/FvXbO3Hs6CNiT3JGj+wZjp3NjZibnowTJ09EY3NbfPzx5zLiXt0M+ThIhjrqVVwnbkqQKKxKTLQ311ajv69HPjzcD3vP5WvXYn1nO5aQmNO4NIixR27DPBbIrqkxFpYWoq+nR/m5gXXk4HhXrNkjqkis8Z08M/YWMxQdQzAfaKohVwiLUawhwFICUjie4B6UYpbklhYhTYf0q6CJS1OIuUH+zVmzXd8kxrBi5LLGYdRxvjM/8JMwc8Iedcs01JEUQ1ZOtSTi1HntldqFAQA02+QY1irjuVlqW1rLK8uWX2RPKHWr5dU1ASokLaXLr3rZVQKjsi4yJnrw91nAf7AhUfu6/9q/5efWNhJqGwYPaybkGq79jvzzgw2J2kbFw14vwFAJuGsBdbVNmMx1HmyOKOetSK56b6+9n9r35ffUjkWu3QfHR3LuMEwlHVofRw4flmoKsVt6fApsXOR2ldMV8JVA0YVdzz5BviBZr7JXEbewLuR7Vg+zcVVxVyplVJi+dXWq7fDD5xOXMh95H/dss+wCRJRvSqe9Yos3LNfQ2d4h+VnWC/cjOXdJRfO93s+Qsn/11Vfjy7Nn1eym1inVmpUV5XKcMeTD/HCGcc2A/qhRZi7Kd/ft6v26UfGwCf717/64RwBGBYuBBcVGzmQnGEv/AYoNHNqJeFNiWWi4LH6KD2lcJZ3cGcs80LUnMQKxoCJUKVhR0MAAe3CgX4ckaEaCNrrix48f1eF57+6Y2Bg0JdS1XLbMlChgHRR+1oUQYcNQooUWXHubNYa3titmSrAeQDX37dqljYDNjb/zvZMTkypeKPDk9/2D2gBujt4UQ4QkN+WUQPI1tWLO1qzfDQ0MxtUr10wPPXpUBzjjgL4o1yM0K6iw+YWSlG8J2UcCQMBIgYJkFTouY0MjAHYDSSubH80MEJpiYSBltLysgjkJJIEW48Cmx2bGa3kdRTECRZlFVhJ5d3SR6pJBLX4Zs7OS6yCAUUJTkM4EbQR2fAcbMxRMCiBZPBBqrkh8GBxlE18lAcXEWz4YxUybcRgZHtH9simDPBdzpxgE2RyuJRZhSIDeLsEwmzfPLQtcmKbqIIN+jKwNB4TM8qqFnErXvZjaEiiRXDBPKGCIdbK5pftT4bAkHtL6FWLD1GI0xCWr0YP591zFNFWmfchFrK6oyZQmxqx8ivo892RUKDlLJHI5NK3tD4rZiR7dcJ5THsyJABb6pwqbL0FTCZ5K8FfbpMid5z5WgSKEgioqjIryq8pGJfQ4jYhiSGfZnftR5jZUc0EcREttsyRjURtE1XQqUoYmg7oS+CVrRcltgwu2jKHklwoSnfUDPdjsEhIfUG9Vs2MXvTKp8XV5gEwnyeKvNCdBnqvYb0QfwYFMSGsMsyiqOtHbERMMELYCkMVi3CwWmL9DyXCZA6atw+ZxwpMBoCnrLubIYJZEobVFQYmS74JozwYi96PXlyKmkbhO5rJImImzCnMPmBZmIJhyaBRLXCC0fJDkgmp0OZnfjClFR/lObIP0dAGdz2dvUqLfYPk2qgVOfluVUIvdVvYnCuRCa1YaSmajSHZgpy5m5+e1LwkNriKgiwz8JNIzC59+hHy/i86JmGM8KKSxL4HMZ7wI/rTHFRqy7knFb0vYObmpV7GUZw2Ki8JksgXVyJAcimew51eRXZJWsrX6Wacg7Pg3GhUpO5aNmmxy1AbYtb9jb+McJYhkb+Ys4/4Sbe2iiaVVPG6WsCDoJSjdt2ev/ou8oVDmog7DkKGwYYkXxsBo+cIG0lzaVEGD8QZVz39diJSgTaE12zjaqFcKxn72btiAknMzYG1tRY0JjQlSEAODbiajEbuKybZlgCTz0WTkz8rastDKRi55aVaLIyS2xZen7E85z7PYxOvTHwj2ToUukE1bGmhd7fJYkM9NYYJJNqQgndh/2ePVXOcs4cxpatJzBCErVkO5OBVVGzhX0AVfi+bYjpadiN0DLfHy80/G0vxssHWfvXwjJhbWY2E9YquhIfp29atAa7PLLOQhI2R5LzemXEjkDOLPJNrMrc1tCsCWlQPpDr2bsQQUkDtp+nutb2zGwf37hFi+c/uOkNsUu2meoK3PZ6Ct39nRqfGnCCD/sElLRaZ5K0X6fMbI77D2WOtcKw0xKhKZPCUCmfjCqHz2QWj1RhyDamP42CMoEhC3MLs4W2kKUthhH+L1KeECY6O1ozNuIo9RfHGyIWE5D7Or3NSk4VInvzExrWBnkhC2thWzzA15g83Ie6ZZ84CYU43QRgqqTdoz1CQtc1uFlg4kNVa1XyhWBPBQfIgsy1NkLEsjGzZFygYyVnzn6cdPx7vvvVeRpGTvSiPFBNtYKtFsRSewgEtAAZvlwFxboaFBA56ZTNGnviEWFpGNqkrkCTWHt06DC5rZqKCxxXiwLimuIRfED40y4hlYFBS0YcPRPDKTBoYujK6m6Ovti6WlBTORV5Z1xiP51NnZHXMLSJ3ZHJtGA/fBXiXJvbJmbQBJrmAZG9aBZEoVt07F4cOHorO7V+9hz6H4x94IAGppYS62VlZiST4hDdHbVRffeOnZeOTYwVicn4nt9c0Y2LUrtlcpAu/E0tpGzC+txtLqRjQ0t2gPYh5QXFygGbu0HDdv342t7frY3IlYWFwK1szK0lLsG9kdp08ej57ujvint/4pnnnuGUnO/vSnP4/XXv2G5s7b774vHwr21/Pnz6mo/v3v/3n89Kc/jbG70/GXP3gzfv3rD+PGzXvx3//r78fVq1fi4uXL8d3v/mn8w8/eivGJWRdwYfuRB9XVxQvPP62m2JWrVwvIQTuZnjP73Dde/kaMjt6MsXt3rYHd0qLCNDEK4403HhI1ajrQkOHcLb57AnoVLyzVeOvr5SGophHPa3tH7O0LFy/q/FhYWvLcKfv9m2/+abz33i/kg9Hb0xdnz53T2bp/3944eeqkzpaUocrYhr2CgghrhwZoatxbagnAhhHSatrVyDhm8dxNA2I6N0DF5uaMLgboxAxZVHP+AOrUHhac45KGQp5DiPEqo0Nm2fKxsD9F/j1RtskSrYIpDDpSw0H3YlAI94EPjrTrKYgjS7VTJ3S1Yg5kFJcX9awSDc7zrEgNlQJ/nneOy/Bno7FjIIGi04b6aNa5bzlR9kfL27XrdzT/kB1LZgVnxZWr1+WrpPhIPoUdiincZNkpDHgXisXmJTcENKUzB5mtdc0h5o3BHmZdJFjBBesqWzIBS9wDbADiFs58NVC7uvRM5ubMmk+wTyYVKtpRUExQHN4qRT4u2VfZdBBwRzGYgVaK2Ivso/0pDI6oVLzVaGrRX6k9iFlW8hIKzKy99HXi92rkIHXEuinjAECR+8HLiXOS++H7OSt5Tz/sXfwUm5picmJc44eMG3NuYmw03vjmC9HR2hDzMzPR192ja7hy5UbUNbVFe1dPjN65qzs5fPRwXLp0IXo62uPokSNx7twFzc3BwX4xIlZXFpUfHjp4JM6evxy7BkZicWU9xienYmp6RntYR3un4nfOKhqo33nj23Hj6pVYmJuJpfk5mWnj39TU1BLj01MxMTsbja3tYigwv5FfFQC0oUGMOeJgfNDYZ4hz5JO4zp7faXBPYUbQbGA9KFZg/he5XcaXugzPhn2/TZ6llt8WELIoKHC99quDubAjZoUUDwqLmYfc2t4aPV09aoIg6wr/Y27O8uKwDlfXNuw/UHxMmAuwXpHkYv4zO5ZBoQuUVC+AztTMnPZe+RORx2FIvhOSS+xEIlO5m/MqACnESjJgbnIzEEaFms0VdvjDGxUPa0bUFvizIF/Jy2uS5q/6t4c1LzKvyNwoGwEGRnh9ZFxdXSuV9L6yfqrxtVnkD/upbUTkvWSjOv+eOW5eTxbm9d1llTL6qRiR6zaZ41Z28DXknpP3Xfv9eS+V88CvltSogFVF/YG9VcCjlOWm2VaaxdTudF5R5Oe8lD/cmuaqvSbsv8Ley3og5oHlRYOLGM3S05aR1Brp6lKMyRomZmAvdX7YZcDOhlljxOXcL3VJSY+WPJV7oQ5I3JLjmbGmwGawfsR2q5P/LqBs9geu/dDhw3pPSr/yuZxB1DCJvZCYRZlmfGJcgBbqY8jnf82oeOhU//qXf8wjcKyDoqy9E1iYVXOkHSVKNtp2cSTRcASvlSZBKUiIKl4osUnLNKUXBG1SqlxUbGpocuCD/FBza6xvrKrYTTeQRSlmQDFKI0hnQSP/pE2jhULAugI2FcCkI2q9fBJeUdGLJAaHGQs5kUCg76DCgvYlUeBauCcWPYGZ5FIkAeIiDpudCuiSCCFZIylpiD0ju2NyakpFPDqsjBGbIN+L/iWyVInkZly5B5o43IdkloKDtyeug4YAHQBygNd0dyvYsya86ZQwR5AsosBGIYvggSCXoBSEncy+d3ZsGiYqGVqO9n0AWVx7IGhMQaGUDnjt4cWz4PW1ckSVg6MUxpSUlQK25Hso0hQqtIJgJe6WXMo5gyYxRY2BwUElcNwnCD+KL5J4ESqmGPIWyY5E1siQXF1wawzyZ56/KL0FVaNCaDHTJbkmUEPjF9YL89ramfPR2dkuBGkWFEG9gv4VzW7VDTMKTS78Gq3OwUMynwU25jjMHRIDXmtkOEUI0Ltu3PDceSZZpHIxuhjVFrS90VDl4C6F9gwCkqKocS2F4AcDHyV/pVCfh5/YBkqKapKoAlii+JyHvxNQm2VWkN36cie+XCvrhkI0BzzX70DFz4gfI8xrGR9GWHMtXLN+ijlZBlXsGaD0ucD0oeD7k1HAvwuFJVNr5qivh+8Uq0CyIFXkhoO2KgrEyC4Hq4yN5TMsxUSBg3mXiD+CbhU029q1D5AUqFmUBtRF2iv3jSzsCvVc9Czt2YMJsBG8iTJnD0gpNFHYS4AoRAcF9oLgVcBZkHBq5GRQT6ETGZ1i1JXBIPOfIlUmfRUWTHkdQyZfGkkquamTKJcszBJsqUEm6a0tNSxZn/zA0qJIQDGC4sXhI4fV8KWQmQjNDKBBHfOZMpVn36cIURCRYnSowD97H9XWe4fXqtCEpZid89L/ddMiGzh4BRG0sb/qbCkIOr4vkVwqjpRnzvuzgcKcR9eTYI79nB/uXflI0d7nGaiIQzFPhW0zD/guCj6SCJorzIRk+tQYk9+3f+a8jx2dCRQCofGyV6shj7SECoxIcrj5KjmycrbwZ34PYogEeX4OI8ESgGPeDvtwx827svjK2nShwp9DIbu9soZzr7MEmJtqzGHWGWNshp7nrxofxXROzQoMfFsporUraKaggl+VCkCFrWNWlgvu7Hk8i0zIsiiS+1ruA7lfPZio5B5XOx/uT4w8Z0B2aw8reypJAwhrzhgxCKBZ0yBEagvggHwz1pxMl6yKMSKRJmlPmQ/+qbluJxrWN2Kgtz6ee/JkzE5NRF19e5y/fDvuza3EOns5TbpmCk4NsbNJY6UURTo7yrzdFtsim5yc6Xw3hSIK6FyEGlTIN25uxMBAf/TvGhDCWayXgubXObwTMTQ8KNAA5sg6KoqHxJ69ls4cvzeumEna721timMwPJVkoSTXkP5ZrKiy536ODARz35IIljZMaryQjB3tFelMzrrcX9nH2MMbKSrIy4xCJHuBvWf4UTNWsYd9q9QQbWiKsXv3ZPAs34iUUlGTBCPCxmKGzBlPUQrN/Q4ZaFvT3nJk2aSkgGhdeAzNKZquyUxbe1ExWDx18pQKUFzD5UuX4uq1ay7gad9CcsrybwmiUZOmNAUdd/hHhfaenjh56lS88+67LmAi4dmK3BZyojQhk7VU9QPyZg3Dy59EcSdNt31++IfnBuJdnk9FDjXlC2GuwUJoIbEm9pEU3Kp0x5X8E/eub+g+YeI2NDWJ2UDcwnpmTnXC0gAYwD1vV30SaGZIi3l1rfiurMX0LIWw9I9hLdkjjs9hreRP7sfpteS47p4KpfIOY84vLUZzK4jItliYm4uR/r5obYjobG2IkSH8g+7F66+/rKYFzQkKEKByaaqsrm5E3+CQQE0UnwDNKB5bXpZXRXN7R0xMzsT7v/5dLK9tmAmgfdVRwGB/n5pZ3379FTX5Ll+8GP/j//Q/xDvvvKtGERJJ7M80z848/kT0D/bH3/4f/zGeevqMCoz/53/8v+LM4yfjxIlj8c//9F4MDu2qaEjXNzbHRx/9NsYn51ToAsjEdxKvHj1ySI0hGgjE7/ze5s8umICKVGyCtBhyWIsLKoRwhlFE5T2cu6wt1lE214jZGPOjBw9JFmp8atLMTuR1iFe262J4cCCef+65+Me33oo1cqgsJBVW3V/98C9lQH5n7G489ugprR8K4Zz3FFIpurA2JLPKMy9oarp+MqVnLhdgQ4X5WzHTdnGZma59t6C0EwDHfJcvBwjvYn5t8BNN3OYqa0osK59NYjHDeEeqrrA8slhH3MXZw7wE3W5fBxuP02SXFGFYikx7rvYY1k9biQU2VciWvwUNlx3iFrP7U1OfmcRZ7sYgEl3WRie+m56eKuw+S+TybDIHZk0oVyu/E2tVkju+F64rPRfMNtkUMIS9jevlv8S2swsw9cf1WdwYQDYKyZx9kj/i/E7ZlfLZMKloHCJJwvMwyxyZwoXSVC+mspz77C0FKMIel/EA70MCiYa5dNsB3wAsazLLMiU7q6mLwUwUvolB0z8kAU4JpMqcLROEjAGyWeUzxlJ5mTP5mqrAJCTUiDsYE/Y43iPEc2HF6hwrzS/22mSUDg8Na00BSuKZ7t2zW9LVyBWxDjiHpVTQ1yfzWuoRMLj4t9Frl+PN77wYj58+EdOT47G6vBjLi8tx+zZNo+bo6RuK6zfvRF1DYxw+diTOfvH76GhtjCdOn44rV65rjgEgQfoIvyLW9GOPnY6PPvok9u45EAtLq3Hp2rUYm5iO1hZkbDg/C5imri5OnzoRTz/1ZDTVR4xevx43OMfkP7YVSygDrG/GVn2jvC1gEDQg+bQF+rtFgBViNwCWyGOzXjgLyLeIj1V/KOAU/aHkXcojK15fFIULMIu4qzCXiJ9yjvM5qGk0N1r6G1aV5EbJ00puSqUZLJMkndpbtSdSfOYZaD0TsVCjMOHbYERk9Uq9wmj2pujtsrwl69VeqEa8c2zhV8QeBQCNtIw119beIcZiFra5VqShWZM09ml8KB4TsC6lydxAzTlZOwc9R6u+D5VD8Sv+8GAxXu9XXOEb5bOYs5mnqJko4IbnfcbVyfeo7TmkcXxet2PmB+GDD7+wzOcy5q69ztr4/GGxeu71lXjgAcBi3mPWGSS5XBqsVkSAPW+2anpVJmAlQaganXrHsAB3iaN03nE2lb3e+78VORg3yZ4X1YWM24hx04tRTe0G6jilhiSJP59X6c/imBXgGEwOFDcsz6t9hSaYGMDeq7Se1Pw12EdnEOxKzWcD77jPrKdoHhXWcn0dNVP7OnF9x449orqS/YXcmCe3oiaIag3jw9+72jt0xt6+fVs1SJp/8lHcMhDx60bFv7Qiv/73P7oRONreZTmdYvTLosjFn4VEmTZLpoKNpSHmF+crAV8WN/LAS1QxgSGbWWOzEV1K1IoWNr8f6B/UIWXdNzMBDhzYp2Do5s2bKiIjo4SEBgc7xW2SoJHdu4U+JCmjOEEAtbNlKQAWLZ9HMZnOapoc4m1BsoKME40Lkq+bt0aVoLEBcc0Ed2yGNERAJ+3bt1/arSAxSc4p7LE5cT28jqCHhonYCVvbalxI+qClNe7cue2gb5tg2CwJUPory6tCGlNMUAAEy6NsYowPn8trKVr09++SvNP4+Li6wdwTY2Pk3pI2P4IrCnkUtUh2k3nCIcimJi1iQ8B1cqkQIVkEJ86mbqINaTS40aEuBitgUFDoZkctEry2w54Hdib7MnrFdBPvjvW1EqBZR5yCF4dOmvS6EOyggp+KFEyRd1BRpRizcfjyXNwcKQFNkc8hgYbyTCHXEicuYLsIlShSLgAAIABJREFUYdmEzq4OFaY5/BmbbM4xtgRWoBCzkGddbi9lGkCScRCCy+MPSom5x7rh+fIdmNaquCEpIRImj3GlWFgKa5UNokgZVYKFCjKhPKdiXpiJhAOQpLtXG1CJbkpmQaLcFbc1GC1v5oTlk1LCSW2KSnG16EmrD7FjRpXMxm3WXpkHxWysUoDPSk4xsFMDrOYzaZuwZ5D48cxhvgjNpWLRRrRJhqgc9tIttoGhGyI5R22CpmdKQl7mY7VIbGSWf4xedBHT85B1QYMKtgz7jJEXNo4n8KVQAAU054ySxDJ3uLhkHGRAnoEj80aBrKA/DuoJvDPYYizYZ6rf50A/i/DZPEiJLSORnCxS2NY9F/SbDe53VLBXIb5ogivQRccT350A2WTTbiXGBX2jYhWNp5LwMe6grs36cdJKcWJiYlzv5bp4z549eyvINBAqRsa6mI3kjpCXmBiWtUsyJsTTzo4SSAWOrBv0cNWA9DPKBoPmYiUpsHZ17Xrh32k20rRxgdxm27zH6Cg/YyVCKjDAeLORZwbvFOxAmljjnyZRMYxWs81FyTTTzTnOM+Be2ItZ1zOgtbiHGqRfvjbXcu06YkwpJrLfcWYJkbyxWUEbZlIldAw+EzQeMDItjZCt9Y3YvXu3GkTMA++JdTbQLtISNJRzf+LehRpVAXwzenp8Htmvh+dpJgrXxdxkr6y9VzfmzU7LeSP5CVGaXVDhrAPxKVJ8YdrwepnZFRZKFtGzQfGwpCe/N9dAjt+DiVzuiTkfPL5l7dNQaDGYQahbzHNhtG0hZbaqea4mfX1DdHR1aM2IvVPmCmch+7dlLdm/PWf5hkYkD7Y3oq8r4uUXnojF2dnY2GqKS1fvxujEXKxxdra2qKi7MLcSy4sr8hLY2PQ5Nzg4oNhFcQHSNJNTsWfPbhW5iT9AEOqeihQJawR0FOhm3qcmULjgJV3zrc0YGNil+TS/APPBRTyK1DAxLK9lFlV7C8Voe1UxbygoJWKbo0jrpDT92aORFSJu4BnqnEW6RWhnsxUBA1C0SfN0FRXq6nUvfLaegZiI3D9SDNbwlZ69zLBtXiiZEGgp9fXyA6AoChLU57rnU2qfaz0g4SCgCSyGjljlMwtymr3fEpHFDDflTyjwra+qEJqNDNbdyZMntddx1pPUIYmifb6G+ac9qZiEM8/ZS1986cX44P0PdN5k8ZFm2GOPPRpvv/NO5dxMoALzT40UMV6rcihqRHtX1f8XA6QZTxAkMsyecKPeBss8T/YdUH5q6PK8efe2GxWdNDs9SdSEauvsMGNP26IlCvAoQWbA+769imgiwTTm83v7uhTL8nrHbOzXq5Iog/3B2pmdmZOUUu4VNMmz8c81ZbNLMUZhBvI7xs/5wFasbtj3pA0pBHzXaFZtbURfR2t0dzTGc0+fjsXFqRgZ6Y8eJE/W3cClKXH10lU1A5ELYx7gVwGghflIzAXacX07YmJ6Nj749Scq1nK68h7iS/Z7ZFtuXr+u4tmLzz8TH//2N7Fv/36Be2io3Lx5K/70ze/FZ59+obX3N3/zr+OTTz6Py5cvxw9/+AOhom+N3oj9+/fG3n1747e/+VRx+J//qz+L69duxr2Jyejo7InmVgrZoOcbJe3Ck+GZ8GzZezKeIDblue/fvz+mZ2akLw0pk7hRRfU6FzVefPHFuHH9uuWdiI0KYpPiG0jrF559Jj7+5HcxNQu4rEHNBU0JGhUD/fHUU0/Fe7/4RSzCkm/2GUdxngbIK698I7788mxcvXZd5wf5Fmzzs1+etVSjCkiOPzOPY+/IZyzmUdljOIPIRxQn0hAtc1NxVXu79gXPD3yBYA80Fx16rwXnFenVZIAPZz1rkXOM77GMX1WKzPPVxU819WCFqzDkgqI8NhQGuvkueY2iPT4yNGRWBHmR2KsGhyUCdrN46/G8bEhtPybug3nNvGefsu8ijGgD4oTObWpSA8pgGOfK2UTRvcjnzXJYsE+Ic/mzgDZqTjpHqWUTcE+whASIqm/QM+RMFiAGwAbrvcTp3Cc5IXr/7FcrK3hDOR+xLFidisGFgGiwmfbkspYVQ5V4qsQYyISRHwu5XmJCxhimucc047lqQ5f4LxtT3B9jmflG9ZmXuL7GmNeNmcK2zKDAnI1SEIbZRdyyHRtr7Jf4rrTq/OYHD6+CQVAdI8dHjewCZBweGa5IpeDbMzI8JOAAygoULXthfBX2wd2xMYEiUQTg+d64eim+/6ffiP17h6KvpyOWlxfjzujtuH5tNBoaW2NoaG9cvnIj6pua4uCRI/HlF59Hf2+n2FE3rt/SPKdYrgbz5jrc1jh+/GT87uPPYnhkbywsrMbFa9diYmamIg1jZjQ+Rs3R2twkz52nzjwRw0ODce/unbhw/nzMzM7F7OJizC1vRFtXZyyvGlxXv+O8uRsZK86aBoCL5FZuXDN+8uss9QTmrNjINBMFICi1Hk1kH19iWpAnFdAar+Wz+SyeOZ/H/OymUY2u/8qyiqrW7zfAgr1MqHWZfLNPtEZLE2A/F4WZA+QaBoPh6VIwOWq0FrP1Ik3NvOb75xcXBapQQ1dNDV+7gIAJi9J8dYOEOg8/7NE0t+/evSevIyQB+a/nYcmVK/tU1U/wYU2HWsBSZfrW/OGh/15AWV4XBuGIoVtkVVnzbg5V5Z215kozWNtcYW8l4kGRTUV5IXPih11RtZbwYA7zsPur/YTaBk0l/a9pUvjfDRbIH0sKu/ZAQ5gY0T+eXMpzi5RYAvvExkfqM2yKzTpWs7Xk2jxzAdZKXJC1GwGhy5xU44Jcrng7cP4SDzmPKWcc583Whi4lQSucWY4zLcsoWcMtf1bKJqsBXhjgxOlsm+wrXE+uMZ6pFUucV7M3c6YICF3kSa3kMaX9n3j12vXrqv0R52t+y+/KBtxa0z09agYyJhPjE26EFE/Ojs521T2/blQ8fM5//ds/4hE40mZKvBaj5HEsI8APyMD0kOAAUxcf9NrmhqjcNnSm8LypTYTFz4HIgtRGq2KszY7FJoCO2GRTMjYZOqQsvtRbe/TUcRUaKIpduzEajz/+qOiwly9fiZu3bumQefLJM3F77K5kkwgaaV40YVpY0NU0EpQwbm2LCk/B6MiRI3H+3Hnp9p46fkII6rG7dyUjRXFfm1n/Lpm3kiBQJDh+/HjcuGE0hILm7c3Yt3efUCOgIym8cs/HHjkWd26PGbnW2anGhXSnVYDlv3W+ToLYkiyS7Ft7bkEFFDYxDtnh4SEd+Ddu3Iz9+/cp+AdFQ6LN/fp1mzG/sKiiyK4+kDMr1gZfXlEjJhERRoE7sEjmCc/DUixOiio6sxQba4r71nB2s4Of7CazkedmXtu4yCKiAu8waje72aDEhOhYWIj+/oGYnZtVMi5UA7qaaoLYVLZSrCv6rko+siPdbOodv5N5sZD2yPdYwoIxzfvi+2FRMAeR4SJJIchic2ecSE4ykVRgj4xFC0lJmtjtWPaojIFMtwryOFHdNKRk4l4MuVSQKYZkZgWYxu4Ct4s63HMWBbc53Eq1MQ//CoKzFPxT/iqrkgVocl+ikA0K/psFdgc01gaVh0jp/tcWAN2oKOFCCW6s5ehgNvW7Hfy56eMAzu/Rn6tRTuWD3Dbw9/Nf1g+HtQq9+LzISN46jTQc+fzenm4ncJIiMkrbxZ1slt2f3LhvWopVMsurMiuk5V5khFJSy4mjdYrzGbBPiaFBAbMELhkIKngUe8ooBX6EtgWhhzZ6KdzkmAstWORDeE0G3fZdcPOGgFpo3fI5olGj61uSBRmsV0yaXTB08dlmpYyA6K7Fh4K5bfkeB0EN6HRLisEFXBvCFyYBLIsie+XPNMvNyEcXiPJzZOAHuhApO1Cf8qqxSV59I2w4U77FumkoBtdC36MJWoqWfAeJcGE7VFAuNQ3PaqOiFKFrGBXScK6rU/GXvRO0ce28SBo3v5P3B6jVNpt1M4bsvzQpWJucJcmwSXQdQhIKZsWmsjRQNooShUxAyPug46cEWW3TVuNR1tX9x7/nOGg1mszyBIG+i/dA0cYVUrMdDxCz34QGLAg2IGcUodnzOQtADrpsYvN2rblSpEnmn/T9i6QFzW3OGRB0PFf5T4CQLeie9EBwYcemoswNzpFsxukrNt1cZi7RlE1zTdOql+3rI5M7S4pJtqdIAWYxs7axmo3vnNe1e9F9+1JpetY2f9xEdFHVTDwQsptKDBi7kcFhrWPObqGgaFIq+WlUQT2NpY2c2lYxmsJfNpAYXX0eEolrS9HevBHfef3FmJ+djqnplbhxayZGJ+dju7kpGttaJG0zMT4T60jSIM2zvaGzjSLolatXKtIbrFt+ByuF4r7NtK2trTMK7eqRkeju6hG4gedFIcaIUK9rznk8CPKsEGNK2rpLlb1avjZCP1uyA0AAhXkbimIYuaOijOjrTU1q2LPnXrp0Rcm7mqllTWQBEfQ957SZgfYpS9YFn6kCHo2hJgNRjIw2+pXPoNitpiZGnewxLa1CB8NwAvUlyaRGival4SsPFxdQuN621vZoaWqJzR0XzM1YLHFL0aWXxB164hSGaZyAOi/SRDLoLKCENF9lvyMeoelg1qA9YWgqGcHueMcSdiGZJu4bZjGyLadPPxb//PbbFaRlzmnpedc0Kipzt+z9Wbyk+cNn8d3E3JIzKeclSGuugTVHsx6PEZ49BtScPJ2trZLSELJue8sN9mbkC9qsSQ4rbnYullZWY/++fcVQd0vMMOTvkOmSZBryT7t6BawB5DM/txBHjhyN7t6e+Oijj3U1lnw0QxFZKK6NZ5rPFmNafrh/YuEsDHDfxEQwWlvb0ThvlIQO50Jvd1csz87EztpqDPS0xA//8s1YmBsPjsN9hw7Gxvxi1JFx1zfGzRujsat/IOYW8B9ht65XMZL4WuzQxoYYHRtXYem9X34cjc0NgU59BznJ5pbOizOPPx4H9u6OD3/1yzhy+FAcPnQw3n3n3RjAi+LMmfjxT34Wg7u64pvf+mb86Mf/JU48ciieOHMmfvnLX+jeyDPm5qbi7X/+MP7sz17X5/7jW7+IF154KoaHd1uSpw5PnrWYX1xSPIN0DN8FIpIYU40KtPdLw4ow+7tvfDNGb92KCxcvS9qQuMANa7NYvvud78RvfvuxmtweY8daaLC3tXXGU2cejwsXL8TE5HQ0tboRQZG1vblVjX10vG+P3Ymevr5obadpU1fJWRg/TOWRlrp9i/2hMZ599hnt/2fPndVaoBnCGc8e48a4GbDJZlX81orRbatex72x7oitiBcAn7nQaIaiGd+cyWtidnEGMs8lP1PYBPINQmqmMCUN7nC0y/0TuytPKIxUD0wVkawiTgFMAEZhvIjpyZ34HvI6nhPvd6EqLAs5M6s9kntifuUZqfy1sDoASVAUUxNTTXHHkMQY7HnEPWKDLeN5h6yMYzDGxM+9FPXrfIY9WFxMOVhLxgGcsPykZFHrYH1Zmod4psLkYI0K1OJcLpkgsO7JY2nEcW3EcPgm0lSCLSAQU9nHdZY2mglL7OBmpGURFXv19mkesz9zZhB7ck3yrSrM+gRBpIyTWaOO+cn1HXdUfzJ+yr1DskE1stDZsEhmXoKHeB/5s5pIkglEehT5WBuuU4/IHCeZy1yjJEB1PVuxt7BUZ2Zn5AXC3krMQ7EPGRexmiTh0qGGNvMbkAH3OHrtavz5916KrY3lOHRwXwztHZFM3aVzF+LmDdbaYFy7PhrtnZ2x//CBuHjxQrS3NMWpEyfj+o1bOk9g2NJgnppGcro5Dhw8FJ9/djaGBkdiYXE1xiYnY3GF/b/TgEIVcEGH2wEHfwr8aJ568ok4euiQQAaXkKK7cjW2GxpiYRkJYiQN16Ot2aAFivUqykr2E7S55T+5f/YmmtLk15wDisLLujWQsEExIPue2IflXJfaQ/GsoYhrGVjnjFxzb1eHvYmKjChxomTHikffyhrW4QQ3Zld0dQDmMhuHOc53M+94rvquUh+wPKgBlEhctbc0Fi8Ay53x/TY9drOCOHFjbUseScxB9mFJhLc06hnzHmQOASIh3by8bANkIPMGpxkMmTWJnKcPazr8v2lU/EG8m8DDAkhMkFoCStyoqEqo6v0FZOp6S4IxC8O4gIkfQmy4Pz0pYLTaXz4YaysmqWGT1IK0KrWKkmvl59QCMqhtaN8rSgG6Xu/mZR5Z5lisvJITVljvpd6gRh0qIu2tmhfEcoB61ExTDRHghyXOOM+YP2p4FUUSnh9rDllQxS4lL0z2sWqEMG+lugDrekXrASBNeh2RC+eexX7J2cIP+yDjr/i2NFGy1qbGcPG9JT4mN2OfZb2RC/LZYsWVfInP41qmp6bjueeeiy+++ELgOj7nwIH9ej/nJmeVcqCtbSlEOGbl+uriyrWr+jvSUdNTU183Kv5gxn/9iz/6ETjYima/C+sEiiw+irlpGiZUfkGGq2Ap82FLWSR6vVJALoVty9e4wOk6omlebErNTab1s9jXhQBwJ5LPAOEj7ebFRWl6Uswh4CS4BLUktGspHKqTiHkziW1JLPkOEqWZ2floLAUYmhRslBx6FEy5fpATbAx8BwE0aCNQ1ySSBHTygBDbA1oXhzGB8o70I9kwCXqQZGLjoTGSQbKNpesU6KipsOWglcSYJofYA6VgzcaKQTiJdurlw5CQfnkpjHK/NFv4H59HoMyBSTLLgYYMRprIWrrFSEyNvyhw1n/W5trcpGIEG68TbCcGFXRciSgtTeUf07RND77v9/o3B1MVKEt5j1B88o+gsbPX0mGFGs21cMgQLHKt0gwn8Gxo0nOkcCf63bYLEgpIG33dMj7W4ejAKbvlmVQwbwm4eI+NmU0BpNBLApc+HRhOMpag6a3DvKOAXhIg0PdKwUfU9cYGzUUVNRpBmbbp+aSni9dFhZCp4h1zhkAw0VKW0/C6omDG3PL7LTkh1GVKOdV0DsQcKOsuOwoZEGWwkGwK/V1odbNjmOOWlalhVJSHqqSioGTy4VXQ2aKRe8xImIyuMdqqUvQvRfw06uUeapORuhJASYZHRVKzGnI9MDfMSHETjx+j2m1CqjEVxZJAnT3DyNLqvVcNxx9kV0haqBhy8zmmWZJ4leATen1ZzzwPI3jdqNA8rGFrKEgsRXAFbjXUfgINikxpPu/GiNkQblBZs1/Fq6LVq3VY5BT4LOYfYyjzWSG+CWBsKK6kH+QtcjYbGwrIa5s3bhgaceNg1kbWQvc1NAkhosZakUHJhJDxSFkq0N3JYEp0XyJwsyDJNRAMJTqS8WBuy2ARH5kdo4T5fpp5zAMxzdbXYpoigOSGHOzLTwFUVUFuJd3XBbGqZFA2a5g/FOwpiluz22s+g2gnTm6LSa6hxcahiTjkdxQqYIrIYLN4AZGL8Cn2nbGvh5BMQllZ3kTjBDoRPx3MtMUE9N7+IBvgwQBADbGWZgXOIOo9PrzP9F6ukb2FsyYZFTDvshm1sWpUtdkKFFOtPS3Ee1lbkuhT49TNw0QlURgYGhrWekL+hzmu8S0ScOzJDoyrJup8BucYxWiPLY1VDBm3xKJgnxJ6KELMlnx+2kfKnmJvAe/P2bzJZ6VzpIYJln/Pc6h2/DJhqk3q8vWSxioUad4rxmQpbO/V2boj1gLjapDEjvb8pRW8OnZkdEvDhfFkfSFtMTU5LdYjRRnusQc6+NpKtDasxnPPPBobqzS11+Pi1bGYmF8Vo6KxA0mI4ZiZnIulxdVoa2+R7FBfX69AG5IkAOG/uqbEKhlENMyQmmgqsnOsIc6WvXv3qnEwenNUBblNkH2FecXcHOjvk9by3MKcmg0UG0A5c7ay/mnOSLZgbV3NehijACjujN1x4VCSRPbQImGiaEMxlbG8cf2GYxIQ9uXZM46snZHhYcuVqQFhJDX3AvIahmpKu7S2Ypy87GZGMbJmDQmx2NisOSHgS0NDjE9MqmjR1YWppwseQqILAQ1bwoUG9lb2PJpHO3V1An9wjqQ5uuYwkksUl6Qzbx8NSQVy7pVzlII698Bey/hTwEvkYrKD1QysNLDNclJzsUg/Eftx/b19fXH8xHGh1ZlPrBGhkmvMcJNRUTuPfYrbD4cGDe91o9ixWRri6oykicV+z15atxPTUzPyWFheWIlO0KBdXbEJIralOeYWZqO7r08xBXJJI3v2xOTUtOQ/jhw5pHnB97CHgv5G9rR/V5/GFkQ/4wkKHLAA845Crj0zGizjVtiLlkFwIT2lFGuZV4xfNmq4b8BEsFcpdM8WjzbJsTG3lxZjdW4mDu4ZiG+9/lJMTdyOtrbGQD+eonlDU3PMTc3E1ORMNDW3qRhLMQwGha5rZbnolO/EwspaLK2sxc3ROzE1t6A/r0m6iP9txO7hwXjs1Ino7e6M9955N1566QXNkw8//G28/vqfCBn+2efn4s/efCPujY9r/dEYP/Xoyfjxj36ie/jWN1+Jn7/1i9jYWI4f/OD78f77H2o+nzhxKn7+T++pkQLqV4Ut1k19fTz/3DMxdmcsrl4fjSb82oqUicxe6xvijTe+FefOnY87aNoTF5dzgbVA05NiBWuXNUycxJgzvpLdKuwICiCwaeRbhL8djJW19dhYW9Nedu3mDY0/kiYr+CvgM7i1Fc8//1x88MEHYlFMTU2r2cFZ//jjj2tu6jnKL8CxBPGsWdglVi0xFU1R+TXADCjyMI7fLSvDOZoMLWIKniOnvJsxRg9XzocavwIXCH2sZGHT12LpYcnMlf+RM7CG0kicvd2MJcesnT1dsbTg2J3XwcBnP6CATpOXvUNrv82+RZwDeb5n4175blm3WbBkz3axzJJPzhMBd9hwmPNTfoKw3VLWqUjrqMleZBP1XSWmJHpnj6KhTTzIc6B4OnrrTly/ccOa6c0tYv9N4qmAvFZzi8bR/jHk082WxW1vF0CCeIIzjzXOc2GfSE86gc2IU9XQN1NpYLA/Ll68VCkwsm+grc6+wOt9FjTE/DxxncF1BrC5qcm+m/KW7IuZn7k86Z/aRkX+ubYZwWcZCFbNKDKeSEaF5V8cBxKfsRZMKHMwkowK/s6zTYYzwD98HAGuwQhGUpFnhMcOzRz7TNpbCa8l7gUQAe+/d3s0vv/nr8fd29ejs60p9uweid3DwwI9zEwvxPTMfFy8dDW6ersDScaLly5oXZ4586TYVwIhjuyOufnZWFzCo7I9iFm+/PJCDA3tiaWV9VjBhJ44ufj3kZ+rYL9e4m/iXXktWbbqscceU1H17//LT6N7YCAWl1ejqaXN6xcA1g6y1gYx4sEi02DYtcXfrTL3icdp7kvOGH/FDc1tHu7OFs1E1BEcaxkEtK5GhFgZK2YxgOTmHON6yYOQr+rooPFgeUlqADwnzvMEFq0LMNIosBTfy7WxBgxiI/9cUx6hnKnGLN0eqQatIG2FxFR3d6dqIsrh6upicnpGz1MNL/JZ1kiRSEPyUxJsgIm6u1UUZuzYD2BVZT6SczDnZ+Yd+ffaM/7BHCD/XvuahzcqnAKLmZX5Y9kbXZfhepJV4rgmAYZildWoJVSuoeynXiFf/ZPXVgu2ysZMxp9ZZ6gdg9pPrM38Hef4R/l6yfs87v5dytPmPYkJWGF8O8f3HmyVAupz5J4oq7DPS7IZqfbiTatcscSXri+YDadzqICBzDo2+CfVNZgP8j+STB1MIRrClmeyb+aOje0V57mBaU+3FtVuiKNzP+Szs2mhulPJE5W7CRBlRrvqMwVMRp2KeJkYF7AS4wJ7Ak/eu3fH1PRmL2d+kn+zdy3MzetaAfocO3xE9TJYmZz37Ds0yVOe7WtGxb8w+b/+5z++EdjfTEJYKIMFbUvQB2VPSDbRVimyFVQxRrcySzI6HwSnGhtasCkdZB1tFzddbFRgJMQ6mr0Nki1Cg5gDmQ2I5GhXX48SKZJKocu6aR44ob91Z0xByPETJ1S4unbtmg4VDOOgR3IwsbkQ4HOY0YXlc2lAsOBJkPlc0BMkoiStHIQc3AQ0bBpcE8VrDtbdIyNKYKCGyvB020kliBV3eC0bQjLBZs/1UGAiUbty5UoJ1G3+SgBLkAwln8/mPSRFvI5Njo2Z//J+eXCA/tneEjoS5BNBZtKL2ZzZpNjYRkaGFVwRhPA9i/PWtuMAIPiu0gf97PTcShBYKf6q1Z2IeSPwFVTe54+QhmvVgyhnug6xUqzmEGUTt9m0dU2tv0xxokvXyoGDrAnvWyuFM5KOlGSS1ELFeIliN+gmF2aNZLcRaAbF3EeiPfIgkB5iMZRF556AiTnMOPIMeR7ZgMiGBvNgbn5O84B5p+KKWEU0p4y8Z/6hBS1PEhVcjWZgDktXtKBlk8VC4sFPFpN5ZhS3VZhGr7GMXS3ygNfXBjWJyM/fG5HlxoQfnZGu9pdIA08nlsgJiE1TpGFUMKwkhtW9KtG6NLZMvd+oGN0ToNLI4XdCpGdxVLT3bcl2ibJerinDFQKDlBviuakws4UkQpOKhKZx0qSBDbQsZEIaHHLtKbeT/hRuWlhKIMczC9WS6ioJtcwKi2wFBXh9bjGQIxBO9E9GgPIn2IE946DIfh5OlPlJKQmxTJBGoVgpWTf7GzDAjBEySELoQ8cvjRUCFTUqcn3UFnKLVqWKZJJ6MioepK0KssUs3nrRbhoasX6/LBbjKZPrOorqs4XF4Mkh82k1ZNyEYe1xrfydYI35SKJA4yV1NlNPmz1d3i8NNgkWbbW1OXq6uqumaaBFi28IRRE1SHdsuEcjRLJEKh6y/9jXRBR0eY9UmxMZ3CqBLs0I9iH2Q+1vi/ZJ4neez36d9goYaQW1aH8OigEOekFN0uTNBpSaVEVjP9dRrjX5V9SgmxhTZsDcvJkJVbSfUYx5zbkuK6upsCdAuPDdvDeTATO23Lwxk86N4jWkWVL2a3E5BocGdf7xnR5Tz33p9aog5oJqJhti10hKajPY7zjXCICTGadxLfRlnw0UY43mtT4vAAAgAElEQVTmVvOY5nBJfJTYFwaP/UyqxRjdcxnrbFxWGxNGfNUmO9l0T0BDPl8XgCz1VfuTiRHrqnYPrO6JeFq5EEXSwH8p0lGcoTCQbClJgdGkqTcal+IO5wVsUViVYlQ0NMbc7KxiA8aJRn9vR0fUr6/GnsH2OHZ4JFaXQPY1xfXRybgzvRgbNLdam6K7Z5c8KuqjMVbXl/z9W5uB7xF/Zm5yLYmSJb5A05x5bPTecsVkHZkvmotjd8fMXlhFRsnjw/Pcs2dEQI7rsDs5P2FYLi7GyZMnVLgdu33Hxb/1DbF4KEwBPJnA2JqCg4qoTpJI6nM/FbOilQL+rGTFapvhrM1Dhw7qPnytnXodc9bNwxXdC5JBfb3dGt+enm4h9ZO9ZJ8yfy9mw+yFsGLxHDCrp7qX5xwwk8oAEVPdjUbHo0JrszB/BJ4oDWkxaUuxlDmZ0oPMPWR0iKHYkz//7DPR6in2UZygMCsN/poJqMYtcUnR72YPVHF+c1MxwfGTJ+JXv/qV76lIjPDfLLrlPK8FEmThjLGgiaZ5XUyLGV8VSPR5Xg9iKNEk7Oo0im5rM9qbW+LVl1+O8198YSDGxrqa0W4G4LW1qmL/3MJixR8gzzcn3luxXRrlxL/yatrY1HlAo4LrhomBJBeFoqnpWd2jQCDyBnCzkrhVcVuRnMl4g/XjRtOKGm+sOfwpOJdbGGeaoIwhiMS1lRju64wXn308GhsoctHwB3DTFE2tbXHt0pVYXFyJ3j5iaeLxVbE68N6QFxGm3dPTMb+0Em0dndHY0hbvvPd+UApf24DRbZNkTLk311fjW998LS6eO6fi/1//9V/Fz376ltbok2dOq5lDfP/I8UdUrPzRj/5zfPtbr6mh+av3fx0vv/ScWMtv/fztOHPmUSE0WUOwg37xy/c1ZsiZKIbYwjS2MU4/dlJNfBrcFILZZ5hraui0tsl/iPhRUnqNZrUxpswzADycWfwk4jOL/5xt7GtI8ly9fk3Ffwp2NKHWVtajbhsj8oE4dfJkvPuLX8jHwwhc1seOEMQ/+Iu/iB/9+MdaW5wxACFu3ryte6QZaKAHXk4wyJkjjvn4vyz+iL1FIbrEPtqbiU1EW3XeoCYxcoJqxCXr0/PbjDDPF557bfE6ZWcMoDITmRhPBR+xHGzKzfpCpoy9wnGiwRDsaayF1fUVg38a6tWg43nIxwjPheKrxRrkuyvodRqdBSXsM9osETNOLdfm9cne5bzWABEDvrTvqxBlOWGdlSVWxkMDVQFYn8kWFdsvpbOK7wJ/F2AFA/PV1bg9Nuamg/xPzE6Dmd7ZDhp8qXgvWn6UeKG7t1fXzHvKFYhRxecRD1QlV7wvJ+Ke++N1sPZ9LgMSbNO98MP9ChyHb8b8rNZ3+khW4n18LNrbK9JPKRH2VYyKbDgxvopzSgMqC5UZR2RcwtgoT0mfvxIviTlX5l7m0gnYUkFzazNaW2g6DMfde/c0HwDr7D+wL+6O3a2cxblPM8agkomT9+zeo2ubnbobb377lRi9cTn6ejtlcK0YdGsnhnfvjcnJmbh08ZLitJE9I3H1+lWtORqaFy5c1no6cfJU3L03Fmub6zLeHRnZo0bFwACMipW4NzUdyyXnFMhtZ9tsNXmt2fcHJlObUOQU57ujr6cvLly+Eus722KU0TRlH93iz5tbbubjebFtGTXGg7lAHMG+wxnjpjRm7kgY469lPzhAnax1iqYAIjN2oznDXBZbX+BBs2pZ9wYUVQGOzCtiF6Hd1RRaUmzigjWKAvhwdgmAof2krk4+hsw9M2Oco2QBWOtVDC7We0RXd4fktCVxpqZukxiHxL/kNMyHWWRjS16Rc9UNuv+Hvff8svM8rnyrc26gG41GTgRAgFEiRSpRyQqW03js5fHc+9/N9zueO9Ee2xrNjEVFUqIoggkAiRy6ETrneNdv76pzXoAgr2et++FqFlumkbrPec/7Pk89Vbv23rWTeUVnLCwuR7dmA3p2mJWVj9YnlY9+WqOicvFPJLUNok7ze0rBIneRnN0g5UrmNY83KgT4u+hwfCmXp+rsZl7usjUVDO3eQaM8adcuj19zsyHRymGq8dAY5N16sRbnsdGk8NtL9a3Xy5+HXMVFcybUZzaB0LiF1lPOKDWmA15ogrCaFeP7dC6bGGonlk0axDs0iIeUn1q10cZPyF9k85p2z8LqIGJhnwyJT41B19q+7LL3W1HuY+tSN9XtEmJXDN6FnFINdbkHeEi3yHBFOlQDsObpUY90ax6k5r2lkkw5pBrnS7oeFFyoUdWwTdsvFCG8P2Qmzmx+HgUlMV7KXOysIMaNDIuYJ/VS98EvN+Puk9bk53/3+R34vboDx3thU+Lz6eTFw5hDBy0gFgcFCSMHcyVhGmyMJD6ZPgDA2nTpIaphyi1ehC1fhO0IlId9DHDVIwYSm42OPRv/6bOnFRywQYB9ePz4cbE97t69qyQDOTizCLiOK1eu6CCj6yrmf4fZNQASag4MDaXctTPwp4TlVBZMFNVT0/da6gYx+PoHFAhgGRKMTp06qeSO93XcZfjsqAIG8yZgb5L0njp1SoHk7t0p+T6TTHHP7D9s5iqvA9uR+4OSQ9L5jg7ZM6g4EDDRIZCBgEgThcSQpJOgZsZgCGgH6JMUGPkiQ0FpXGBf0t2tz2vPWgdyg3I+ROxt3BEbajrl/AZn5C25L6/bYpKXh2JZcZTBaQbnGkTJzSnbLbOE/H58LoJzse84iIrhouQ3G1edeRhwGLEmxDLUAL0EebOw5x4RvKW26QwlUH4fFy4cQvxabHaeA4AU95NfYVzyjA4eOijZLA0hkrS6VoBbd8u75Y3N4UOhR2LlIcNuxNGIwrKLoqOAWF339lbMzMyqOaYh4TBKKWrS/1XMeAZ2r7UHu3KvKwFqghvNpKiaA2K4NADv2l8CbAFLdOildLuGNSVIVfLyUn/4vRymlPtLYm82PqAJX9ybssdpz93YbakIBNKX93kxIVIFws8DqvYmU53X4bNTzlJYs7Z5lrBqDYhgjWXbOO4p18LfKSHZ9Z/LDsUgt69ZMQS1VWZuKnoDhdagGo6VYLD/iqXOXiFWVVHMtXEtZV9Rz6QsAkh6m40RtYgaw+X5N/17pjrcUNYQ79MCZvM517DaKswoDmnmAWiTrNfwdF2Dc9KG3YqHf/GfiufuHu0nvjzcy0kRn2N2ZsYNk8YAau4RMciMLRctt+7cSTDFns3cE+KKixc3o2uwphQlPQAZLhYFtqFE6scWzdYBgLBisGxtqdAuibhB/hoy63XnhqqTdNZgJetah2khs0eJ3boAWcB5W5K0bbis9nJKZt9lgwYqMjJGkrjxfaXAE+CpQbre36UYxOIAIFHNst2dmNi/X68naTgzVtKqoslEaib61bwQiN7TK3C3VG5urvlz1ZotZpvmeGDdl7EHFiigo+wxAIqSQQ/wDkCphkaBpBpObiDBKpjtmNg3IaC1mJ8aIpqS5Tbbx+CLLXvaShWukzOrAFsXkx7sVzIssZiSuV7WFmYU+zr4qsbk4wzzAnibDalmsvR4o6IaGm6qe49RrHNfmD3A18OHD3Qml783/+ZZKajAtgXCw5qUYi7BVFiTek0xBD1slbjdw4dY34z9ezvjpS+cje11ZrOsxOUr0/FweSM2OJeQotN0X9+NudnFGB4dVIObnACbJzyPPYPAFkI1j4o9jmKAOA34CmDMM6I4Gej3IGIVRlhkYoWy44YxKlNWNHYxxE8Y2AD3AIvcdGZeSTXAfC4Y1WNjAgTYw6xvYo5thdZV6AGooviRMnAJOXqfrDCxDZEvcO6Vs2fPxK2bt8WEPH/uaeVb3DP+fmUF60yDPvz5w4uX49jRg7F376j2KI2DGhgPoKhaurszbt2+Y6UXLPJsZJRyFbYphVYNCCYfYywo1Aq+1JRML3YNmpQK0lZZno1AzpnDfrMBR25WcwK4ds6BaiAJRKUpsI2POw0b9nl3i1EM89rMPTf1iLVnzpyJN958Q3lfreGy8nNjySrfWsdSmDQUY5rPtWV1QimiiEMsbDXedndidX1d14OSZO+e4bg/fS86dzvj6IHJeOWLL8UvfvYzFdeAT1ieyF97czOGR/co5ksx0m0Vl5qZApJhOG/H+upq/Nm/+NN4663fKj5/4xvfjB/96Ed6VrPzc7Fnz5iAJ1h7stlIr3IaTbXvq4HBfeQ9SoHGmY7dEXkY8Wx5FfIBZ74tE7bX12O4tzvGBvticnQovvDC07G7xVyEndg7Pqbh2cyY+PjjK7G0tBIHDh6WrzuM7v7+ITW+Ffd2d+Lm7duxZ2w8rl67EcdPnY6llY24+PE1zUAxEzLiwOSELKSOH5mM5599Nl5//SdiJrImfvvbt0WO+Ot//dfx9//w32J+bjb++q//Kv7zf/47rbV/9Vd/GX/3X/9OceOb3/qGzqA333xLVk3f/OY34sMPL8XVGzeifwCrkp0Y2bNHYOgWqqxRD6hFgVPEgyJwkRNyP9jjNMuw78J+hC+USny9/PJLIjBNTd9vkRMsHMQObSi+9PIX4tdv/TbmlwAUUaj3xNrqevR1dcbJY8fj2eeejf/0t38nX3rldzshuxPizl/8xV/Ej3/832Nq+kGMj+9RM/LBg5m4detO9A+Qb9MkpXawakupTtpXtsDkUrdSc+V8EsWrrDfK1s22hJ63A4DoGtJWP9i5VW2gQaL599W0qP3DmpNiA1CKRrQY3wCtW2JnC4Ci3lpbs4I51Uqcd6jcAEGtRHHjR4r0JOP4rPMgVjXGia3EFcgd2cjWTInGnub6TDbwe9WeqBqn/t6AuT9rNd3ZA3iPi4kOWzwVFwLfsL7d3LCiFpUWRBkpQD2IFQUL7H55ls8viEX7wovPx+s/ed0khjydmYlGjXr/3r3GvS/Lptno6LAds2yF1Ewin7NSDfVz2esRszSQe2XV59XKioBx1sDi8mKSimxfUveDz2lrNjPzlbtkbVm5UbMpVfeIv2vmCZXLuzZpg6qQjGTfwjwdqXf9b2rAp0rAM+zM5hbYPoitkAlT5L7kguR3zFp7+uxZ4Qr8mfpfDeMtA9UoKnimnuW2GYsz9+MH3/5qTE/djIl9ozF5YDLu35uOu3em4uSJp+LM2ae1f69evyrLu8uXLyuOPvPM8/HR5atSop47fz6mpqfUYGY2w9FjJ+LDDy7HxMSBWFhcjfcvXdaeVjNGM54gCG3oe2lM9fZQ92yrgQA5ADUzpIbrt27FDvdwy3dEdQvNxg3WsWsjFBXkvLI4k8Wh95Tmf66utqwowQiaDgy4GIjslXMrClhtOQ9s07QwFsSXbRvtQ4iarAg55MJD/VYTqubLofEo4PbuG5fCr8hFNCH6ers0j0mzn1KJQx6CWwazk5jdAhAu4iJ5fG4A6idwH/YZZxH3gjNxHhVUkpsg4PZiC7W1E3tGR6U6W9GwZWwKfe+tBG/PFGw3MNsWw5X7N9doM5et3zcbG482KtouAa59UpGfTap2o6LdlciQnPmFldLV4FHMzCrUgD2GX5/8ajYgao8192fVv83rd76fcabsF8p+KutUf39dQf0pf9WsLaviKndyLDD+QKyoP6uJoXmqYA2WgtNYFLmiMQOMBh65BvUN64AcWKQRzSp0I5z1WHW9bJp0VtqhhXXBuQzxZ/redOxNfI4cnTKGNcp1oSjiTGDPeOYbxBITyNxoJ87b+cO1qxuqsrtu/ErsAYdivYrAlbNIuH6uhf0OyePChQsxODwo+072BValcuBI9T+ve/wYllCdqhl4XWw7aXbw8+QsnzcqnrQTP/+73+s7cKjTIKv8HiWBpbsJw4mDkYLZDGWFIbcQs9NoX0GOR9jRYpqkl3RlTirmYCs3LGhQVKi4o6BTUoyvsGc0PHP+rIINjHvYRQzO5j04XJeWVzwkOz2xGY4L4EBCLaC2gwRpTck2BSkFKu/DjAsAQRoVBGHsGDxscrY16wAQiEBF0IJlweGMNBOv2xZLPQ86gEsG4n344UUVeHjCMneBQoWDlPsAeMD3AUxJQTEwKCZi264Dr+C+uHP7djYZYH8yYHyffp7PCwOKhJEkkdfDdopCmtciYO+b2JcSTQ+G8rBbD/1RsZxMJ55FscRhScHEsoza9kAtMCiHGqnx0PBWLXCpBjUVkNEEFjVQOJsPfTnEkWAMw5N7zUFjZoY/ZzuRt8ctxV6BciqwYX2oY04h4aZXMZvckfb7FaOa5J5EXmCBktYdBXhAG5IxXgepPy+EGgYmGYec2Naac9FtMBT1hlgNJPE0J9YTQPTvKbbo3hfYzTWQ6Orv1vHiXPCwcA1VbA8h13PBkzvZWDr0BU70Cjxg/VUyoH+rBD2bMK2kvZKERsTxa3lAerEX9P16zm3JZTFN6yVsadbV8ulWYkTimcmsPLQp7CRddNLmGJAFcBZqlHje73kd+UcpQfJnGPLHoDUGnmJvAJuQ+222oBkWpaAgkSkbH7G/xZQGELfNB8kvSpUCUpyUWI0gFnUO1PYwZxeTrB2ShAJTzRrzZymGfTHUBX7rM1gFVvdeSUnJVDUsznNNSHz4Xpo8PFPPeLANBM9FIHKybkuOKok5iRWFb19fzM3MmPWT/rEkWLwfr8s65c+wwWtYLD9fAJkZHrAgbbHF97I+6/PzuSsREsNaNgQGJT1k2NYrjhMU1hQfnqliH2MD2YB6ng3gwoW10y2mIMPBvG+I4SrslpfUVG2nrWkhV3NUxGaxpV7zzKhYJMu2LWyMJlW8I9c3y8Y/I/k3+0nP3gUSDR9ZTmTTiM9iH+rZdhNd4LXVUaXokL9zMl+4L+wT9jKqH94TiwwUeKyhioWVzNuuzAoRDRGmsclQQYrJsTGxXgzS2N5LzDPFM8ugWWjEIjXKUia8sbouZR8gdp09NONlpyBbG1HWWmtUoG36VbMuzHyEGWdWkJRf2dAx4N+2nhFohMVdzkkqNqfvodUy1aDITZ50qUYAav02zdQbcaJZ4DVjx+NFXvPf+L2aoJ/4YtZLZ4wMm9WN4lFrDGug4RENC+XvuccqCtTkZ58uC6RgPwBO0vzinkihwlpWo3JHBfQwzYwtGhXd8bUvv6hGxe3bD+Pew5W4eX8uNvEkHx2O4ZE9MTuzEHNzC4pVFNHMl0K9SfHAmU0jG6AHUIP9wlpgrVV8pSHIdUJOgGkFaYG4wz6n2BAIphkX456nse1GOg0RzXzRWnVzjvVG0wCwhZhC/kTjTWojyecNwoippUawlSnkJqwfQGCY9GrGp3qQQaB37t7VtdCMuHnzls7hY8ePKU/ENoa1v2cvPsBzshUaHjFxAssnN7oNYnj9RUwlCwywwMCicxM34A0CcM6S4w2o8bIpwJ7GjJpgCWpZeeLB14ApNIpoYPEcxMzL5rHYdNk45vOyXsgrKg7SBClVU+0LxW5UBOQX7FVAhO0dFYOnz5yJn/3s5+nZ3Z4j4v1vgK7AOa3xzKO8vt1E5rV5No63VorK9kGxkMaGUgfFB2LQ/en7wUkwPjISX3ju+Xjnd29L2QbA8sxzz6j5Q/60rrjrM3Xv3jHlzxsbO3Ho4ITyc/Linu6OOPf00/HxlesCvgFqdC32ZtC5ak/xJTUIYOMSAgrULcsFctna255BUIpc+9tzPyAa0bjmM42ODMcm+RUqkK2NGO3rjn/1l38csUNuCGi0Fben7sXxs0/Hmz/7RXT39MXw8J44cPCg2K5qopNDrq7qLGBG2+Shg/Hbty/EwNBIfPW1b8Ybv3k73vvgcouwcuLE8RgZGoj3L1yIl7/4hRgZGYof//h/xrlzZ2Xd+o8/+qd49vzpOH7iePzjj/5n/Mmf/ECx/8033hSZBb/nd9+9oGbdn//Lf6EGyuuv/zL+4i//VDnf7PxCjOwd0++x24JRCYN5aLBftrDUIAbXAKKxrKXh2xHf/953NQ/i5q27nvm3BUCee6GzI/7oj34Y71y4ICIUS76n1/au6+ubauS9+OIL8fY7F2KFtS6ApEszCACaJ8b2qfmA4oL5JTwvYgPDyv18B+LSpUtx6/ZdsZ8PHTwQR48eizt37mh+jHMnW2U6/1DfosUA5dkSb6RM5dyR7cuQci8DllYE8fwVfzUw3goy2+l6LpeIHtV8INeXWtX2VLwWz1lN8pzH5cHajltZgmpdal+1/r8BxmKSdvd2K1ZWXslz0jXshHK29gwyE7W2t9s5VakmisntnNANyGrMEUeLwCACUsP2oywXyQfctEbNijPAou6FZvPllRa4LoVHAnciqAg4ddOabBUWP7/XMG9yLhS3OYSaZ8AX94T3kwpcue+uGg5WpZIPZF4nG0WAtR1ZPDpUPcqARjkL2agIGtw74sDC0kJL2VRNhmpAENv47JVLk4c2wdk65wssrQZP5bAVUwwUm9hStSJrrnJ54rfmYuVwW545MVC5rUKZQVxZR9Nk2bPHZ2TWHGysY0ePaYgt+3RiYr/WfpFHyAt4L85mnv39u3fij7/3WkxP3Yqhod44euSQmkHYt42O7o3Dh48ox+gf6o9703e1n4hnr77ylbh0+WPNa3rhxRetqNik8doXhw4fjYsfMqdmfyyvbMaFDz6IRQ2nJlfMAea9kDp3lQfTNt7axO7Q56UsvdY24gYYwsZmdON+gdKAxgx2hasmnHhqpP8DS2Gdku+yToipVd8I9K9cMc/PsnJ0vVSNTxPH6llWHm0lm50UWNp+BDSNQkqPkYE+5Qis/8Ie5haWpK5S/oVqLkmOOo4AeQf6ZHsJYZa1wbNcWF4RAM/+45mqOb/Zxjx6NDem37Z5CRoTK8lVyMeIqcp3O4lVJiahZOH8JUZbjeC8t5mnVs1Y++TxP1e62mwE1H16Uu5bgar2nvOBR23WXWon8fNJKXc286Q2y/pRTeZsVFQTs/mjFcfquTf/rfl5pSQVOG/y4ye+WrKxjLtS/VvxTx3Oun2EwCoHhrYzR/MlDXm0LaJMXEMRx5mF7WG/8iHsVWl4sDfBJqoGpnlbOT5PkDqZGGS7p3IhIDauSfVohb7rf/aBZmckyVoEW5p96RBhVZ+bfKwbznPsTmWTmPhMvYdzZzenizRalr5SrssS1QQP5Zhp+WS75I04ffq0GhV879FjRzwDo6dXTYiVJc+UoR4+ecJqZxHKIDmsrkhhhx0s9cfnjYpP2Syf//Xv7x043NWbTAN3lUu6SwHoosOJa9sbz7YsbGwKRTalGW1mJhdDtRoeslVBUZGSLVgdJLhSDyRrhAOHw3N4eFBJMAW8CvEEUAg4bEYNo5HvdoeSgSpeBPj19Kqopsiq6+Za8FoGnNZ1AgAmK+bGrZtmLuawP5IB+4abLYdaAesnghpBdyfcwOG1sWsgsAjYldddt4Zzk8zRFLl46VLa4SSzo39AKgoSSxoKXA9Jw82bNwVsWorG8Ngx/T2NDz7zgclJMQMADLhHFA9YE3F9JF00VzjEC6Thnq+vApSaocyJVSx6zc+AQZOAQB1U9bwMkNvGSMBqypoLbG0ll6WcSWBYCXIOBnJPn24yAzztWcrrVte/ClpAOH4PM1PPWMU6t9mspgLVlXimTUI1FOTPmxYKGuKXw2pJTmRVtrMj8I9rQI7N82ZdAICosYaHJmtsYVHrlcRJINXIcKvwoP8Pc4/nS3FhDN6sWxoRVbDxWmqsLfp7AKckrVWDJUFYgTCe2aIELg8pkjJ+r4HKyVipwc3VfGglPY1h0U9KGFpNjrJgaqlgSNydtLcTI3tAlkUYr1dSacDusiCqg9DNL8tyK22qYlCej15Ircsqr8pqVPArn0+J8CZr3bZs7BmaSbZScrJKXIARxuvxXObwz057AFno5IBrWQPkoGvWjoYrJ5CrBEkKDCuKOPR5JiqKshB34Yk9S5v15X8v9mn750l4SIJ4PxJlyexllWT2Pp+PpKkF4ONlmYChhlFmMgljAjCaBhBNG8mv06qLZElDbzP5oOEptkwyxNq9INswVCOxAF3iB2BFMRBJGHUNOWzRhYMZv2XHZwWGn6mGh8nux6wXew473XUhbcCTZF9gd3qDssYp+lXgZVNGs4QYnokKrNXDcqNCzZ9k4VUxW8oKqyjsI1r2XjRuafhWYmlbIhfDXAeAJs9RBWtakmjeRAJnxMdia9U6V5HEnIqceVOWS26q+4J5ljQLuL/M2pA1XQ7aLbC/CpXm5zHwj9VAr8BC2P4+Uz3Q2mBkewerwJc6h8LUdhfMqJC9juYRGLAvYLqG0QkAbcxtqSYu10Jjlusmxtb1uDHlYq72RO0R20PZVsssLoO3u8wt0P2oYaDe57Zf+GS+UwzHZlFT19gsbP85mVKzwGt/v990eJDZIQZ1WeOyCejp0TkpMFYgBvMYsGVa9wyJdTcG+YyLi1g/mOErVtP2Vqwsr0UfBRE+yV0dceTAcDzz9LFY1yyr5bh5Zzam5lZiHRn64ICAjbmZpVhYwMqpWyxfzagYGPB15FA/CmPAMhQesDQ5uwDwiAFlw0DOgGUL+UOtPeKJlBW7uzE2NuoBfLI8hGW5LjQGtjD7FbsO/n5lcVk5C/kHzSr+nuIFr2jYubyGFIR1lhBjl1daSjZiUz1Y4hrqUOIHoBfWMDS+uNesB3KW/gHbbXH/YPh7TSbYtUNMNJuVzyAW9PaO5PkVc2neFanCzQxsXWj0Mdy+OzqjU68ByCCWPgBYNgt1/goYwfoLgAXmm1WnNRuNe/HySy+pMcW6/vDDD+MqljmbZpqqYZM2AKx5W8KYHafZE+n/XGxHrIFQVPzs5794QqPCjfYnNyp8ata5r9ls2RAi/LpR7DyRJr5tFD0TjOYryMo6/uN5dp1gKOzSYswuLsXT509riOvqOiDsQDx8OK+mDteMaofPSKMLr3J93p1tNSfm55esEB4etUIX+460AISNTkG/sLDk+4FVZdrlcI3k+uTu7LGa1UUs5x6XHScx1qz2agiux8GJ8S+KfaUAACAASURBVJi5eyd219fjxXMn4yuvvBgdO+Tj29HbPxhrW8xjm9XZynufOXsu3rnwruIozSUUCuT8PJvB4SE9p22h6D0xMLQnLl25Fh9cvBxr6zAW+2J87944f+6sZmP87rdvxcsvf1Fr+O3fvR8/+P6346OPLsf163fVoLh166bmyp05c1ZEJpQVzz77dJw7dy7+43/6+zhwYCJe+/pX1Og4ceJITExOxk9/9stYXl0VMxdii/tLnfHqKy9JyYF610OoHU+ZUcE5+o1vvBbvvfe+1B8iBSV4A7hCjvDSS1+MGzduKn6T27PG2d8Gijtk/aQcYnhIYRgbE6xvO4U5O+dBBT4ytscWstiSJhB36PCheOedd5TDMv8A9uix48djcv9+1ROeWwDZo0MNCpEIEtBhFZdSDsWUFJViM7t5UU16gcZYR+WZzLnHdZRPN9dOHUL9ZAVkWtOlkkC5bKot65gpqxPew2cmzfrMR3P+U4Hl+vmOXdmiYRdCPK7ZU5rRtEtTouwN27ax7HfimBrEqbIwWcM1nkhQqa6oc5JnYtYtOSbz9dxAoC4G0OIzk+tyJtm2xMomvoihxLCyIVFTB+Uxsx9RVTGDpNf5FaAtr0EjvBjB7C32G+eImoKafWQlD4ocW7ptaj2rwbe46A5oEnRYkygLjA23AUTFoc4u5eHk58pBdndjdHSPFB5LK7bSqVpAeX4+Q66fzyPbnVT6Vv5b79t+fz/LykMqn6o8y03s9vVyTxWnAeUhOjZIU+SIxFeei8g21agewL5qLWdS7dV9IK8iR0RhzT3hPtEQpnEjEB0F5uKSCIFgAlixbK4uxw++87W4dfNKjI+NxKHDBzWEm/8GB4eFSwCWnnn6qZjYP64z7MK7H8RTT52NCxfeE1h/So3/OwId909O6P5ev3Y7Dh44Enfu3o9bKDGZBQSJJpXRqBF5Ntgpc28BbVHXUB8wo6S7q1cYxfLaanSIKNOpxj0EIhJN7olwCqy3Nd9iUPGcz0+DhnXNs6w8kfhBHd0CqHPQuhQ+cmlIK++sG6x+Bxju0R6XagGr2iQh2MTBJDrb9HbGXgaXp721lPpbW2o8y3o2lbpy2tjizyH1A8+efaEcPUIzZgrMpgGHegPmu89sq6upF8EJwIg0uyrId7CesjMCuQR4wCqKzHXIPGBaJttUo6LWbrMRX42K+req0Zs5bq3rx3PdRwB/5WE530g4jYkP/vL8Gu+zHOj9hJzb+Y7vW+Xsmt8iFN7ZXLMx8Vm59+MNDCuuawbio42K+hyuJZv1gWOJPsGu76N7LamoSEJE61M2Pm81ZapZ6XmvXltYLu7fP6Efs5sAMQbVlpvm7FuUiazrzSQmFmFENVXW+UWwUyxPwt3AkOfY8L6a6dbRaWWhGh59It3YKs05ju+JcZKCVWT5jS00BEasUrFi7uzUOmXt6zV13lmxVecI+aIb/NjmDQkjRIVPM5jPzl7k9SAvoRTi51BinjpxQt+n+WLdXVKkmry7a/LW59ZPn7XUP/+338c7sHedTbil8NKUqXMIOQg7WbAnsIEygxswbTyPoNWUSO9eJykAH1i3WObLZhQoBT9sN+QZuYa/oMBeb/CTJ46LhX/jJon+dJx66oTY1xz8d6amlAiePv2UvHhhBonxLYaBr72S47J+4hopFuTpubysJgGDlSnmKHrKn1EBrKcnjh87rr/nEKdIgQUJgwsgm1YFSaGaCfJ2hLmyYrun7R01HSiK+R4CComr/FVVYMO6H1ZgxfoJMIn/7txBegoj1x1Wkid+vXjpsthOMEHwyyS4UXjDgqrh2zyLg4cO6L1JuLjHJEvyvE02JoVTHUDyt+d/OcDIB62ZfARcNxsMNKgZkkOKCmAHYNH37ZqhrkNiEFa4bVUky0uPaBJ4vvg77hdF1x6Glz58KNkyQZbkks9ln2irD1oKD0C7ZKSX9NONgj7Z+gDukaQXq4nv5fmJxba2pmfN/eW5UrSikiEZxZ8cNczsDGoagGLL+3gdEr8CsklySCjLisrJghk+Yh2i6lDTyswOEg5sGDTPJUEy7k+BsGpwydPTg+dIhqvY4T7xzAUk1mDq9HZUwyaZmUqQPiXAKHEotnraA8kqJQcQ8mNVUHDAtgpEyS4B95L5yh7aNOhbg6TL2z7zDceCUhzUgN/GdZl7Y5/iajgV0wrWWk+PfYaxXwOAJnFmH/J37HVAKYYQ8wwFk2JvoKQcsA0/STxaSRQ8JNaFpRuITiRcOGpN0FyQhY6VObKDScWRbGs088KDCosdxkchMRYYVgOUE8Tm7zR8MeXQvLeUU1h/kfj0WfUh+Woq0grEMXPDrYHysa/7wmfVYPf0ApbUVOx/Yo5lorVOlCBlUwCgQIUHKqDNHAbZ2ZW2U04gK2bzeVXkqZBmADA2JX7+9gp1siVQNGdWSEHBvdTAcT8LyWUHB+PA/smYujtt28AcOpmGVbpuCmlsFrxHeEYWLpPk8TzVdEiP6IpRpewwULAT+ycm1FxW4zqZ0gb0yqbGTbjaJ2YNGxxiTTCvATVagaB+ni4E1ZxLtnQxkmRzxbDr7W39LOuLmFu2WjyvYqUb8PfgRymjUmbM88ZPmviDRVwN6q7CqhpoxIb6PezmUmtsrhn01npJAJO1IZYnMRUFR64jN1Y8nNtN2m0xKPmz5vHk9aoQzaKj1D0FxlRzrK6lVByeB/JJn95Py3Eeby5UMfOkpsNn/ZvjzBMYXJwSykc4U7tVcJblnRqYXZ2xd2yv9te96Xst9VQ/Njo8UwAlchKdyShNPLTaQMmO2H6Lc/Mx1NMZxw+OxOmTk7EpILIzbtyejTsPF2Mb67OeLjUWVlc3NaMiOj2Di/upphSS8wTmWOfOlXaVe0hlkM1KKyfX49ChA1Jj4pfPXl9d5lnDZDcog1IDsPX21F1dqwaIb27EyRMn9T0MAaYxMfNgRqQMyB6aKSTbki19L4A3YFbdP0MGbp7LbkTFrWNhDSI/MLlfeRLNFnIP5nkQe2nWU3bSwCMHOnLkYFy/cSsOTO6LvXs89Jrnwhrk81FksW4BdbFGlIpu2zkkv7opmUzMzBk4s4mpNPhoNpWKhJjFXpZdV/rgY9Hk/e4cRjmEbN8G4/nnnlMOhcIEIJprJi+rfKcXO8KcqcNa0LpgVo0PzLQj8KBLAMCnTp+OX/zily2VWTXiak99wsIkFRUi+3DXUt2iBn+qWwpgrRxEzQrFT2J1T4yg1lxeiS6pYOxPzt9vxY6aCw9nUM9ghXYg5ubm3UjaSHvFbE6o+aJ8tEv5EENyu2HubkL06HFOKHLOSGztMMuLPIrGWKfstlBBV65VFnUVB7gHtfZZ39i1AoQLvN3cjOXVpYCcP8RspOXFGB/qiz/+/ndic3UhBnrJp3qio7sn7kw/kEJpZHSPGoCcs1wDbFypYjSjwumQFJLk/oAI27vR0d0flz6+Fu99cDHWNzyMfZg8MXbjW998Ld698K78rH/4w+/Hf/kvfy+g8Llnz8d7738YK8uL8ZWvfjUe3L8fb7zx2/j+D74TH13+OD76+Fp8/3vf0dynN371VvzZn31faxfLM4ZR//Rnv4qVddSUgPqukzq3duNLr7wU165ei6mp+9HXZ/9rs1NtNUKza2FxQQ1rgJBS/JA7cN+pJ6g3+BkaFW7CMT8pBKACfAN4Moib14FcQuNga30rDuyfkNLs1799K7Z28ANniKyHYdO0R63xN3/z72Sfy/1DJUUT6tTJE7KNoFZaXV7zUN1sQgr0TRKAVA85SFse8pubAkKL4NRS3jaIK2V3aZvUZHg3ACp+2OvHZIACoZtgdBHotNakAiaH6W9ZEpfVmfM5z2uCuc58KWoPzcvYTNAtrw1gkocgYDzPFH6+2P2qbzPXKGCp2QzR7JZgcPZi5mBmNbPmS4FRhAriNuuPzyrCVeb7/Eq9q4aHAHjnbtQ2NCTWNtfk8Y9Sp2b1EUdYB8OjVqtzzZ47hpp1XaAeX5w3N27eVp7NeqJxaVDaKlAIJbDzVcto0K3VC84XQ2cKP8fCA2ADSDPzfVU1d80hrNyxCBtWVLiBTcwwptD+KmC37m8zDtYzr9yjGhVFtOFnAOoFsCdRQ02xtIWs/FrEss4OxQGth85O1ezU3qzXvWnhTI1Hzkg+7pkIbmChwuVacGOgWbOzuRp/+offid/97jcxMjIQp06dkNIWlwZmTbAHmR3S09sZTz99xoS2gSHFM2ZU3Lv3IF798pfjytUrsb6xqllOA4PDMT31MCb2H4ypu/c1SJuMRNZN1GGoYpeWVaPKfjMbWW6ye5D9+tqm4tNOJ6oFnp0KeZJbWyvuRGygFILQ0+G6hv9Yx+SUtpdqz8dTLSu1Aoz1XtWrdhKwhbNqZWoEhg6rbrNaiDOKf6MuwHdqdRn2d9oQJ84gsmvaKnV0dseekSGRNtgv4AH82+aGSa3VtCpVkGr/Xs6uAV1H/+CAzjC6EsuLy7pX3J8Cp91MyNqujwbPkCy0hA9pAP2WsJKh4RHlJZyXZEQtq6TEImq/V05ar9/MX6uObzYqam02c9lP5MGpIhDOkbhK1dUF/peyyPmN9emtNZ41QHKJsuYuZcknGxVPuqbmvnz8+qp2eHzvNv9cNbQ+ZzYs9Iz1TW176RZwocvytfmrnefX+3tea6mqd2JweCAG+5k/4j1fmBr7lngJSbea11o3qf4pwpIwKs0xysHbslMbUA4pZwOUxLITtE0mX+ThxHc5G3SkrTb7MM8LY2KOk8RPcmasm4nbrDHqeT4ncZnYCvGDpqfiVzaWuFZwF64LQhvYIc4c1G3Eh7k5YlCP4nip9NkvxPORoWERkfh7NUi6OmJ9azMmJyZ0Tz5vVDxy5Hz+h/8d7kDf/KIPInWUkSzVYL9kUyYL3HElZWjJBLXthL3bCnRqsas1r4ADl+PXTQolpFikhCVXg33Mk4DZaAYusmz+zIA7ZJmHjxxREkdC9vGVq9qkJ06eUvKJZzOvBzhBkiYAI9kCJJuARCR7JOCwDK9evaYklMKfoGSrJBfMHLx8tAOTB+PatWtK6I4cPqyCgO/V4MkhD80mCaZYwN+SQMIwcZJMEiIKe35Pc8NgsL3+CcIA9tX0sYXLtliWBRbWAHDeA+blntE9ln719grEwN6AZ1ReoXRbScTEyOns9LDwmVl9Tw2hk+Q8B+KZu2UQqHUA54D0AifV4c335JopPKqRAkCvhDubErpvsKST+V2MXVhJ1VQo2ysPAd5Vh5hg/vDBw5iZnReo4kF5+Aoip7M6pZpOFCW9mkFgWxosJgjgJJ3qiotdgpTaXoSaA5IsZBJt7t3y8pLWAfdfgyV33XWmGQPLCSBSPqu5FlSUMKNhdVWNMD4XF1AzOTwU2OAWP8fhQsEnoEescR/UDOaiOOT6tKcSNKxOPNdSyXo1KcT8aDQrlBA1GhWfFm+UHCQ7qZI8rrEsXarRUolTqYhcmG3mAM4teWGzbuurErMaclV/X1JNXDCV3NXQrATAnHjZw9gHstfx9jZNOQAhP2ueg1mdFNQMTUWq7UKZBIBCnsO5Eh3J4RNgL+mmWUcGLyhwiAFqmOXMAlvoeA5ArT+eEffAyZEZP2UBo4QOwCx9I0tRVHJWgQOAY2EWrlUyFBjed7yu4mGqP7iHrOny0Ac4k1UCbI2eHrF8SHJoUvIZ1LShmO3Jlg/FL/sSuxPYxhQgqkes0KnnDQvJvvSwDT1EWHJTAVLZqEFttJrsWnxkc/ZC83njJytlRvpxah0BJqbrqYuVLQOdYj2l+oJCQwxq33spXpKpUgMr3WwA3HcDm73dVmzxDPPsScb0gQMH9ZlhRVqR4TPFjW9Y2G7EeEh7b2sQcd1zPMUpTmvgtlmdJLNm++j8ylkrakYkiMGeGN83rvtOgV+4SyXvVZSbEW7lIddDk431RpEHYCAQQ00V32HeS+cJjbFku/lMbagd1t3crXODNaIB67JWtBUjVy8FkRQ4vv818JsmB+8DaOlBum0FZDU+3IwwANv+LO3B59q/O7U/fGa4+HvyEGyHgE9ro/6vZ0mf1qioeATLCvsLWVai/My3NuMfkIYmjRtSGyTyWTSJodXbpyKfhoXmN3D2h+dD3Z+aju7d7TgyORAvnDsRm7KSjLhxZybuzqzEbm9XbHd1xMT+ydjejOjt6ov1TQAg3yM/X8chM9iZ89Uv0Bw1AWc4+wIAn8Y5Z/ZTTz0loOPevWk9w+1NXoMijOe+GkcOH9Q5f/fuHVnMCAja3orTZ57S2Xzrxi2xb7cAXAb6k3G9Grfu0NgIFXrLND+Qw28YhOc+YKmg/KxApZynIOvDrW3ZPTHgm3V04tjRwGqT8/7I0aPap8wxmJ+fi5Mnj8fNWzflzc/9L9a195bnZzFrAFAcZaj3jLea7dJysGZuEj47IKobFR2xUw0UlFIp1ddQw7V15ULsHrFDe3qip88exMTqYonCMsYy05ZxnvelJnpnRxw8eEh2jRSS7WapB5lq7llK+/k3GhXMN/jlr97QWVLrvfYP91W5VmPml14z82czJE1cEbArS1XbohZTD7ursjNRmILZjHoA0sjaWoxJLbWl5s0aM7XWN2N5aS0G+1EWDYqZCgAp8DjC3s6axYONFbk3lh+2Y2GtAdBMjI+J+cdgaCwNaBCUfSALhXVILqMmfc6H4XOJ2NLwqOe5i5GMfSasQWbj4B09PBAD/T0xe+9h/NH3vhHHDozH1PUrcfL4wejc3YrxA/t0j2Zml+LDi5ekAOoTGYSGjAlEgPoijgCQKVen8bIRvcyFwMqjbyh+/dt349qNO8plWOs00lEmnDh6MM6cOhWv//Qn8dWvfkX1xFu/eUsN3S++9MX40Y/+h+qK73732/F//dv/O86eORNf+9pX4t/8m38TJ06ejK9++SvxzoV3NKPl1VdfiaPHjsX7H34Y7733ge4fJBuxdpkBNTwShw8dFBnCVhFduh5yZ541+521Si3B5+TnHzx8qLXEuYyS+vy583Hx4kXZyihO16BVLDOHRuPsmVPxzrsfiCDBGqGJCUmhKzrlXf3sM8/Ej//H/5AKhfPReY5B27/8y7+I//Af/qMGhB4/cUzn381btwXoDw9BwNgKNpwUqqmSltI1azevedtDsZ7IAQQStywurdTl+4qwxV7hC3KEgKEcYl97tPYd+6LuGa9XKmOROXKoezX9aZDwPmqc5Pwr7h8KMXJJGjTkQZolcP+BGbhq3o0afIWIISsu5ymafaJZDSYaOddoq5+LNMD692f1+uducA+LIe4fck5We0PKRqxD+rHLzIHidd0Ne02GAGM9jPqb3IP7srGJ/WrNDjHRpFXjwvrt7FBDgWY013z//j3VteTRJ0+elBqAWpq4Nzvn5lj7bPWZ3m7w+lxAJasal+b2AkpxP29ZSjLgeQkWrwfL8qV6LW1jy5KX4E4O5TyjKiLnAc1GRWUGRTAsQFwq2azjCvhUnqs6jJzWilqegxpLzSaLuhS2g+YZDw4NaP+RU01PTYkctXfPqNjLEAV5PeY9aXZgsqQ5M1i3k/snFdNWVxbjT//wW/HOO2/pGT7zzNNqKk5P34vhIZRL5OWQcnZidM+w6vqvfvVril3zC8vx+j/9NJ5/4cX46OPLmmExsmckhodH49rVWzGxbzIePJiLNRppnCHMppKFKrWA5+wxa8O+9uQrXTrjRodHlRdi/UczGaIccZT1AXeCGrpqeBRM5Az7xsZUc5HT8jn43IsLVs2QO6geAa/QXKteKXloUvFcuDfsG74XMhDnB/uC5wLbW5jF8IjiCNfHmSIr1pyPiUKCn6NpgpMC93dkyPOMypFjeQlFi2s8gfSqs1GDeKX0dLEOhwX6EkdZIzx/8iQeusgnmmHn/VuKYDYqORifg2YKecXcwrzOSizFZRdtv0VdL+u/1OPViKjzrpqXT8p3K5Y1mwK1xj/x/S0Vhck3hXGIaNpwULDltgkdLSS9uhUiEKcfnj5vxh/2RuM1mnuurrGZldf1NvPuykk+q8HRrAtsXZcNz1QRtt63SbJ8hIPU/kORTKrOs8oLpYExQnIKZsiSr1ITku/gIsDaITbJyULEPezFrU5nj9Zn0hpOu13lnonlcX+lUk7rY15P80/TOYAYonxIVqpWJld+X1gaalvOWc59Yjixkz8TR3gfag5IzbiiULNwrSLpQh7B3n111bPs+nrj4sUPhZGNj+/VHiQuQfDlPSFusL/Pnzun9am5YLNzcXvqTkDIOjg5KZL3542K//Wa8/Of+P/5HRiFtdRICgpQk0VGBskKgNU1dYJWLPgsWrK4K5mg7Vlg1mE3YlsJgQrRKQmrDiQx4yzXZ7jkvvG9SqhJOAv4BcDTLIFuWxNw4LLxkUAJFNS1u6BCbcAhabYLYOOGbDTwgEbarICfSSgesFVc8isKD5IBzx9gUI+7o2LUClRa8+C21VUVMA8fGADTIM/dXTEWuSdI1Qk2Bmd79D1qMOyB6dIRC/OLAmkpVGiEkOTwGThAaXpoqCJA99qamjBcp4aVEyDxSh4ddXFP4rFvvKWo8OHeoc/sRgVqFwdFHU7Vua8BzsVWT5saMx3tu2pWhxmK9ssk8Uu5bScFudkylcCY5eaBd7Jw2THDl8Ok/Gn5VTK91VUB+EqK5N/aJfaXGgIC85CqG1BRIULCKxkgjSgPKtraQkbnIk6gbA4Ko4HBPeK1KES5B9PTU2KZ0TyShz/sJFipGnbcJaACMEnMkrxHYsklAE2hwXvy3vabN6ta/rTYia2uWWGyjVf4gBI2J632NWQdkgwVIFNqpDbQbiBaazYLvhbwX8ziz1BTNJP/ZjJkwMTPnb3cbGCU9L1yOYFsFGpbZffWZjUUE6GZJJVdgRQKNdYub1jxpzTfIAtB9j57a2eH57qjPUNxj/UAYLdtzPYKgGCty38WW6/+/sbsG5gOnt+iZmf66rJsqoDW51Fh7fkFhZ3ac9gxqJoJBpXa80B8L5wRq5hNZq2B4SywtGfwzrQ6g41BnAD41J4VKNa2leHv6rmzv9kf/EehjcKK19Xgac25cEzVvBLkqmLO2s+c76Mw4JoZaE1CbuawG2Y1tLUFmucsD7FwOlmvLu40CCx9h7lHpRRoJ+FmK7oAoPnq/aUGdrLUBPBu7ypWY6nD/qjPqaZDJcimA7VsnIoJI5ZdNhmbFlNV3KtxpPfYjv37J7Uv2aMujg3o82z5HltrtK0HzdrsiN1t22VQiLWUBawpsdMaDfdk0VVRwzUIzNzYiPGxMTfMNFzbTYZm0l772Genr1kDipEgZ6FPg8WgpllqxUrj12oUSBa8aVabgNnNLTFeYehprRNvpDrsbtlwwCp0cV/e9h7UTVzmulmzABb8XXlg4+FcRVaxxmu98x585kq8+b5qYtT3PKmYeTy1+f+qWfFpjQo12AXg2ooSQJY5AjQuagAo/8a8B4oY1iz3zvHYjLsCWT0g3GYYMPKYcbDBwN7diCMHBuLrrz4nX/2FhfW4cv1e3JtfjXU2Qy8F02TMzyzF3CysvAGdLah/yFVQc9DMlPJubU3FFXsdsgHPgPXAmvIw7cXYt29C4BCFtzYbFi548Pb3CyjaNzGmpsLcAnaQPvMYUkxRo4ZcV7cYoFjd8O+cU+QiD2Zmda8EE2mwrpuDiptbnI97rBRNwLwGX9Zzphi6fv2GbCbOnDktpSnfg/c/6weQhmLpwMFJ/V4DQo8cVvO/VJZ9fVY9KkbxXO5MpTLXajXYvWbPpidxBw1+MzilUkNBAXsaK6ycy9Fi9OccLj4ZORmxkIGhrVjd0aHiD2CUZi37ARaawBuBAT7r2H/aJ/p7N+mLvYiio3zSyeuYZ/DGm29q/VXBz2uJbJONijqPfRblrLAcrtsGOdr7tuxfRBjAfistOwA2nesyHHU3+vN+YDnIYPIAhNbh1xGba1YL2XPckwYcY6xsBtzifbg3muuR5AvZaW1uqqDn/XQeas6OVb62UGGopT9frQ3lNdm8VJ6ZSupiR2+sYUU1rCGunFf7J8dj9v79OH/6WHzl5Rfj7V/9PJ55+qnYNzYcI8N90dk/FPOzi3Hz5u0Y3TuW89g8jLITBvg2A29hRnbqnsjmcHNLrOTt6IyN7Y549/2LcenK1ejp8Zp75pnzsb25EVevfBSvvPyyGq+/fvONeOHFL+jM/p8/+WV84+uv6nO8/rNfxV//1Z/H3PyirJFefPF5rZnLlz/S5/76a1+PX//6rbh1+7ZUFrfuQGDajtGxMd13AC81gWQZMyAlNnuTnJfnCrBShJdzDKb/+Ir2Qmc3eXzlvRBLIr7/ve/HG79+U83WSv9EqOruFOHq3Jmz8d4H79t2Svsd28eu6OnoiMOHDsXBAwfj/Q/fj17N7wPw75KqiX2AZe1vfvMbWWzxuU+cPK489Zr2OTMMaFIqoWr5b1t2yrP3mcC5V8PsTVSyUojXk8o583jPPzMhhb+jaSZCEWu8wX4u1YHO5lQZVi1TjT9+VUNCw32tFuM6ec62CEnVfzF7AfBHRxV77927L4BINUXa11ilzYwtmtlWeQL2m5BrYk2pKApsq+ZFgeqyg6yBu6hYZUmbVrcNm0UB6319qeRqN/PLMhirHnJNsaWJ5z0mvKC0o85ZW2XWT08szM2r2SNFi2aUOa+gRmQf8/w4B7H7Y49zpmETRqOZ52s1GioY27jajmQ9ldOZ14q1bZWq5vXp+XqWlu5D2tNVrlw1BX9vhYUbB6wTcpfsGbTShDrX61e+v9Qnauzn+xikbFvjaNi6lF27Ir/o/E/CHe/LfB59Js4ArjkJSE2ixsT+iZidmdF9In4xWxKCGddJ7Y96oeaGLS4siIzIeQ7RbXNjNb73na/FtY8viaB0+swpzQ4iNz904IiaH/emp2Jy/z7NwpmbeygygpoV3X0BAE8z4cKFd2JhcV7+8339g3H58tU4fPhY3L83G9dQmdIMPgAAIABJREFUN9GEXt+UOqLUBKxjiAgocgBAaSajJuDZAqjemZ6Ssq6GSqMw7No18K3ckYYeYKzs39yslrKYJpPU6VstTITnBhDMHmUtatZiAuG1/st1o3W+qendo5jdjSXlQL8AVPv5r3hYd57xNCuoSV1f+xmPDtnylvsNpsH70EgR8FyzUXNuhNYgOtZOFD+u9ckXUPvwK4Ss9XU+j/OeOsu3t6hF3RCgqcI+ZQ9h+bQkIilpF3HMObbOscQcmnVznYFNgL7WbDNPrgX/eD78yJ8b5D7nP76PIsEVRpMK4mraPJ5v1z704eyGYDN3bl5Ts3ap12l+7+O/r3O9qax4Yl4u1olfsWKlrJTSocVWwn4W2r/55nW2+eecT1Ve4r/zfzTpwAtppFXTiNgp8h6q5CSZiGxInM0zoj57KaWqqUXloL3CjLpSBDbsDXlvzn7VavocNBpMtPSsLlucGSdzTJKFWcY9EVzSmk4WUeQq21Y3iogk3MyKY774PTGaRhr7xo3Eldg7Bsl1tUUcZpGyl3CbeOVLX4pr165q3aL8J0deWl2W7Rr1+OeNiiftlM//7vf6DgwtexhsK9lLb17LzDICNdiSSgfS69oHga04KpkUK0HApxkrFFYGvdm0XWK1iCk2NGwGA11zVBmbNBXGldgiBWRDwwyh4GHz3X/wQAf22Pg+HaYffPiBJVo9Bh+5JuwgBGCR2HR2auMXW3Jqaipu37odp8+e1t/RABA7TYy/QSWBSD1hPREokOSSWAMgCPjvdhOAAIXvJ+AZgCHBEUAedgYzCgDh8ac1EZ55CP26Xtj+BL5bN2+pYABIv3b9+iNsJAIyn//KlWuxd++oPFabioFK6jiQPedjnwIq94t/Q8FAIirPeiWPyBzNVpc9Tlq3mAWeAr3sHHPBMB7k9ZiDpKqBpcI8mVX2/NuwFD+Zdbw390UKhlWYFDCaOpTouQCxhQ1BGNCG7jJ/J2AFEEKHc7F12wcfyVVv+pFzAADOlMJDh1kO962klffjmrgO7i/3RezrPBxgrot5uLCg4o37KM/XnLWi2QDh+SSS/uHVTAMKNibyU9h6FAGbm9GTRQOFgcBNWb6YNeb73/aeZo3Zkzxl4eyNBiuTdQYwVfezqUrKE74ygU/GmuqoNPwoC0gpqrEaFfIPdfIphn8C0JLFl4pCOJYBLc8rKIVHxQG/vRMOMx4eV1SUtFODpaq4yeGKYo7veKihkgwY68sUWDDQ9wQFAveI9cG/sy95tsXyZc1ZVZBgfnoh1/NXU0UMXTe6yhrJwyidYJiBb1lyzZhQrEurKjUi8j/ZMqRUXz6r6YFLUcs9lF+mrokBdQaG+KqiupLcui7eQx6WIyM5Z8FWAyQkJCGsERV72Ad02/4IAAl11b37D1RwE0vdZLPiQsA/QIEwJisFlGQBPKtJhfKozY7Xsxcj3+x82R9lsllFTEsdl80TNTVgKaXNEsWPpeG7eoYC2GsGUaoVqkgVazs9rUn47OXpe1TrtIBKngnPRk3urk41ZQHN5IWejKIC53U2+cElWOGbD8BZ+43G4fLyohJEDbtMplgVSWZS2qpLOvksfnkmMKgpXm3lkAlpfk5iGtdaa6B+JQ5q7XTYegZ7gAJiCtB0nPOMlNq6bkR4IDxM4cOHjsTCwrzBkjxjVYjr3lrtY/DASb7mBGSRQwxkvSn2NRpqpYIqq51WkwowVLHJjYra3+4zGdivc/5Jxc6Tkp9mQfbE4uYJP/R4UffEpIrGq+IS6x6w1wBV7VefUZwrzK/oFgioJrMKBDfXKUJq7WnvJGhDkt9LPrKzE0cm+uK1V5+PtRXmUKzF5avTMbO8ERsU//09sW/fZCwtrsSD+7MCDjhjue9+5ratK7ALsJx9jdoRBrUHBA6qwKLo2Ts2rmHgNAKq0eVhobZ1GxvbI+AJoFWMMWYhyJ/c54UK7pU1xTrWIY2qew8faL6P7n0OZiUPY+ikY+COhrOibJSNkFQgnNFu6BLLDh8+LPCNJizsLhQhnJ28L3sSaxiAPjO+Kegcd4jVtpwEgLO9m59DR9yHGSYigZ/ujtjb/t48WdJqwooIzgBil4ZpZyOBfc9rOK4xp8LsdbH5e4oJbX/f1177hlntfb3x3rvvxaWPLgfM5ZolUaztsmxqKd/SvqDySM5DpPmoSX79618/AgZorT2hUdECCTRQ1ABkzThT/BAw4sIXdSdxj9jF3VMM7DaQSK7JXl+T1eiyFBadPZ2xSkMHNSpWqhl7uRbP8YCFO2iwUPfH81hg4Pb39GidAgaR45JbE58B3foGIAN1yO+5LCnE1s25bZXrFyBbjHblYgUcpu2InhHN020UYqOxtboURw9OxKtffC66ttbj2scX4wsvPhuDg30RHV2xsr4VV67eEOgEu9X2YKhtu5VrcJ2QfWyxuRM9HZxHzMIYiLvTD+L67Ttx9fpt7/+diInx8Xjh+Welan77rbfi61//Wly+fDHuTj2I73z7tXj33fdjaXk1/vAHfxBvvfW27FRQzBAXf/rTX8YLL5yPiYnJ+Mcf/fc4c+aklAr/+W//MV750gsaAPvue5dinfxjeyMBdhzgduKlL7wQH398LR48uJdNI59RkGP4PF959ZX45a9+pXtqO1aAMQBbAJSd+OEffj9+/evfqEFYDW3IWyJ7UKMcPqJGKMOyiTFSIgAskvcnI5wPzb4G+GQNKY9HFbR3b3zw4YcC6O7cmdZaOnXqpEA+rHZNPHKuqxouZ1SU8kCzr1C50qzo8AwZrGXsAV8pqs9FSGNipeaMOisfID4x38tK71Kf8j1FBHAt0J4vxp+rWagjnzkV1ZhIsLPsh8oC1LqPEGse4oDsf6iPlpZbw751HlYgQhnCoPdue73bBjPnWOS9qGtsg+mucasxyt+Tb2gmQDYwrHK02pNaI09XxSu+aoYI1+chyQDUjmcQ7GIXi7NexXaa0YC5rWtWYuB9R13CbEbU3RtbkGZ8/bwOdqrYlfF8iaU8P5EW1KDFEqjOd8/nqXtY9q3kmnWWWaXrRony5bT9LUKjWPhpewrAn7T4R47yAjObYG/lyW482au/nWuwntIuK2eimKDi5omuRemb95IV1Wlh3N/nHLqvT/W35kTBwB4eUe1M45qzD5UzijWeJ88Ku1CIRUcOH9HveQ7f/c5X4/LF93Vt588/HVevXNV9PnTI9lDYCw4N9EtRMfvwYWxurMXT587F7OxCnH/2WX0vxMRLFz+M4ydPKA++dXsq9k8cigczc3Hl2g3FE+ICzSEyHVlGj4zE6Miwn7VUBV7L1NPUTvdnZvRvNC2xHF1dWpFThVRWAKKA7txPGnD8WY4Im7ZwlKISANXzCIpI45oLRbTJj/Wl3zdIc8SAIvdzXxXnyJF0xtBUsd0SigcNvUYJueF95eZ2h2ZWMC8SnIT4JucBlDLk/WltUzkpv5Jz8Mw40zQbkFkToyOOOWurqYC2pZtUU9S9W44IIs8x0yfVbtzjxWXX/OTgqPM1gJo8M8+zInHx+vX7/7emxJPy5MfzWzdLnb9WHClVdOVDtVeUKz3e9Ws/lUefT+EAjV3XfJ2qfZr4T53fdd31/cJncm3U9zQ3sxSh2Rx281Pf5dokccLK61xi2nq8tZ5aEdH7NU+QFonE+75LzdgijpG/mXTcobNNOFIST8hvIMTw7nYTsPKq8KoiarD+ZFGq887xXvhn5n2+llKHuHGlXLCrUzlUWc4+0ljJup/8WtarWXMrb0VFn4161as6Ez3vhdcl94IApJkUsvzdtvJifUMqS2ISGADrltwVC0nIELIAHBmOweHBGBgelr2nmkSfz6h45Mz5/A//G9yBkRV8KCtENKJI/l0raFoq0ep8OoC5AJN6IFkdxUTWQL30wIwOBm/3SVYOgwcWJF98L4kPh+/6+qrkyID1sA8B70ggsGAiWSDRAtA8cuyoMCWGI0oGjqx2AAsGPKPdMZfUtq83rZC64uChQ0oS6EbioUuAmpKtE8FgXYc+DEdAhekp+64DPMDeIuFS8p4BiNfnVmDRwIGvQbvYEs0vyFvcBTMenpYlU0Surq9pNoYP0lV5SaPUwF+S76HwozDZP7FPQXN6eloqAJhs3DdAAnzsCGQ0TUj2AfFITLlG3otCjsRFh5+CoQGbnq4eBT0AGsAKDUekyO2ydy4FKyyMsufhM5H8OXibhWoAz89fYDdFtSxo2nYgFJh8oTzhGhhaOrZ3RIOFYAcPMrhKtgyWjMIq5b57gJ8PDgXZBljGQbBCIykHfMFWI7nScDENIcJaA9WCixd+lKQRaT3JKPeR+wSYxGEhwCQbItVh57NuaBCnkxn+TDONZzo/O6dESIB5DiQ2I9xqCViaSuizscOzYAdpjsEGLEDL/gENScTWVlFO2Ldfw8rT65D1xc/JYsEZgZlNj3y1HDSTEfXoXtXhmshnOwmx73ZLqt4CHRvM90oQBNyTyNqzt9UsyYalGbew+Q3Slz9+AUcq4FrXDoZgxpqeaWennuHOLmwXM+JpWJHczjyc16wVLJ8AYijauf5aj1IWqAlgOwANS81Cl/ekQCspuhQ3YYCEf7P9CCAuAIyLHyXkSmBsA6NCLP0ouesaZpifkeSl2OdOct3wUcKdIBm/tlUyHvLK/ZG1GEBfDo1k7XmI+Y5iC6oSz9nYiAf37ov1TJPQygurmEpFpQHeq+tp0ZW2Mo1ksJJPy/h3FU8Vo1CwWdggqxsNaE0fTRUwyfAuuwYlcNm0MhBvFZwLOOJIzrDYYBAdfrQdimM8W34W5ZBA1fR9b81xEdjgBlB9CZhosHQNABh4d9/A94lkrdie9TmJG6WccULswYtiYmIPBYAt71ya3ItivappnNYlXENZPwEsqLhVoUtzzawzIVy7EStSYDnWuBlj9Vc1GzRzJu2XvL7c/NHcgJl2o4KfUaO5BqRLuWP1F4wz7Gn4M3eIs4KmXbFT1fRXo6jdPCSGWink5hyfndenQPS+sO1UASv1GrLrkFev97N9wc0OVaFSbCYxTdPz9pEGxidzBN3PJpkhwZ36e987f343EttNqtqXzV/rOT+eXgkMGujXupPlQ54/2bFqsehKAy9GeRZbgOz8PIz/GnxXllFVi3NvenZ349j+oXieYdrLi9HVPxK/+u2HsboDm3s7xifGo79/KGbmFmN5FUs2q0YpGMhdsHcijup+qPnvOUnkMBqCK2WZCznW5pEjRxULbty8rnVcLGUxhzc3NasKVjrPk4Ke58Tzgi0MgIgFZaGEKANPHD+uRgVM4rL+q0HRXA/xnVjA3AqaYjxvW/vV+jbLC5APYIy9h60T788aEljZ2xtziwvKWWBx35ueVgNAgIoG/LYVLAJDYI91dsa9+/fFGJWFSY9tFcuqrvYVOYpzEyx8AOAWlWPxfdjksUZNVqjZFjVHhebnpu5J+f6jVhGBRmeaGXSAlcSPzS1bTPFaBaJKuZEAJWtV5xwKtJ3t2L9vIo6dOB6//OUvW2dqrW/WtPZxDhVubAWf9TlzByBJjZlcqcqtWr7wBjrZ52JH93TLsuvY8aOxssQQUHzmV8WgA1SBQDG6d48AKdSI5Km8NrYafM46k7DgGISN2M0aWo6BPrPcYQEznJUzk3viM9E5H2z9iqkibKAqY2+kpVaTlCQQtnKCnR3NANO6WV3R/WBWwMbqSgz1d8W+0f44sn9vnD11NBbnZ2UFef7558SSvv9wLm7fnoqePvYp3v/LaoyxrmgivPO7C/Hiy1+Mzp5eKR8WHs5JjcSckRu3b2tWxb0Hc3H7zm01OjifWKs//MM/jJ///JeyDfned78T//Zv/iZeeOF5gZCoY2jWPPvcc7Jbmpp+GP/yz/8k/vZv/zaWlzfiT/7oe/Hzn/88Hswsxv/5f/xVXLhwQWfg+L6JeP3nvzIYn0NiAd2wTWJGxY3rNzQXjXuO9RwPHEUEueCzz5yPK1evWrW3b5/WDbkzuTz7S0pAiAzYXcgG1SAK4DdNQ/IJYovYwxsbAlj5FcY9TS32yq9/85vWTDWtS2bw7BuL177+Wvz9P/yDaiCub24BJdg+zc0oYK7mlVV+zNp3g8o5FUQRbNd4tuQ+YjKnSrMap9z3snMpK2Ffh1mkzh0dZwC7BAolMOhapUeALevUr4myCBAcxrxtv1DFeL0zvHRUzwH1DfePvIs6hj3f083sOQPYbm6j4oKg5hmCBYqXypi4wt+X/Q+1WVncaL/mV5277EviLnsDwMnxh31t+00p2ajRsAFMm+E6DxU/qEeUF7rRS/7IuqGR3NXh+33wwKRqYvaVVNLhwa/UfcQyzjR9xp7emJmd1fVAwFLc2dkJLDTv33+owcujI3t1jgyPjDr2Za6GOs6EwW3Zl6iJlLURsVCqM5j5a+gKfQ0V/+pcl2Ufz25jQ7l8AdKfALsbB3tTHdFuBln5J2W/38RkGPI4wL20AxaonAromifn52zVCLko65A9gTLhwYP7yiellhgbE6mA74VcSJysL4hsgIGckTyTpYX5+O63vhI3b1ylLRwnjh+L69euiWQ3PjERDx7MWA3NLMn+gZidfRg8+kNHDsWVq9d0Ld/41jeV3zEbgWucmr4ve8bxiQMxde9eXL1+K8j+AMs3N6lhevW5+wd6o7evm9Z/q2HEHCtsC7nH92cexrrUtZ59J0Uv8xZU0xu3AH/o6evVmcKz4b7afsZND5MZbV1sgqq/irDEr2AisnNbT0IL4a6h0mW9qVaW2hlsh/s6GgP9VvkRJ1hPPsOJASYHYYM1P7+oPw8PmT0v8qDOGs6BpdhEZaL6CZxgKzbTphmbKeo/ahNmYFbjCpyFZ6FZATp7leU4h09Cl4gQzASjRts0EI0KSWmbJ8y3VB9NoP/xXNd1b+XEbcVUM3dtcwmT/ptuDXqt/Maqj6ouKtZb1dSP59fN1282RvgcVec2v6epDGk2WpoNCz6HMZh2HaZ9l8qW5uvx+3Lp4KZVrWL8yTWJ5kEKjKe2cR5VjeAiRKrpXDiT77rWi6+35r9R1wzqrITgI4cAsIAtz1Jxzb7ugevgkZBmsTxed/OM/Eg5C9asGxt20KCBr5mMbQsmiceolXOgvZwKumw3yfeq2UbDPW27uFo7kVhp6JrEJLyqvVmHfQP9sbmJUrhHNWgRYKgLwJD4LKOje3Qtd27f1loWKXdzQzNqiXPGFPq0J8mLuH/k/tQsJhF2SCWN8vTzRsXjK/XzP//e34HR5XajooKjglAFUXXQHU5LWubi39PqqyiD9abgQ7JDUNIwJQceQBiklxQfsjDZ2FLA6R/oUxInX+Le3pg84EQbX03AJYr6GsaMr6qG1WaQIHmEYYVsnTMP9hDAJEXdzMMHeS07KqQnJAGG4RRKWAAMpm6bwSgPX2wC9k/qGqRO6IHJOBaLy0tpseHgSeAiMT129JiSPt4YVpKAlTyMuaaPPvpYn4kikkSXxBMPbJhYeSMdlO7c0esvLC7H3r3Dsm/g76v4gw1z/fq1WFhACUCw2xBDBiCEgh5rEw0fvv+gNciZ4EaSIva3/PHsTS25WVpHEHQ5ZFz0GFjnq2ZaVJGqRkWyHbUGsKXIeRMC3NNioJgwVVR0d3vwtfw/R4ad8MguqS86pX6JeADbGAZ5Nio4mGRdkOyqkvLpEIYVmM2K+fnZliewvEw1PNwqCoMMnXH40GHZf7iZAUCJndhyWiP4WvivAAp5+cpX3AxNSRGZSZYgl4qsTTdzCpTg/omZKen2hj+LBo0zj8JWAMXkYd3LO3agvwVkCvSpJCfZy4/qIh8DBPM5VHKgNVd+2DUn4LFGBZ35VlOh0JFU01STqane6OrsMVs71QZSQsEmSIljHcY8dwH4NUKjwbyuJkc1GwqMMitrLaJjuw3qzdknVEyC5VVJIElY2YfsG4Pl5etrJn6bxWb5d3mal/TZw2bt5VuMLxJZEnjARIpJK0aaVk8kAgYXKWyGBofdZKBhJ2ueZBbthhLlYrmLeZfFt9l+vqaxvXsUYwqQ5Z7qfsCA7cJ3fNjAcCaGeAnX4HHWFwkRX9XAK/a0ADfPeW3J8d2fcgHd0+sGsADmtB3xejWTiF/ZCxThKgpNc2mFfROw3cSqJgXAt4aWzTPzwFYtGj6dA3ORnev32MHt7KoRwvXbEiqZmTCE066H923toYbs14lvqkKSdQIoxzmBRZgTYIrxts2K2XN+jsSYslDwwE3P0KEA9XVbwUV8qP1fbCExC5OFV9cnJURnh5ovNFfrvrZfp9jbZuSYEWp2uJmMwzpzuG4zd7y+SlFSxY+aDFsJvLKW0rKB803NB4Be2dRQqvp/rMlS4BQTzg1Uqwh5HxVpCep6bkhbEaNBwaUIYU3p3lmBY898q9CKQVbXWk2PJyU9n9ao0HPNBiG/r2fffI3HgYzPalSU6qjsQT4rAfMaTtvAesYZqxRHskqsRoWa0Ts7cWr/cLz64tlYnJ2J1e3OuHRjKuZWsSDcFaA4SHzAc7l/KNbWYHqPiCTgRspga26XPpfylV0pZOSFKybYRrJv12Ny/36dSzTVK6Y7R3AuBamBmAZQxfOwfeGawFU8yTn7h0aGk6TA3IWDMc+8KproyXJzY8TxSXtANi32zRehYRd/bN8M+/iGwEyaKzQK1Iy4d18x9cSJE/reazeuqzFw6OAhqUTH9ozGoQMHVDgxcFWFtxpzvD7AU7cAGa4dJryAybCFHme43lve0m7euUA00EQMUi6S513tDf6eL4ClYh47E3MM5DnpbO7p0f1Gqcd5IXAGxhvQUKnnEiQ2ScN7tuICf0c+CAj/5ptvukjOdaW4m/HFDZS0ocnmXAGhFXsLTBEAnb7IzqGdw6yur5rsACt2yypNziw3/Dty1kY2ZzUXiVwDUGZJeRxxF5BWRa3sN/Bz7rfNJeD/AIShPn0fZ4TnWOAf7matAD5mZexsax0JSIA5nWoertPkGhQbfs6s28oNaB7QWAM4WFmFEIPabzu6YyueOjoR46P9cXDfnjh67FB8fOlynD1/PvoHBuPSpctqVuwd3x+bW7sx83A2zjz1VNy4cT0OHZhUk+vA4SPxwcXL8fT583Hto+tx/fpN3ZuXX3059u3fH+++/17cuvNQwNuJE0fi1s2peP75Z6K/tzc+eO+9+IPvfkdWoDQSJvbvj2effTb+7u/+q4B65uP9u3/37+OlL74Uk5MT8eMf/7c4d/ZsnDt3Pv7pJ/+kuTT8nprgwYNZKRNWVvHHN7DNWTc82BcnT51S7K3mDaAooHqB8xAYIK1I5blhtj1z1wTCwPbes0fXKEvR9LmWR/b6uuzpjh07Gh9duhQLSysm9WSDn/VKk5IG5s9/8Ub0dAMweU4ZFioHJvfHd7/7B/Hv//1/iMGBITE4OZ/uTE2rWTGxb58aHlJhJ/nJ6pxtxQlZVK7ZwqqAMa1f+d+74aYzPi1na0ZF/T1nSjUjTSTwvAHy+lpDZWckZVOCM/yb5zNhf9Wl9arbnTZB1ITEQJ6DZ24R03ZF7AIsOnT4iBpxxG4AWvZagfJqJGTuQK7AfWav1ywKdqXsQdIWlmdV4LtUPUnY4e/44vucs3r2DvfOuVnbg74sl6p5XHa29X38rAhTGxtx/Oghq9w3NjRrcXZu1jVbkir4Pc8EcovWD4AuuV5PV9y/dy8OHDyo+ABoNzQ0GpcuXYr5eYaL98by2opU3xs7KFjJo5yPEopQm3PmcGbR1CG2ulEBUJhWwg2mfTUbfO2OvWXR1ySfVS5QZ3ato4qlum9aGyaqaH1zdmUDv+pM2Ttl7q28o0UiKRFHWwnNtciGeGhIhDmuZ3gQZ4Zxzaxgz0GI0XzGJH6wf/kZFEh8LS7MxQ+++/W4cumSZsI8e+5cvPO7d5SLHX/qVExNTysP3Tc2HkzEfnAfsuNKPP+F5+LDyxfF2n/llS9p/R0+cFiWqb97+51YYs7S+Hg8mJ2NZWbzUWN290d3D0ScEJuaAd1YT0G242RBrUgzAzUIeYOUk1jECiT1+bCVXvY8Tc4/nikxn9hTavlS67LuRJTL85U96YYp6w7bbufW7C1qKO61iAid5DEmmdIg4fXAcqrWL8Cdfwf7cJ25o9cgtgnfGeiLTmyjlKMzA8M13tieEZ1NPCc1ZVHey6JpR6oTz63q0s/TzFds6OpSHkaDyeflpm2nci6cZ0S6BqBvQa3U3eU5TcqhmdFaja+WBZlri8p/m43KWsOPNip8jre/mg0Mx4BSFjye/yofSsJDMx/+tPz2STmzcqiMRY49idvlXq3P0bx2XXHiENlGSUtgk4scE57cgDHps93Uae5vb0sTu4Sd1fnwKAfSdW9LqVPXa9IpsZIZM6rlcqA7e9TzZ1g/A62ZFeQsnJconjnH3NjkXPJnKBIJGFSRw5SbiszHTCWrd2udGWd049aYl2so9ko5gLhBS71UMzhda9CQqCagiJyQizRbizM5CblJBKvzpPIv3ou1q4YGKtyurrSV7xLRmbziheefj6k7d0XKBq/UHE6U4EePxtTdu583Kj6rKPz8334/74AaFSXZanASW8HMkayFZgm4w5KnFwZWm0lGAGHTEmw1+Im5Dmtr+r6BQRdbsnFaXBKzi8SZhIqAwsYEnCSBJ2CsLK2IBUQSymYkiZiamtb7HWBY3c6uh153dLhYQs2xthp9SG3TWx7GP8wcWEuw6lU85KFNgCNJEVMmpWpIbUnQ+OL7SNYJOFj74BVtRcWmOv4T4/sUQFB9AMzxWQEakOJjX8XgPYEzFHc5ZBuGIoDknbtTGuhN0Xvh3QtuvOD9ynCpETx7hxV8+IwkmjBrH87MKkHnHhOQAQ9IDJCv8lnousp2aXnZfvWyxCBQmx1fbIhinVRiKIa3MAIfSh7w2D58zEwx0FQHGr82wSZ56usZuuHDMG0YEbr343ikzuoecQ0wdUg0ensB7GmmdEtdU00DvU4mFvV+HFAaIYtUAAAgAElEQVTcAyWnKu493KgYj4CT8t/v9QBbDjGaNzwPwAUNHUxWGA2DiYn9GsxYgzwZEkpRLTB7DUY4stURPVvuMWtW0nNqeIAC2Mf4olLUiJlsYAUJNQcYhyrrjS+SPQp6BsMD5JZKpYA7eTDX0DNZdxhQ9dejjQp58SbYVM+jvrcS/koUWs9Lzpt+nSomZNeUAHVrBk2+I0zGAvyLJaU1kMUHiba9Fnt04LpBV36y7aRICZEvxkzq8v3dho2zpaJheHBY7C+KAS5nYX5J38v6VlwRiGZLBDVKEkQRi6fLlkYaVjc3l6CA51ZIGrmXAXfrtr7AkiQTGzOxN9Uw4lloyGwvRXF7LgLrAgCM50UcAChiLZgZbEspsfdokiT7VpZLmYhx37huS+DZF/Y7FZAOMNFnW7ICikmMANqIdyTrNbSdmMD62Vjfkg8+1y6v2wRF2mvE998skHwWmUDyDKzcsU0OzwXGBU0Y3ofmMuuh7N54TQpSXScJYbLTtL4ZFg1jBZ9bDSwzO5tnrCSuq8dMDwbVzaEAeyjIsAr2AuoVn9JSTMl5AvBi0RjvyXVl/00A4GpU8L1cF8/YVmvpq16MyXxtW2Ax08SAnJ6JGD0eRF1f/LytnRyDqlnEd1D88+s8ip1kGxeAXqzreuaKtalIqMKY2EMcf7wBUkBPC+xhjwCYlhXZFgzpPR4qv7FuMET7PhWNyWTjbK2ipH7lNYk9rPtqVKgIkeWfAQQl1qhA0rJRz5CiMwFamv5qWKRfeLNQazYjPivbaRZRdY/41Y0iN2web2zU6z1+1jTfx+scJr3XY4HCn34tfp8q0Fw8w7z1QnuSooJBlIdGuuMbrzwX66tL8WB+NW4/XIy7M0t6Dtg7wKKcW1yJpTUaoqE8gpjDUN7bt++44Y8qKjqlTGAdMsdBg55zHghANHmU7C77+wW2VWFH/NP+2tqK/fsn9MwAntgbNX+LfIX74EHzxDDHTnIo8gNia6s4TBZz7QuaYbLYyeHsGygKsXtQjkO82o0vvPB83Lx5U7HpzOmn9Lko1E49dVKg6e27t3U+Hti/P+5N35fVzp49IyJJkE9oCHKqDEgfNndCYLNBdPIBgBU39ur5cL3EWJ5PR4cLO56xSA+5dqqRUGuAWASgJsVXNh9YD/zMM+eeUcOQ3OH69etioPn+2w5T6rtGYV/2DnVe1lrjvQFbAAurUVH5TgGT/Lka07Uea50XQCE1UPq4qxGaAyhtV2ZLjLJcIp6UlaTYgTS3BmwNIFsD7gmNq/4+scNhoKNoEeMdgoyYrFYtl8VVi6maTHbWFa+tgZxSpbkhUao23os1D0momvCVdxVoKBZ42o5VHqecMYdAQzbq6+2K5fmFeOHpIzHS3xn7Rgbi1KljAoeufPxxnH3hhZh9OBvrG9tx+eNrAuqeeuq0iEq/+vkv4vnnnxNICuN4+v5MHDx8OG5euxkX3n1f++HFL7wQBw8fipX1dQ3Q5jXOPX1WNQdg/DPnzmmPXr1yLc6dO617/NZbv4tvfus12fNdvPhR/Pmf/4lmUkAe+spXvhwL83Nx9coVzYX4whdfin/6p9d1rv/B974b7733fqxvbAVMScgdfF7WGD7yNMRQSvF8eS6aw5VD5QH1UUpr9ssqTbNtWahtrjOo03atX/3aV6X0gClcLAL2LXsShvLZ00/Fu+++p8Ga5EYVRzkbzz59Jib2TcRv3npLeQYNSWICqmPqhzNnz8ZPfvK6gEJycYZvsyexxOGZi4ShuT7t2V3N3NJ5TXnf+8ySRUwxaKUk2NWaUlMVdqdqB3KwVKWLRMWe7nW9IBCq3fR3ruT5FiZsrWsNll0N85l2tq2yZf3a8mUtBoaGNVhYszH6+kTIuHHjRjAnh8YMXxqSmrFQ6xilqqwrXeIWUO18wHvSSoeGMjEblKV0cR5IXmhSBvlN2bp6tki3YqtzRz8vq6ysLmznB+R/boRoriN10PqK6mTu8YA+E2S1Ta1N4hq5I/ka95DaknOEwehee6v6vOPjY2pIjI2Ni7WLzRl1kODDTrPItYeJr9jVJnOf69a8vVSAs9Ycx9oN42ooVT0j0oVmv7npVrlf1SWPn/HV2GgRxjQw22pX/V+uQ5TZilNlESacIZvcqQxWzMmaQ2B6zvwDIORnuTeclcRRhj5TmwL2k0ftm5hQfFCjOOMr147DgpriG6vxrde+FDeuXJGi4vnnnpX1Ew35w8eOxez8nFwP9o1PxNDAUCzMzcXCwlyce/bpuHLtqpwTvv3tb8d7774bI4PD8cz5Z+PSpY+syBwcjKkHD6QSWd9kzUFAswoRYHJ8DPtTZt2salYVuVvHLjn9ruYr3L13L7qZPZeDxft7+62oyHpR4C2McM461hz7XEzydLVIi9girHGPAWw9F8PDs7mv1GzkFWU9pYYfqoy09eV5S/GUVqT8yr4q1TZNVmKQ9tLOjkgDyrlpiC0ycN5OCawlqz7NHCdHVx2imntN+5VGBbGTWp09qnWi92XWheca8rOsQykytjyPAlfrvp5O3Sv2DXNPOSNKDWD+l2H5x0F9gcwNRdUncs4Glt/u4X12o6KZJz9eu39WPvyk/Lpq9IoplR89vvcev+5Hcvq0c2s1Y4sI+RhnspnfSCHRaFpWfFWurv1sEhe/Lyvpmu3TzN/bqpR89STZsO6wP5VSIBOpeg4mrzEXx1ZmnAOd1NCZ5yvmSpThh8Ne5jXIcWRjl034qrmrUVpx3GRfO2CU1ZysU5N8BPbGtTgn9X5i7/Cl/C6JvuxBNz1smScicBJaSv0KQZsmmxTSHaG8H2t4cvIa0M17QUA6//Q5NZ3BF8f27FUeAl7J66Ly/FxR8VnV6ef/9nt5B0ZXzN59PBZV3FVJ/xh7QkAxLNHcnPJ8p5ufPrwwVgA1KZo58GDBHz1yVAf27Vt3W3ItissVVAtiLEecPHVShfuD+w9VYMAO5MABTL5167Z+f/bsWYF6WD+x+Tmc1GHv6lSjgWKMAoeGghmzWwKba/YEICTWQLwe6guCE4chgYNBdADcAJTHT560D1x28gly2AlxDQcmJ+Pq1WuyYzl+/JjuDwk/0msN1sHDPocY83McrgSitY21mJudU9GLGuLjK1dU5HGdYn0MMCTTCbbsYdKTlMTCtjjbsbTk5JTvhwkF4Q1QliD24OEDWTLpYNDzMTMQuasYhzqIaKBYbk0xw8/KripZQGKAlq9sefk3B3FnMlJFPM+egrqVROZAM5okz5w/L0CDRoICupL8LhVwAAxrFNE0Kxpsphp2zppUwyP9JDkMa2BceU/yPXxWMUU0QJtgv6fFjOK+cq+GBgd0byRB3DFru69/IObn51RIwrres9fNLD7q8NBIrK6ZOVRSPcAnWeAky5MDqZJyNbG27Z0s1lV3l4pBrMAoDu7evSOPa4auak2m727LgiSTINtZuFGRZ2srpjSZC5VcFHj/pEZFNUWqMaEDN599qWRaL55vVuKAUhuUvY18zNOupQ5WJ0LZVGn4ljaLBTWWkmHGHtvepVgz64A9qeKgp09FPsPpWZPcM3xMiTE0KUkyywOcf6/5EtxH9iIMHYABNQTSl3Rycr/811X04gPOEMe0E9CzH2C9bOs5KKlpWBK52LK8EyamB4ruSMnE9Uo1A6iUID7Jd9lfyb+517YaBbqpOM1mCYkRVhOSqq6v63tYc9XwMJMOliEqKDPcWQi2HjK7rxWLW2afbhaxh/zvqE52oxev+LRdqWHzqFZ4SQpi1gIsrWIZiWmlRoDZx/wsMZP3c2O6N/ZP7JdNDaxfYkoxtLkvJHKadSLhlT+X/KUTWDYgaG/OSqZLoddkHbZV1LvyaaZRwWt5OGdb0dQGx2yzIEuuGnidljKA9rKsSXWAGqEMWpeFl2XvHs7uWRW1dvn+ajbOLSyooGn6xhrwt/WMCxoXhvW5iM0oG2jW8B7N/cmeaxYTKswUZxl02xdb6+sCFTSIdZ1ZQDBWc+BwSpJr7VbzsYoRnj9nUDUqan+XV3F5+ysWuI+o56EzC9ucnGlRiXSxsppA8j8nyXm8kCpAgusrcIO13yz8mj/z+P16tDBypvLPuaZKW2yB5PXBRmrlNk9UVOzG8fH+eO1Lz8bu1mbcmp6Ja9NzcW8eZU2PCAV7xsbj/sxczC+txtBwv4ph8haaEij5YPBSXHAGwDAnRpBX8AWjy8/V1gSAITQAmaHFfTcwZP9zvg+VqVhhyfxnL2JTyRlaDWPWD2cg93eTgmhrS6/HV6sJlzFOoOfWtoAu1lGxyxTfs5nJzxw+dFCsdgAvVBMwlCkasUBifz+YfahGz4GDB2JxjuGjA1ItEpMBKCgaxSpPuyDAAZo1ahRjDbS8koNbscfCwpMZYNjIEO9RlVp9WMoGrpPPqyZlxiPWUFk3wVonZrInADTw9oYdT9zme8gXPUzbKkENeRSYXkN5/V51thYgXw0IZnaQjzKjohSvtWYLrK91quZ8NkBq2C+/ElsN5GBh4kHuzr2TTADBBNA3v0cEjzXPrxKYB8kAQGoTqzGDr7LvXGHmlxUZVThXc6L1XHOekchBqabVNSrXKxu4jGHeYLqPsOUBMMkdnasyo21C7y0mXzIE6/1khZDrSpYEnJ1Dg7G5shTPnz0ao/2dsWewJw4fnJStE+f7LoBp0CTB6nMTSE3AEznk8OCAgFsNbB8eiS1s7ZZWYnzPuO4DjFhYxU+dPh23796Jm7duaw7F4cMH4sSJk7q+99//ML79zdfijV/9EiOKePmLz8dPXv+F9tEPf/i9+Id/+FHs379PMyqYNXfp4pX4wfe/LUszhmh/5w++FWvr2/HTn/4svveD78qqhO9jra6ubnj2TJJZnnnmaTU7sHYh/nDWFPhLQ4hGBPZhq9iAyq7QjHUsBrFY+/KXvyy7KZpElfNVPKS+YbD9g3v3VANR55jcZVUj64h9oNwIskUSKaiv2I/szYsXL4l1iVLw1MmT+jtqIc453kcAfCpDBapnDGEf1znJ3/MeBqKsqhCxAdaoOG1uRFADFtlBwFWCo6w5WS5CMNO8OmZ9mNVMDkGTgdSS5i97eg3iGKShwSFZ4GigvJoX1D2o2AZ0PwaHRuK9998T0YT8jPVJHN6VUHFXeT75SxGOONNXV5ZTMcxcG4bs2gqumuJiW4tAZMJONUzLSqr2m2aZpZ97E9jy3B+zwk3q8F5zXHYNQV3C69FQYv+QT/HnocE+2TQxoFmfvdNEBD43hD+u38Cvm/GyIQW8zVkgqGCxOCJ/JA86cuSYatZr165HT0+/vp/a2Xmc1XoijIhU49ljyj8ghVArrntAdpGX6n5U7cfPc/1cS6lQ6nsrVj6OJRQAXPmATueyGk7CTw+DzxukmWoMEkPrTC9WdtloteN4p7AA9gPNfs00GBj0zIqHEMg2dQZDKuHMoHFhYk+XcikwAMgIf/SDb8XKwnx8dPFSvPDcc1Ib3pm6E8+++HzcvTdtq+qRPTEyNBK3btyMvv6eOHT4UEzfn44bt27Ft771zbh5/WYszMzFyy+9qjmUiysrMYkt9dSUZuxs0M1nRtFWAf6bcfr0yTh79mTcn56Kxbk51fdLi8s61xZWVuPW3TtsQJEkW40xcjrZzZloyR+YNUTOyv3SXE5IR2mdxt6j1lJDFZso1iK2iOQTeaYqvsD4Vx1ogmkVqpodCCm1ryd2t002kO2PzrK08cGmOa0PIWNWXYFtFfaxjp8m1Wi2WqrCWd/sZ6knd4j9zFTyvC6+b2WFRia2asxD2gk4KIpHqCgHB+2qEDuxsLCUs5cAqrejo4sZLX2Ki663PXMF7IPn3yb2tUk1jzcW2vVznuMtEK1y1KrjrSoowgIFS7PmbBMaHh2G/c/JtV2LtFWcdVZ8Wm79SGOi8o+MS2xuqQbSMs4qgsctqNtXpbwllQ/6bDup+G4pQ1y/2srYFrl1r/nBVk3Y+AzNz8y1glGxVyF+qZ5NIrLsw9eYv+TZbJwjKHelDk6rOPaKlDKa/9XtXDQbJqwf4iLrXPlgkSOFb7mZoZrPXSv/HN+TeZBwBWykRCB23K76vAjc7DPyZ5EG0h5YeCMWowytz9yYtc9eJb9kHxGXSA5pSvAcnVPtKB5RZ3Cfb9640ZoFJ0JbX19MHpi0ReLnMyr+OVvn8+/5fboDjzcqKhgr0FXi2mhUmEnbBmXEmsjp9i3QJTrE9ge4o8O3srokH1ESR9kBbO/Kc46NSCDj93i4HTx0UBttfm5eViP4MFJM8DMwpUjSSDwpdhleJYBQjNFO2T/Z27gndrd2lJQADONFi3rho48/Fii9/8CB7OgvK7GnuFai39mleRi379xRkjW2b7zFCjOLnDkCnTE7MxPPP/dcXLp4SdJI5FbyfcyBaQTXBw8furOZdjuwmmjYcP1cs22v+ltgAoAFBQP/0cCQfDMBeNj49+/Z2olky5JyvO76VABy7/h5gqKlx225IveZ58W/9aIEUKHrgXhEYIAQHrPsXCTNzkHALbAcexgznApws6rB8ZvgTSJDQkB3l8JNDRpYVttbcfzYcRUh2FYQZGk4jY3ti/sPZvTcxApaXmkxhYqFU2wAHeCyjshBnbKy6klbICepBH6Kj8yadK0a7FUyyA4aHtWQ6pM8GqY2Hs+w6SjsYLc5OfFgULH6YXV1e1CqGiM64NxdX1zAF9NWT1yrpIGyPNuK8bFxrRUOugOTB+LGzRu6z+yTGtokL201Tfyz+jeBnQ1aRnumeIuFVYd8gXRStuQ9qgRExWYWmrUW9B7aw7a4anVBGsmmlypMaydrAjjSyqZA+QJk6pC2PPNT6RaPMNENvvG5/fY0lQBIKMhZ7+xpWLY06Hhf1rKGnDNXJdlTHn7tZ2GGQ6jhIVadhlGbHVr+yCQCKvo0BNAAHgkvDapqPpDI86w0wLm7S8kP7CuuyQ1ZF+g8W/mh0rTZpTlmCanBcaTRbophRUfCYi9LJz08D4p4qcpgCaVPJXua4rmGffFrKdPMbjQTUaJp1meBrYaZW0o3cklbUFEMmBWmZmY2EBWf0u+3bCeQgi8uLrSKlmI+EaMA2YnNFGncL54R8YOCj7UgtQGzd9bWFGNtjWU2FAoi3o+mtD5/zuVoWT+k16wKg1w7xVbh+j0Lx8ACRTaxkvjGvldcTOWWFT2NpLml0oAx5Zk8FF8wws3k2VWTgkJGZ1Ay7bnWsnrg94qB+BaPjmr9zsBY73ajrn6mipp288LM8FKHsB5JrrmHBVjy83w1mU5aF8lIVQzu7JLn+KFDhxQXWcfaa9zfXEO1N2vXFWux9iQ/y2e2hNkARgEolvkzrtfMz/pSE4xmSRUlFHuplqzXqALoSYXOZ+U7ev8EgMWga1li+Nqe9PVZjYpmc6Zd9Hz6FfCZm5+hXUt+UlHBed21uxOnD+6J504fja2N1ZhZXI97C2tx5+GCm/v4IY+Nx8O5hZhdWIqBQSt8IB/AiLpx82arGcfnRuXHnhZRYmXFhdPWduZGq5rPA/gLeFge0UUU4EyiYSBFAvEk1YbEF3IFXpc1xj6sWHz8xAmxa+/enUrGMQUVxZzXvIdLbot0AShRYH3Z23HvORM5x3SWdHXGmECdGcU+zc3Z3Y2ZeeduFJAPpvE+H9GfaxYIZyoxjxhEIdXbNxA3b94SQKu4jsKwqxqP7SGqUlhIgWcbF77coMQiEPXAmvJIA+PORNRs0SwjDzzU2SGwdjiWFhaVx3JdNHe4Fs08as7myH1Sa5PXq4KS3/N6WHAdOnw43n777WQ9285O6oZsENT+biqHHNPMYhWLs+ywiOdprMBzd37gQeetvU1MzcZmeeXL+iyJOXPz8y07D81jSuWezrMGW1vs1lQ7C4hJa59iBNYwbrPBYZp2xxpgaM6uwKKI+F37WLYhSeKoGEUM5feoBTkLiSdSwqCg7WYBr8T4UG8c3b83YnM1jh2aVH7Eeb6wvBI9Q6PRNzgUv3vn/ejs8pBU1AF3bt/QZyRfoMlwf3Y2cHQYgeG7ZHs7Grl79u6V8hgl0a3b0zpjWS9/+id//P+w957PdaZHlmfCW8LQE/SuaKqKLJWRqqRWq9RG6pmI3p2J+bYb++9NxMR+2d3ZHamdRmqp5aXyJKtoQA+AJECA8H7jd07mvZcoUr0d3R9GG3W7FQXC3Pu+z/s8aU6ePBk/+MEPJKv65huX4v/8rz+M9959Sz7sn37+cxU4kDa7dvVqrK1vx/vv/0n8l//9/4jRXUPxF3/+bRUx0Fv/T//pP8Q//OgncezEUeU/v/zN71RkkA3LB0ZXxNfffksd1Y+fPM54zj18zIXBr5I7fPbZpwLqieNtmwzsE3fu3b9XMYjYnQW49fUp3uRjkAPjMzmLvK9AjPJN7ZYEREITKTCeE3kU+xE51JOnTsaNGzeip7tXdoNO8RMnTugM05UkGYyUbGMvSwYmmbFFiiG+YL+W/BnMccDsQwfHYmFxXn4X30VnNVr6VShlrTibPsvMtjIJgiIYv2tgzV2ojudWYtfQoIgs6Mir+13nwfK7xClFVKshpL1I+oyOqtDTN9AvmT18IUx3gORdQ3QquqjnmBhSBwVEyEUUI4gdXUDiVf6ZdSxihHMkui/5yoXOBqiZA519Dy0dZbxXvmfF1xRE+HuR5NI/ShpQxccuF9SJfdOeIYPDevDiXACAkc+yCSD70R2rQa+d5B50gg8oxyEPGxkZ1b0BbkPCosiGPW+jACkpN89ck6yJ7LJnUrBWjkO3GnlmFRQqB2kFRF1EcQxVuVxrvNDq71v/3vGU7Z+IQduOE1gD+eSMLRvF35IjTimV6vTBzhcponJa9gp7AlsEWY3slbyTrgrkm3m2xEwUsfERxOOAoYDpFDCQdertbot//1ffjf7urph6OBFDAwNx4+Z1xVUHj4zF+N07mneAr2P/P52e0TM9euxYfH7981jdWI9Lr78et2+Ox/b6Vrx64bV4cP9hLK6sRv+uXXH7/v0Yv3tPs17a1LPhQfXM7RwZGYg3v3Ypzp48Hvfv3Yv7d8kn12NoeCQeTz+NWeSswBQyBkdOkZIlksqAs+uba3q2MJRMzGGoNTNDKSyiq7/qQjlrl6QaiJXYI85bEdOwIfKh6i43sFpEgSp8g10Qv/LsVVzPPEjypZD4FIMwV4D5U91B98fc4rz2jHNhdyDREVjFvrIJYB0lL87+ovCHvcLOFQi+ssbsTO8hrk2E1eGhHI5tYJnnq+KWunR6RETlwyheFPmytaOiigg67RmvvjBuTUll/16TfFCzHJ8vVLjjsLVIVxHsl6SWWhnDO8Lc1gJH4+//uc6P/MUX3osSKoPy7s4v9QzHYTtfzsdztmA6wfq318ESTn4fbGVznphIOVnE59mri7Px8mezRi70mgDKXpRdyefAGSGWgdArUoCKUnT/IJu5KflanjVnUn4HBZZVfGuHZrPKzuMz2dPK4Zlt4VxPpAzZUnAdKylgdsCHFJ+n3WdPkaPyPc5HzXjVnFw6GXt7nAe309G3JL8/dvBQUwZcHUTrkqIj3963d68wz/Hb48K5iOUpEEOsJV/vbO+MixcvxMyTafnE5cWl6OjuVGcc508xyVeFihfu16+++Ue8AsPZUdFqiHUod+j01fesAexqqIYqA4BnW74khnp7A0azGGAp30Q0NfuU4XkYnB47P7FtLMlBxZvgjDZVtbeuAQ5vKrBXS2FbuwwLwTIJCUkMgQXBnmRIkmmq1q5tKpGzCiQJTtBeJXmiy4GX9OvaO2Lq0VRsCBw1Y2141y4NHZMsEMC8hhBvxb0HD5Rw81ncN1XaQ4cOqnWxI7WWSarvP7gvCY2zZ87G1WtXc0icq8ywxAtQpf0UozsyOqJ7IJEAGGBVNTxwYCAePZqSUYfFR6D9aOqRChsAu9w/xlkzOnYNqsJqSQM0Vq1fKmeXXREFLit5RBqhraknjDPgOZRmfTFjCuzWgpler8BRIFcxMxMMx1AT4DJY0xVnt0vDJDtx/Liu+/at29HZ42FAA4NDSjDVptfu4XGlBc3HiU2RTK6GNm0yLPBGYvpIFxCmmq+NhMpSNXZGAJsEo+whgG5YILDUkVPp6x9MljqyMIsx83RG70cAA8NcrA6SA+Z6ACpl8iEt2QyAcFisp0AKASqsuxn9VMUJBikgCbDVsCScVTI2cyCvW60J4NxaK0mplqFVBcIq0G/MIUhH3yhE5HD7lFJpFDBakmfh2S0FEAL4rJ85oso19Fo2GR2cS1g4rG0BMko61VXiM1/Ja20TvUVLdxbPlZflJLhWEhAPq0JeiyRROqipFcl/6TxRW6YG3cPaR17ADB6vkXV/OXOsN/dQMlHaRyTbuXEdHDGjpJhym7IJpSWs69YQRrPGANfoJuAemqxZF0UIFgrAAghnr9deLdBAXU8MEF1da7AHa50clLooyzqasbRmiSqANdaawYf795tJIe12s5w9lMyrrJb2BpTlc+A2bthGDFA2KAYbl+KCCyTWPTdDBbai9yIdXqUFbMkrF1H4PCTbLIvgZIXEbWR4tPG3FC8IvEqLmOvj+RBcAcou06KdRWTtpeyoKPYfd9OQWkr7gm+pdmE+U0PQ1pDP8HC9GgQtZlcC7dUF0WqX1KHX0SGbjn2tPVmt3QrSxfDM4YLJtOGaa29T5OA9KLi0SrJ5fat4lk8lW9y131jjbusb15yASihUWMzrLmBGAHIWMLiX9dXVODJ2REOZCwRUxw2zi6Sjuq59U1rA9Z6lEU/SDSOnmI0KqFMKsOZb4CMlDqiiAWfIsh8GTMzabrDaGtqy6VP+UPv7C+KgVkCiAJ0q2vxLCxUVo7SCsC8ramh/vWwoYrX37+ioYH91bG/H6QPDcf7kwVhfXY75lc2YnFuOe49mxHQcHh6MwV3DsbS6HosrgDuWEcAOScebIeWyU/aD8hVIc8zxPJGXQEpuyT5ha1MdF5zFmqHlwoqNKKlw3/4AACAASURBVOdwbOygujgo9mtQuwpPnbF//wE9Y+ZUEL8A7BFHoL3PngWsbHTVZYeRChW5BykswMqVH9tE27yAwnbZjsNHDsfU5FSsrixrfhcdGgAbSNesb67HxBQgz5oA/IkHE7Fn96hkStifXHtJGWHw1UnT1aN7MLhr9nez0FhsQ3ermdVtUL+SVJ4n/1bXSLLqWI8qXpj95qS5/oY1xs5637TrXPBfFYCZ2aXh22a8txY9FVskaOJOjzXNWGPNP/7k4wb4WmdOnS0lAblTaiyL+ewFkm5e2CeTEzzDxN0yXo/2HJYrAH5tXXMJ6qW5YhQJKCSmTJPvP/XViTGqsy5njfj82Xe44IW0FnG3/TqfT/KrLld1W3iWGTaDZ0W8rIhfoIMHXJYNaxRCU/6Jzzp69Jj2h4YsJ7t6Y3kp+jsjjuwfiaP7RmJXb0d0bG8qKeeef/Hr38XJc+ejo6cvHk49ie7eAQFbkn1dRr/c3Uftnd0RXOvqmuJgSEZmCrtLZebprFizd+9PxbFjY+pqeP31VyWBdP36F/HN996NJ0+m4969B3HyxFGdlZ9LWuo17aP//uOfxnvvfUMd3//w9z+OP3v/W2Ky//2PfqL3oRiJ35udfRa/++BDxfvra44pOLLEj3R801FBrEvOglyX5tQRO1OQYKYTjOTs8mIta4g7wDJdhPJZYvZuemD2avrAzk6tGR3XrC22xmxVyEhrcf7cK7Iln372mYGe3Cc8/rHDY3H50uX4wQ9/KKCb34MVzt9ig/D97py1RKL2s+Jngz0uBroDgPipvkcZhr89dfKkYp7px8jYeAApAI4vxIEhayDWfhtr1as8h9iMc2iVH9tSPoPvO/bZjq4ex9rEQzwnZg2Q15FLcfaI4+lSVcFqaFjxO8+APc1MBvIvJIsqL1JewPw5FQRsbyVxRnd+ntNWYoF+N6U86iyWXEj9TEStnG9RcwA405KZ095w17el7nJQrAbUm6RTMSzPxTaa2SAuVPA1NpnzCIjFtSAPSXEJST72wtGjhxsyUAJiJS+FtJVBOGwJsw2ZB0Ox4urVqzG/uKQOpaq0YZex25BNeFaLCwvq2OeFLPHyMrNXTLioeKuVvAE5o+RVKsauQsVOYLRyzCL7lH0XqUSStbbjkqlsIU00wGTsbBZ/nENZfrPIQdxzSeVBeOEwsG/4LyA9km4Ua/BhxEz4X7rfyS+JX9mn+/bt9yyIzvb4s+98PVYXF+L82bOxOD+v2TnXb16Py2+9EQ+nJrUuFIK4jpknMwI9T505E9e+uKa99irkxqufx8riSrz79jfUxbRMAbi7JyYfP4o79x9qzgQs/7YoPfv1GOhDirg7Tp84FhfOvaJzdO3KNcklzc4vxuz8guRu5jXIvVMkTWJYJCwlPU0uteW5E13MO8LOJ0BcJCh11WWnD3tWRcUqdGfBsjW3rKIj91pkQZ43exNbW4Vs9gLvLakpzSoiR3DxneshR4fcqPemE3KNGZEehK55oBBiIbjRjdHlTlN8ArkIagvYYoo2RUZRnqiOSsfHdFh0dqCewFymPuV2nBX83xKywNuhzjLe1zmbc7Da338ottwZu5o65oJP+dvylWWLqwjhWMPBZ30tCaUkPjTD6Ja45AWcnjpbFQ9XfPyHyEQvi7l9Mf5k9ofyaq1Fa0b/fIDfms9U17LvuUhI/lvnyZ4HUYSZ6vZzPJbzaPLtW9enumJUTM5h7/xaxXXyUTkUm33uYqUJh/3K+y3/xJmQ5DG5dI7FMD7UvD/jYLbPLiQ3Zc69bpY5LptYhVP8urt93SUIVlR5O9fEvsSns5dLtpy1gywBxsk5Rc0FDBG8T0ocu3aJmIx/x8/xTIUl9fTEK2fOxu3xcf0O987vrG6uK3e/d/f+V4WK57fpV//6/8MK7GFYTA4ZkoEjwAGEUzXRbAolcwUmCYix0XDCZya+jW7+DOAsq7Fmo1AJdTKlwkIaGgUdmxuxtoZGa4cGVRIQkUBzODnExdC7fuOWkrmzZ1+RdiOBhQOKfjNlc/jhCowZAP3hITEcuSbeg/d7OPFQQUnfwIC+JngTO7G3N/p6+sS8gKUy/XQmjhw9KuY8jAqMDcYPhv2eURdTeN/ZmVkBUtzXzfFxtcQzE+PhxISAR6RjpJO/zRBvDzlFi5puEwzqszkYzbT5mqkIY4AA5+bNm0oeSIwwxGbHhvUZGd6cM0J2jxrUZR1wKvyeCckZCEsSxZqQCig72sUgYD1I8iyN5eBcYIsY9w4SC1SSNnpDU9xyCcVsL715ApFK/gl0C+w7cviwBl7xrGCaDw0PS/YBzWOzms1oqv1Xe6iSoJqDQLKGo3CC4UAZv1F6tuwj7kWM7wywmixpV9AJgPi8vr4ByXSxto8ePUkg0vMDCKI8cNxMAZL2pmM30MyLJEoyPZq3AXi4GhvMwsiA3m3PFI6Y0cLsFndiuOZQAYqdeQUVCsZbGOJ2iq3feO6HjTPXYGUkG1LOtbSDs6W+EXxkYOl1TkZ1Xpjd9ZfbPIt5XQmAkocampdaUcXEFjMiAdACTHCeBbgyrBz9cZguDCiu514seWwEiTqBpfRRccLr7jIodoafgYOhCpSKqcezKyYRz9PJFKx+S3GR5BZL10W5DRc5E7gsloTYcx0G+SmYkMCK4ZhgEgxAJ4OewyPmw9xcdockWz/Bk7SMvl51HHhwPW3mnEHOrFjNSBf09+v+Hz95oj1Vyb0C6WRgmjXsIirbQ50GWaiYmXnqQlJ3p0H+1TWDRQnYSuYnC7gk6QCaSLYwq4N74tyy1jwzkjrAoSpmMf8HEECF6a1NsSZJFCqB4Vq4fj6fYq8GcQq0Nfjd2M/pR5TgJHhjeS/AHjqTHLTyDGDosZ+wb/I3sMSSvexZPF7rSpaqIFJBMH9P4FcgAOtenWECCZPNUolSyfDx+zwf1lgDZWVTXGDjZbkG26+GLcrOGh4aCaGlBWb0bJxc1761Ldb+Sb1vFUzUdcVcIQN4GorL9zQM1fr1Lqjhky05VeeG91HhSzMP9ui/rFkjkTAealBUCIBthHy8hmgbEOYsqJApQLs5S6I1uXlZEvSy36nvF6BRdtzr9vKOivIFO5PFLyWILUOWv/yeTZvZAEwalrO5Hnr+qTHevr0dR4a741tvvRrLi89yRsVCTD59Jib37tFhD2neilhe4zlQ+G0OJ4e5q240gURo1ltm4smTxwLUSr5IA4s3NxUz8BxKGgrwEcCQM8Oz3q+fdwgwaa5JSB6MF5JMBYLy3ruGh2SLADKa8n9NX6MC1wbSZsxhomBC1yCsywSug263EXVy3Ll9R9cMAIpMJf6VuIpEb+rxI/09ZITxW3di357ROHTogKXUpMsOKcSAJoUbNKWR18AOU4TQvCNEo9VxYKalwMitatN3xwTPDfJGxQScvdbEnHPlmAAJIwBVDy7ER7/z1jtJ8NhSRy1scsCkatG3vfHaqJiSslsF3BWzEB9w8NChGN09Gh9//HHj88v3thYqar8293kVM+nG6ZY9q8I9X5c8Z3UIFnHD7Hn8kDXo+Vt1ktA1mNI52AYSV5Jy/IoKLuoAgcCDj3AsI81vCjNiS3uugMgxKS8myQb+t70tm7u6vqZni/3G75CZV6Gi7EMRV1g3+2c/K0kJbiMB6E5ndW2sr0bn1mZcODUWI70dsXuwN/bvHpat431+/buP4uyrr8fy+mbMLqzElrobu+SHZiTXRTGgO7q6++LuvYcxNDpqqc6FhRi//SDOXzirvcNepVCBNNOp0ydjZWU9Jqcm4vXXX5PEz6efXotvvveWCg1oxP/5n78f1z7/IiYeTsV//I9/Hb/61W+1Z7/9J+/FlU+vxOOpibh06ZI6hn/+y99I2u3yG5fjww8/9owk6WZ36JmwPisryLJ6fhegJ+/FGmMH1IG4vKQCC7Nf+B3ATc1ko6iZ881ev/S6pKE4+6w/e7Ts2oF9e939cc3gp+z3GsCyAcjz585pD1y7ei1JDQyYNrkDIASw9Ef//cf6N/fCNTx+/ERxkc6EunJyVh0gVcsMsmYXggEbXsSEvd2dMTjYr711+vQpFyCmHkmOU2BSFij0V5JcNZu6CFR0dQAoF9mNPVREI9ZSNrSvT6xZ3lNnhrZI/GlbCLSE+MQexT/SUUOewXsg/8lZIN84sB9y2aL2pPx3dmdTGJVWuXIRS+9hT32GKGbCtDYQVZ0Vsj9ipZstyzktgLJ8rmVdnUt7plqCdSmHWflz2Xl13qYklItCa4rGXUwpBQLitX7NOJQdZF5YR4dmBHV2wRDvcsexYhN3iItRLHk4Oo57tefGxg4r97x+40YsKbeqDhITk8iReD50yHBddDjwDMhVKwfa6ZdNMhp2Dppr3OpqW/12fV32swhgyjlhmufz1Rwe9iUyrOkv62+EU2RMJIKk5pkgmwWWAH4BGciyjOT1PG+APn4Gkx9sgK4nziXd/pY/zo6D7AbjDPP3ne0R777zaty6fj2OHjqkmU3o5v/jz34aR44fFZkRzODY0eM6B48fPY6+/l0qDt6+e0f77t1331WhYm5mNt558+sx8eBhrHM2urvjPlJsDIBWkQzdewOiyB10daJ8sBjdXW0xMjgYb7zxtThwYCxuXL8RVz7/XIWKJboi6HCQUsVgbGHvkXHt6orFZfa8wX7Y4crflJtCJOL9XWQvkJz9VsQoyc+25KgiaqXEnM5/4gp8LcKi5pMyuJ25ju0qJmhwvRjqng/XJ1lbFya7IYNmQQ2shzxAxfHVVZ1JEfey0M8Z3NR7tMUuFVXdFVlxNMRH4hrH8i50qPBP/Mz329tEhHV81S35WoqX6qBJKewMkRs5z85YszX2LXxE33suT8+ML0NP5ZZJoKiKrQsXRTI0MF7EBXeDOEeoV0st8Q/GzHW9iuXz/Ss/az1jrefyuXA4OxsaRQcVsCxzW68vheyJ89fnVIzaxC+exznK1lROWL9fNkv7Kgmb0POIRckreWnuSEqKVZGA58x+Yt9iD/C5/IziPnQY/LRmQ1DUl4+z72rk/ImJcP3koMbErL7grl0XixzjpU2XbCj70ViUB2x7xqift9/fhBvPCUO5AQyqnrWUQiiwdJGrW7Ic2Vh1sq0sx+HDY+qmwG8PjQzrLKFIwn8hB01NTIkMQZ6+e99eSb5y32BtX3VUvGyHf/X9P9oV6JudV1BiIM6gXasDIvCkGl0SJmbmryvhLM23SswNHsPEaVZIJQEgIBkArMcB/ZJbgklqSUJJRGZnZyTRRIcAjp6ggtZLAGWKDFevXRdz5/LlS0pGrn/xhUB3guHOni7rfHZ1hVpkBwf1HiQEBORnz57RMEUYfczBQD7q/sMHAvLUxoxMALqVBC+Pn4iZdeHiOQUYSH+wLrw3ACvGCeNJMA5Yd/zYcbUmF3hN6k33CGu0CViajGgGMdJ1UJJBOFw6Ieq9ARcOHz2spAGQ1TM+ABEX48njx57pkMB3tedhuIdHLNNCsipAX4w9MyIUlEjSCeO5FQMwjJ89072Q5LUWKtjACvwSwCrGTGnrqRKdle8Kxvmv2WAO5l3non2aAWRrceb06QbjcWJywtfV1RPzi4sqMJGkWFbHrcf12TVoqAZls8/Yh4DCjFQ028hMtAqYCFQJplk3sSYyWAbIhZXNwhCQdnR0i221e/deDblGykssHjnclG9hH2dlvdjr9scuVhAAcw0EVWIfaFBZm/ZlzrzV7wFClQzVTgMhtm3x5JNZWQGMf/d5EM+BSxP0aH2/Al2LGdMIFtq23TadgL2AIEB3mL8VYLUUKmBc7QQiCxAuFqgDx9SabGVXZ2eDrjzlZngOPKMCxFgntZUDXqtNpAlWVjGO4EBDnrdcYCRQ4n0IPLgPOljM+mkOCXUg6IQQqYlGUJLFLbHZUpqninzVmg5oBDBTwbr2UBfFJzQkreuqs1Bxo/TXbb/4XFgPgJCrKwA6LcF7sbaTNVfnCQDcLKMNdXAgI8HnFAsYiTi04QEfnEyYBY2sBOvhgVwAXAauHSD64jQbBzuuGSADOuNKwFIvvVj4YizFdiwsLEd/H0NZ3RnH/UiObdnzEQCK+DyuA/sIm4mEkc/AD0xOTgXyI5JqodiqjhtYUO2NjgrJwGXg7NagFpZKMp0NjFtCUMm9khLPieAUUGxQB03O8ylGrwFmvwoYLkZiPRv+tjWpqH3fKK7VcEwNsXRBgM8B7CBg1VDT1M9VkaPkWZL9VJI7tX9U9IWxNzpqacMMihtFkOrKyuyjUSDOeUD4jBEkr5aWxe4rlpc6UtosO0H7cSUi3FuBPPwX6TTuEVC49qiedyY+LlS4K9JgkYsuDHWV/8/AvMGoa/xdDQJ9cXGhmaA8b+l2FioaSUJLx+ZO2/iyokf93otAj1a71fz580O7v2RV0/7YftJlQkfFVpzcvyu+/c7rMT83G9NzS3H38Vw8eIKUWSgG6OjqjmeLy7G0SnJi4JkkGJYmWvoU8Lyft9UhhZ+F+crmxx/jp2umBPENNtLzEwy2NzpbNrckh8lppZABII8tM4FjQP6Qv9HsmyEX1vgaJiNJTRWH6rwIaOCCtwCkKVRgx9yt2tHp/cDZpQsSNppmrLS3x6lTp0SeAIhCNnFjeyuezFjfm+sHUOG66O4Qy0sdHCltkEVKPgsgWYztdUtNemvVfjLITneHmNf9g/qvz7617suG6qxnQcQddvaNik+y+Meavvrqa40ixC2Gn66sKi6R/JPiBKQyLedVQxBli2RX3SGGr8GGAu5VoaLsae3HYvmWneOaGkXCdByO88yU1QB7yAQ5VFedxRmr4WrYA0qA0WZnnSg+wITt6RYrlI4FkR/y2vAL7Kd79+/HkcNjsj3FtBYRJuOnmadz0d3TqRltPDOeB7Ev87i4TDp0iak1/6DPs6NYM3wPS4zPxa9glwHwquhWsnisuTq+1KGDxCT32CZGcvf2epwY2xcHR/ujr2M7DoyOCFyceDgRE4+fxqHjp2JqZjamZxfi6fxSHM95dR9/9LG0zQ8d3I9jiGtfjKtoNDKyS/Hb1NRkvPHGmwIriCc5izfH78WJ40di/4GD+veNG9fj6++8HZ98/GGsrG7F5csX4pe//CCOHjkQb7xxKf7mb/4hLl48F0eOHJG0F7bzP/zPfx2//+1HcevGF/G//G//a3z80Wfx0ccfxb/79/8upmfcuSGt9PWtBuuR54ic1c2bN4K11jPsYAbRdnS2t6nI97U334x/+tnPXMjfhGhgqRPOGWfpja+9ET/92U/1vNnV6rxIQI4i9MnjxzVIs2Iqnh/ycpqLBKMZyQnm3SHPGCaOcW45R/ijz699rr1OHITsE+fx5vgt+VvNzEhQr4rzAs04UykJWl2q1RXC0PauTp9HNPa/+d7XBaZ4TpcZ8ZxdgBr+y32tbazJhpGbkZfhL9lglQsRU0HicAfhhmYPTj6aUjcX7w1fYGZ6xgUOzeQB8PFwea5V3SbMUJlfVBxOp8royB7F6nwtvfskLSCbxO9SDqI4Rhwpjf20la0FuCL3KJ5IoLa6Dx3nUHxyB0VJVZZUo8+3Zy04Z2K+CRK1jt3cYefBrIqfJfuFhC5FFBdURQLLwhPAFl9DaAMAozOct+rr79X+5bkA3o6MDgvMolOZnBU5PIowl16/FB998kncffAw7aoLUIpDu9Bd7xaIi2+kWEZhE1vS2vXd6rerUGEFBMfn2MFWAHOn326Ny/h7+ak2SDzMT0q5XeKU7KhwMTZEANMrGcrEqVV8wv8R9/IzzgZnC4Yy50syoMgA9vVpD5DrKy/WPBfLuVIY4z7ppCIGpGuF3O5b37gcD+7eidWlpbj8+mvae2NHDsXCylL88te/EjHk9KkzKgAtLSwFMmRIbt17eF+xFdJPt27cjGczz+L9b38nrn52NRZX16JvcDAWGOC9HepkUkdFm6Vq557iwykWMMFnK/rpxmrriMOHDsd7778fP/vJT+P6rVvRTbfNVnbZra5FN13XW+4Kn52bFW7AHB3wBBZYOU8OO8cX8lnVaV6F1oorWWZ1cSdZip2vPZhSukX8EUks/S92HdKp5XNXJCHW6ABWVx92wRKT7G06Kfia58B18AzAQzjH+KKKEjY1GJmB2B0qKtV1UbwrYiA+oDFjgnk2m3SR04W3oUIQc0CZR8T+eDJt2Uz2tLtiXTDQrL0XvCqOqriqtYijprFiA+Xf1r8rr/f+d/eKCvk5w9Hfd3xd9rURryv6+xIc0ChYvDjuTSA+Y/eKm+rzmrlAU0FB5GTlNxQ3W+ZPZhdBHrg6dvpv87Of79qs7zdrLUXObBxbr1UWwmupqziArZMaQxadIBfjwzhjnFEpprS3SSJexIrVVUmAsVfwedhWfg65boNCvrpSTZwgTqUAWvKqxBTkli5OI58OMdJ4Ii9smG1yU2XGkoOeMcGa8rsQcU0Msv/lLJBDm7mJTzJhufVcDSFNiq2KiH379wvfRIYK+9ORQ8G5Z/DKixcu6jwz7xT8BOl7SArEhuQbPQN9WgvFC19JP73w/H71zT/iFTjVlxI5WUV0O5QHmzlgcoKoZERN4DmgsWUuRTHbi+UDsExCyIuDg+GCocxLrftr1ooXu6u9QxqbHZ3tKlLAUiGBxPjw2QBnDkiss05yAGAA6E9xQIMEt7fkiJEbwlE9m5uN3u4eJZq0fQ6PjrjdPtvlYTDBJsYwafg0oFgGzgXkCxTa3FLlXay9rLDOP3sWJ44dVws514MGIkUb3o97g2ExfmtcwCpGtcB3DWfNQWQ44qNHjmggDkUYXgB/OHccNtfJQE7kBjCAAjGSnQxgKEAv2mJg0FJR1SqugW20MWc7OSyt0j9V0tLTHXPzBu4KpFCnJfI6ArPtuCQVktdaRYPa4mJvNoYl+fcx2jVctlg+OIvDh8Ysv7FtPXuY4gODu2J2bt7JQVa5tU9Sr531EsMpAQj2Eq9iRROIiy0kXd+eBniB8RYDi+CcwdXJKIal0dfrlnYC3c6ObiWZGP3p6acpDePinFgb0q/MzocWpm15aGk1twM2uUOI62DdYZPyHjBclXC0sCFfGPTUoKYMQp6XwnhBZCIg5su67voesly5bhU4uv3Wz9/MaeYmuIIvvDgTUMFEWaywdFczMFQwwt5EJgjtXthmyQzzFboTQAl1y9At/i1ZK5hrNWgtWZfSn23MWrAtqS4u9g5JFee2gF3OQ4M9UQEgrJhGh4MDP82YEOPdsxLE1kyAnuvnvgAzvL8t+8HXAHqlQemBgkg19OsZAgaWzAgfLcYETAgKLikxxmcXYGiNZw+k1PokqN1aHALsV5GWobDJHMJOsE/RhUc6bHJqMuZmZw2cU9QR8OcutZLeo1hmgAtgrbR5PfwdoJJ9ukIhJCUT1K6dElqNwFiBfOqPCgSHebhPA+sowhKwFfhmtlSvZCOezT/TPSN/150DIKv7SCBcSZTkGlgv2KycYu7KhmRBG7Ysa1QBpgdjbwlMJTHBvgHESdIp28TLBpFE8z7shwoe65xwvQxape3cwKg7cfTz2kuao2Gbho0XAzm7OVj3haXFLHpaN7d0WZuFldKatf6/WJldXQILAXqrk8JJiIvHre3OrIsKnpkMbqyuKWhdzdkcNROgilKAlOocUXdPcwguf09ix+fyGTUfw8m/C1OysxQZxZatod4ULrtc5M7EAICdWUO8f2tS8yL7U7atNWFqtXet4IRNTVOu7mVh0x8qVLyoSFHvWXu1mUA2WWn1WWXv9N8sFlWhgsCinRkVB4bjzYsnVahA+un25IyGaXMWJV+4ayiezi/Gs8WVGBzwrBc0ZgEi0f/mDOBriVnQR8dPAB7xedhDF0vNcqXAIf3slGEpX8ge5H+cR/avwTEPtmfzsm/MHKMbwrKUPGOkPUh0mJNVe67WvQpa3CexBkkR+wvbg19YW/Ee4JoosPBZ6jSQvTRgJoCysz2W11b0M4DzmelpFTEpzHvAsoF4xRGZjONWJiamfA/Sq6fLkSTPUnXV/aHuWg3pxd4AjrljrRjNigWye1QdXJlIivUMAzplWoghkZa0H8iZF5IrzCSY99lYt8yRul94lsw/S/lMdSVaix/QlUGFe/bujU8++eS5LuJ6Xg2greYJ5fmpc1qxNKAXv8v9iLmYrE8XOB3rMIeA4gDdxop5NzY1eBr/s7i0oPUDdMKHE/9ylomTiWfx097/7mLDz1Dcx5Zj1/v7e7OLkER6PfpSCpHOn/ob5EKwSYvLqeevNcNGuyhkYA9pM8cKtqv+WgA5IV+ObsBW9VLw31iOM0cOxNieoejaXo+B3q7Yu3u3zsWVz2/Frj0Hoq27PyYfz8T03GIcGDsgksvjqSmB+QDbzDSZmHwUwyOj0duHdvWmiDzMXHAHWMT9hw/t/zq7dC3vvvfN+OHf/l28cuak5J5+9KN/jLff/pqe87VrN+L8+dP6vQ8++CBOnDgVJ08ej//rv/4wLpw7EyeOHo6f/OSfYuzwobh86VL8/T/8JN5481JMTj6Ka198IUAMMm6jG6ujPb7+zltx7drnAhJ4IT/iroI2EZxee/Vi/PwXv8yzabCNfSBpv66uOHHyZDx4+ED3wzln3bk+7R8kI9VB6bls7GvpwKcsE3tVsovLsIW39TNADJ4bn01sceXKVcVB/B7gOMxN/BS2CjvAdSB52PCv6R8NxG03SCTEPeR4nLkOhvUK6FkVq/u111/VEGjJdbW7kwhSGPeDrWOfYyfoVMGPavA187/ITySN6xl6nBGIAhrk3dmp2EwMWljaxJY5nBsw0t2AJglQLOCMAGRx75q10tEVQyNm1ptYRzcsRBDHyKK+ChA3uN4KKFU3F9+r4r9lbwxocm2sjeK/JE+I1Z1gXNnA8l2SYEv5OsuS2saK5Jd5SH2OwH5mkEFeS0IL14+91Vy0LHxAzuO5Ppl+nAO3VxRPeTaPbSrxmtnuHbFv7/6YmX0ap10s9gAAIABJREFUN8bHLYWqeIz8okOxFtcq2yJikklDvE8jXtzhvLl/bFDdF+er1R+XD2r9s53xhHOZtgYxUuAx8S2xfXu77JfyQrfn6J5KNk0kHc2oRIrXXTL1/uT2fI2cJmcRW0JxA5KazlI/pLlnjVmLEJEoVEh5YHlJ9uudt1+Pu7duRtvWZrxy5oyIkm987VLsObAvni3Mx+9++9s4cfyk9vHkw8nYs3ePZllRPH469zT+9Nt/Gp989EmsLKzEd9//bnz4wYfR1tkd2+3t8eTp05jj3igirBMHex/QBTY6MhiDA72SoRzaNRDDu4a1r48ePR7PFhfjwcRUdDNnUYPO22J1eTW2NzY9AyqJo5ozmcAvcb1iTfZy4gB81ujuEcUDvFg/SXCv05HN0GF3QEopQIV9x+slCyyCnIqEjjJV5Gu3hCSxvWSYIAggGad5gHTp5CyWNrAcz9gi1+O5GPxtT1nc7JRoFAIs6ek5VvaN7P0i3ajrKeWUFScsm6ToPJZYx3JGA7vAvVwkkT2oeQuppvCy2LQ1Ji7fV2f++b2tn/qDGwWJKiC4ozl/qHuvIkIVCZrFjSxlVk65o6Wh9QxVDM65qHxcz6VBvnDsUXHhzji75v6VdBXPoHAd31vmtZk8Nburnv/Ziws23hdfflXHheVCsf0lyVnzsvgbzixYGXuqFDzYL4q1c64EBYg2pMW4Ac10tA2WnHPaVs8cNTbAbvV6592l6kUjlgO3bHQ3U4Cmi91kYD6TPUicSS5uu+eqBDgLT00+hKKGOmSsFlDxIvutMAgKKsi8E7PzdyYZbEkphq7jknrfvWe3YlSUWtizszNPlY8scw19/ZJ+lv/6qlDxsuP71ff/WFfgcLuTozLAxd6o+ymDV8aOA8fvqPrZ1S2HVoZR/0VeaBEtyzUZfzkBkupsH1NL7HabWF0koNgUtC8JJgjICMAIkIqJDuuGfz9+PC1gjtZpBlcRcJPPOnFv1/A/hj4+m3PV1e2yg5KSohoLo4fgnBeDstFYnp8nmWiLHg2nptK+V86U4BhWIYE0syw0fDoZZdzjwb375H9ouSXhh3lx/cZNfY3u7Z27dyzzkgYMhgFGbXjXUExOTqjNi2SPjgoxkdbWYmRkKIaGzYhiHQg69u/bJ1Cwt4fW537JSlHAsERBuwBNEhECF4IH2B9KGlMihWFClXDIlXS0q3MBp652dBlPd1IQTAioTvYzfyeH1jKcudUpFhhk1gzBQ8kkwY62rjNJEMwedUsQkE1PK9mkAAQwA6hS4Ek5zZI5aIJNTRkqtaWLAdyughYBmNoEVZzhXt0dw7OU5E3OtNjepqreJ/b3nj37dY/Pni1YKgCNSrUDGvSTNmGJuCeVQeAzoHwCWzhLAdQkX+yzwQElEdUKKMmclGN5GYDn89YEnn0GW63ITubyC0C31uAldUbrHfT+KRugIIyKVEnE5DDMYnV8qVBRBZEsYADysp6AWeyHBugdlsoSG65lfkldg55tMc+VCLkIWnvLy2kmbbVNtg7+liPPgFfFBUBwMd9ymKMKcbYtbgVOXU0FKm7j5yMIkhWo5iwCzgz3AaNtdn5O4QU/k21Tka9PSbE6QhiQx1ydZNmpaLnlORQank2CgxRc3jSJI+tJ4CKZDJ0vJ1S8VDQRm9VMPmmwbm1pf546dVK25tHUlNjJCvhhvYttT0HMLa4ejO1ETZ1T6jrxeSZRV7ebChzNZI1n5DX2AHAB9zkY0p/DHrGWMusuxlRKDnH/gJ+AJLoO2rw7c0B1Mp7EuqRtVnKBjtlqTVzA5m+bbb3lb0rf0zIFHljNizUB+G0Pt+xL8iSBANsqrxv7h3UBzOL8YxuwN6wzTBSCORXCGgPZzV4Wmye7XqqIUtJRFBnpruNVHRlKfjKB4u9VbJOtdJKhghGBKQBLZ7d8AjaufKPBvGR957m1PbXPxMJI/mZtXa29JJSWkGM4uANrAVOsUWrHlvQTn1+MOArirLc0UaswUqBJzW3g9tPOcymAYfhPJUs1/Dy1/P81hYoXFSla7dPLYqb/L0WPne/dmqTxvk6K/gWFiryY7raIY3sG4tXTh2NlaSFWNtvj1sMn8WR+WTQNzvrg0FDMLSyrq6Kry/Jy+HPiBcUYkhFxlwHgCfuruh6RHagBrsQ1zMUCRKbLr4oP3JsIHevrmvcFQ5IkTVJ1GVPRHci/6RzF/0hCpbc3Dh0e02dRgK2kKAO8xr8B64m9ALbVQQTRQJr5TrLoHNg9MqqOKfYHUmSPHjEceCsOj42pUIsuN/MrDh48FJMPJ3RWdw0OOFZq816Xv+R8IMXR3hXjt243WLtdHUjIZYdJAiAQV6p138Ob3b1bDOgCx7kO9jh7nq9dXHAxVMm1JEW34tixYwLPOPtogiP3CYkBW1ZrUprsfI895IKnYwnstzpgczYa6/LZlSspA9AE6QtUrETcYKPnBhmAcAxj6VMTQiQxo269TP7lg5jBoEhA/y+pphwki10lrtDshmGzCC230SG2O/GtpApS4kNdeDnLS8lzdqFSZDJ24vij2MoCKRmSStKv5H1bNsEMas+oKPC2VaanYsI6f3RFU+hAG38V2UQkGCCWbK3GodHBODg6qM4KGMKAWcRft+9NxIGjp+Lp/HIsUHjbCmnnSyYx2Ys8F+L+Z/OL0dHJIFgN3xKRB2AV4B6QkG7omdlnsW//3pieno13vv622JY3b1yPP/nWe3H//j3Nbzlx4rie7e9+9zvJsgDu/+rXv48/++6fyG5/9NHV+PPvvCd29q9/+0m8/51vqpiLhMri4opnVMif4d8pEqJ93xWvnD0rcNID3Sls9mqfEj9gmx3T00ncKX9p3+tuRshXFMOKyY6tN6t4U8QA/D4se4hLPBcA+RquzfvTwUxcf/PmLcXgyrVUGIs4dfJ4nH3llfjZT/9JncXYKa5j1+Cu7DR2LAegie3i/dh/YieXrJekaEzSkSyn9h+govcHxQN3V3fGpUuvipCGH2KvU7go4LcKdS6wtsfY4YOyX9xrxdAQMwYGAPFTIrGLbowVAfrYmsePHjXiHXUxlHSS8qcOac+TDzEIHZtmpmyv/pYCRcV7slWyUxnXNAaFmzjRmg+1gn8645nzVKxn+wPBr4p3SQ7QGbccDbapwH7WRTkyw+0zjrJUrDXSC1DjHLtY7PgXoIq9Qiy4Z/ce7asrV67EyeMn5EtQDqCLgK4ork3zDVNXlthQ8zognvT1xsSjKRX/NAsDyrqGTe/SZ6tQYUMpELkKYC/y29g5zmt1Vykvz1ezQNPMaQqYbQVO3bHapkI4EZGKOLwPs4gyfiYeo/Og4ktya9lVSGp0JqRf0LlJYgtdzOxb9iL5AvfHv+3f2lRUoLCIn3Fnt4su5Rupt1+6dCGmHtyPrbU1zam4R3fF2kqcu3heXY9iNXf3xMcffKQZFqO79yhOwOc8nZuVjfnsk89idWkl3v/T9+Ozz65G4ANjW4WKew8fRlvmxuurHiwN0ezQwX3R3r4V22jQd3er07Ft2wSAxeXVeDT9OJbXN6KHtef8BuO0PUxbVkmkqBXNeent7Y+nM46lFW9vuINHHYsQFZBZ6+83oStVgLVvkmSjx5n7qMB51krFAdmJRnTnOQWKl1A66M1irUl9nGOKiyMjwyqGk0/yt+x77CL7Uoz6nMHjjnpLASfu35jHsrBoqa+hwQEx0nlhDygwEQNoXgwylEicK94wxtE/iJwkdq7ZBSUf5oD+haFp7ePKXRr7+iWBbGvsXB0TjThVxRpjF47T7Hst7epv1hkROU2F1C9/UGsRYud1VZ5dHZ6K71q6nFrvR5+XHQS2YcZE3Pzh2V9+NS9iZ5xev/McjtHyD5Mgm8WO1oIG8VYRzSr+4tMOjR1uxGs8N/YmBDbNlgVfW6M7b0j2UsXzrY1Gx5oIAgLTthKDsgy6uj0zjjZhk6K7iRdFLOHanI/WlsC+9atQIXwtu2PtR/gd7yv2r4g3Is7QLbmGwKivAeIPmIbOkYmMnGniCiRUIQzMzc2qM5LclZ/jI8AAtVfJB/btkx9lliHERojTT2ZmNKuLz8IGflWoeMmB/Orbf7wrcBCAhKQyD3Dpw4nBl5anEkOx8lOrk59TABBY1klQiYaombgF/BTYDPCDrIwTHQe+vKQZ2hYKSDE8e/aMOpB/Nh8PHtwXo/nVVy9qpgCSChx8tJl7+/vj88+vKcgjQFCg2BZxYO8+BX0Mf1xehGnmgXRHDh8Rm5/2WAIQChVIP9nJbqgTg86KAwcPqh0U8PHwkTEZEGmcZ+stfyvGBp+37uCXgJBWZYwMgQnyVjhKEudF2EBio6+oEkwyxfsBYPDC0AwO9Ou/DHsmsCxHKrZiX78YTNJ03NqWU78zTqt0V0w9ehQ3bt6SXBaBCGs9NTmpv5FjMbe86QxTzkhst+1tJzmZkBfw11qoKJaQWPECoV2dLufU6kz5XRt5sxoJaNkntGpzX7wHDxpD/ejJTOzdu9/JTjKha+YBAUwxSZUgJCu/AiU+k6qx2Z1N7Ud09rWGtFSLUUGCZ+axgd02MY3RLt63l2Gjc0qQWSE6Y8TO76jBd+jqe/CzWzQrYPB5MBOyNOcBwQ0eW+rCYCPvTeHNUl8eoPmiVxUrsh7wLypU7AyaCuRqtComoN86E6P2BdfSCDKS7aGiRXYAJM7ckHiSX93yQEExabLtUQBItea2BHduF2/qNFb7u4dDWzJJz1eMezOBBZAg59QDQxkGXM6XyE6NAkQMCpmRpgH0mYx5zkqX474M/gjIKaZWMF52TEUsQBI02mXPPB+gwZZD3zUTRsmFSNO4w8wIgpGupm64igx9DGlDGzOZdTlQu9aJ9wJA4MIpJHDfgBE6d8mMHx0ZVXAiYLytLeaezTY6Drh3M2y9J0uCDJYJn80+A3TUEMKS+VGCYR1pFTYVDFOI49z7bGnAnoC55gwOXWd2xFRwrWLTJjJngOYeUCcJNAo4zEHZMKBn/XIzDFk3M4kI+Pz++jq1uNVOq2DcZ6Yp40Yxy0AkLFA6hZi9QQIufdnsPOAaq0iqQfWwyxlOSAdfHjakeOh0K1DeoBCzUZzwiGWTslOsMSAUvqAKFawlMypKmoV1b6eLRQmTwVheVWxSoULP2DMqpImcBd9i0cv/1cwQ6eNbcgJQSAWIrS1JHlIsd+eEW9HRbVYwrz1oxk4Bo1x7Mc75XGwo+4j9rGJGSr/xbIrF7WKHn091VAiIEbAFi/H5zofaVzsLBGXXvpy0fDmraiReLZ0aL7OLrd/fWYRovYZKvvQcMmaphO2fK1R4PoHtu178e3s7jo72xpsXTsb66lIsrm3HF3enYnrB80JGhoeiE8Zve3dEJ+caRrftjv2qh9wWcMOQWxVFV5blF/E5JBQliUdbO9eNPm1z8HNz7SFP8CwmHj508QMG1fJyHD9xXM8fULR02iF5QADhGijKV5GsgLE6B5wV2yyAQZI2x0naL+ubAnnHDh6KW7duSf/96OEx7Sc+f9+evUq8Hs08FniAX300NR0H9u/WWgKaues1QTmtyWp0tHWqqGI9X9up9jYnxNV9i0HAFnPeTGKwHaiBu617kJ9VrGR/YuaZ5D7W1iSj8+677ylx5MI++ugjxZBcI/5ZEhcqhLu4jV3h5eIfvt7FLs6cZHUGB6UVfOXq1QZrt/xoo9DZ0mHgzkYDELy3pFy6AZq7dZaxFWKjA1ir84Su2pQ1pLtZLOtOgXTS607NbWaPWDbSwylhz8JIJXlnnyE5xH5srk0m2u1tSuiJnzzDo9fzkbYj8D10xfDaNTSsvSoJsfR97Nnyv/UMWv1x6/cc42f3tRjo3MN6EAWdP3kgDu4ejN27egmclKTjG3/5mytx5uJFdSmtbETMEj8pnuuO2+M3tZeIJZeX1+LW+B3F22++dVkSSPfuTsbpk0dVgJJU6/R0zC+sxDtffyuYawdgdfmNN2Jm+lE8uH9PMyeQUUNy6K/+6vvxu999pELG97//F/GPP/25pPPe/cY78bc//GEM9PbEK+fOyf9cvXot3vvmN5V7fPTRJ+rU62JuRmePuqnko2EFD/TLP+O7FIeuIrnS6zlyOV+OeJ2vyV1MVKIouSYAAqLT559/YfZ6xdua/dcRY4fGZH8++fSKfIBi8i1kSjHb2/Haa6/Kv1/7/Lr2lIgh25beOn3mtCTc/u5v/045AtfH705MTqmT3UBwW6whZ6VZMQb2eA/tv2SpYylxewA1ZvOjOb8mglnNviOuYn9fvny5MW+Q38HPQOYij2G9KATwmZxF5tnhL5kbgE2R5Fh7u5imFHGxeXR5eaYfnfYD8fQp3bBVVIQdzWd0S8oOlqtJXF736rSis0JxwdysfDRzRWQXMy6VXYDNvrysAlLNpXIMnLr36hK3y3CXkbsSC+gTiSQ7ynw2/Huan5NduSU96YKWcwq/DA7KZosk5llUFKGlANDVpTkVyOnwwi5/5zt/qv1y7+69OHrkqIhy2FwY+I6lNnRtmkOk2LZHNpVu2IXlhbh583a0tRNXMoiYodCD+po1KKDXRIiVl7Ci3eFn0M5xiYqouably3fGDjtzSX4Pe0zOW1Jk2IiudufQ/D22FPuk/ZEdwnxeESZF/qFIKyC4lBB6orOrw7meZmEOagYZ3VzknBAAkWu2XKcJAaWNj03p6++Jd95+I+7dvhVLz+bjzMkT8WhiIuYXnsXX3n4zHj1+FOfPn4td/YNx8/rNuDM+Hnv37Iv+XYPx+fXPo6unR/LTX3z+RawursRf/MX34oMPP4y1ja3op5gxNRX3Hj4g6tZ8Cs5sbPMs3EWxdy9zMDuEJ9DpgV+gqLSwtCTC5VZ76DOw08SRbZvbyv0piku+b3Ul+gYs+6ScXyQfCv1WJxC+oGyK4lCvchP8qF4iLxg81yyi7ZJWQyXD3d7KKeQrLU0qcoKjy0ZOS1eInqXkRjfUMUxBmxdFxeqGpIjW2cZ1WOYQMJoX556OD4ZvE7nK/nR1qXDtPNL5In6a58gzpGMVJQfirWLPs25Ez8PDuwROo65B14jOacZwdTZ3xqatmEdrTKqvi53lJfNJzmTUUslJjKoENcmAepYZD6tjKuWLFM+qOJGyrS1d0RV3tMYfrXhAa/FvZ9xeOUPrvTXuKwfSK+7IWVrC/ESMa7mx/PJ5YuXO1Spz1iQL1R6rvLDWyMQOk5orJ4G0ge1B2g47AmEZW4nkn+SJl4i7e+SfpKIhn7Gis8DzZk9jplWYlWqA4zwKBVInkayzfSQ4gSXPXADlfNR+KKUOzg3Xp8JvzgPU3EuKcOAQ2YElieo2k1SU4xJfZrFMqg7ILq6s6PqIw4jBwAXxc8Qu2Lel5cU4/crZuDU+LlyV6yNG4AwQtxOD37x1UzL3fI1iDPE+78V8yK8KFS/Zi199+493BUZXzBopyRezvFwdtG3yoeV/Oujra3JmsPiqRZTDSAKGHiJsFQJWJcEwaXF4acdVGFALq4Nb/g5WHuxc3vvokbEYGR2JyYlJ/T1AHAkniQJBKMGDJKG63OKsgUnJZmxnCA2ti9vbCo6X1BXRJ+d4aOyQmFcqaMSWWAOTDJ1RYrwhY0WgzeAahmdzr7RJI/sECwNjwX2gP8lAvBPHTmhoDUEBbAwVTJaWpEW5a2go7t27q0ASI0eBhgQVBwpLlyQZQ3jh/AU5VBJHwDExnbfcVsZAuHkSITEdkB6AbeS5IMXGpBugd2BA4OYDgRVDYrGRXPD+BGAEpGJc5TBnsYI7rcXngNKSOQ0d/nLULYzfMtqt+6DAN9ZTibjYLA6iCTh4duwR9CClnZ1tuICcDLAmJFIQmYwHHJ4KDMglZdBuOSmYRW4V5WduC5V7kwPn2UqjNoeHUYnmOgnm2F/W5KTzwe2uBEH8Kck+bPquzl4VTEruxYAsyRP7KrVh0xvzHF2wyYFN7ST7MM1hr1sCjPskKHGLsa/RMyxe9Crd+CoL8DxaQLMd9AkHE02mRb1jK+PLLC8HN2rjF1Dg4YFmojjo9ID1fK/UEncxyAP/CoRwQdEyEnzPDCMz3DwA1UlVq33gZyUXVnakVac36WYNppoCAp1jD3Uv2TgNiK65F9lOX4w2WDClk4rjJqHie2glK9xOEF73KOIl7EwSVxjEza4hPq+7y89HCXgCl8WItv2zpADJfLW+s0aAJdgiAvoChNmfmqPCWkr2YVNnmzNKEbdYWtiKkmvjugGWPCh5XY/YQ7xrkJ3BLop6laiJbQtzMQsdCogEeLvrhFbt1dV1JysC7n3WquW6ihaOrT3noZ4vv4sPKJ3WOv+9mmWBrjLnxR0oYgDTpdPbI2mFYgayX2CtCrzJQc3qbqFwom4OM54NEjuI93u5W6UK53TPkRjBJm8UsnKYdp0vCopmKFv733vPRTc61wAzBBzoHLgLsFpwq1ghBnYWLbDZrCeFRi4QP6NOkbRh9axVKMiikXVlU/pJRYMe+SoS4UoUZNuSrd1qS+1XPbNEvheG3+7d8mGsZ6NQoWftghHoVGnZ1hkjueDMFwBV0nfuaPQMHknm8Rk6FD7/PG8Nvlc7tAFJp5jNLsuKA/w8k2q3w6RVcaASplZQYmcs4QTly90O9ZY7f/bPFSqqSM7fl33yGn/5c+Q+GpVhf2KjxgoAFxFHRvvim29eiOXF+ZiZX2l0VGxtt4lMARtwq71LTMa2ti2dVZIJfB4dj5IUyAG6AI/4YVhR7GMXVgyscK2wmwEAPEy7JHtsU7nv3aMjsjGAdSKFpD/BHvEZ7BPiGb4GvKPQS9JCoatANq1Pvh9fQ8rQvJtkbNeAZAMMbYpV2EcMg2dtuEZmCZCgUVghuX/89InOMIUJEkHZnwSrZM1FNW8On19f21TnpxmaZXF9Vms/VLGh0U2hmTSWLWKtVPAtbW1sL5IyqYVOki+2HEWStPd01FbngRl7kEtWxUyXFrMS423NnyBJpAiIZIb8Rw5ULf1qNN4ZVH716tWUnGgOH694qHUfeiAlMhlV1O5SwUP6x53tsUnxijlFxHUbG7GmYoTXApa6/EZ3T/T3dMZAV1eM9A1kRyrDm3tz5gl63T3xTPKhBvi4N3wd3as8S4A2d3J4gLYK0e3WLyeuxF8gkwrpxlJby9Lyhp1KZ5riY7oC1RHdnCNQNgHfW2e9MaMiz0MVfrc31qO7vS1eO3s4ujZXYnSwJ169eD6m6CJq74grX9yKg0dPx+pmxJXrt2LyybM4e/4VkVw+/fQz+cdLr1+M+YWluHbti9i9d0+88sqZuHnjVkxOTMWRwwdjdGR3rAi8bYvxO8zqOBSHjhyJJ9MzWou3vvZ6/ONP/ilGRgfjwvnz8etf/z5Onz4Re/fujt/85rfx3e++rzjiiy+uq1hx6sTx+OD3H8l/fv+vvhc//OHfy798/evvxN2796Kzp0egAcUTAxBI2jLXqUdnmT3IXiUPIMbEf3FWjh09poHs+H2B9Qkc8ugPHtwfp0+fjl//5tc6W5a+6ND8K/bhvr27JQV38+a49gj+p4pd+AMNyKYTRkB9j0AUgc4p1wKJDOkyniUgPddP9wjXrm4R4nF8sAofO4Ep+wyux2fCMph8ruQ5W0ho/Mxkpe64dPlSPJqc0rmT9EtKq1LgqHkOfq9tSWyxdsTaLpQAVO2Jffv2x4OJB8qJsHGzs0/jMHZofV1ApJFRE4Ukebm2Giura7G8tCIgn8JokSU62js1iJ04DRtQfrnp+1yQqLNc/k5rk/erImTK8OFTBeCWnGn6NYBbdTWlJFXF1NVlXHG2CnmAwHSMKq7zDDLfknPu8p/4AXXNdtmWLCEXlEXaM2fOSKng6tUruicKWvweBQveB3tfpDfkbvgAJP622rfi1q3b7lTKWA3mPV+ztjVAtoZpl3/dmdGIDZ8y0VWoqNjkRTEB33sZGZIz5O5phrX3qEhTMqFa6/Y2dQNxfQ0glk4TzSg0s7hIOn4GJeG3ID9Yczc1s0Kg9XA8nJiM0ZHhBvGRYhD5OR0R58+/EseOjcX4jevR19UVp44fi/GbN2NxcT7eePNrMT5+S2f54rnzcfjgWDy4d1/ktUdPHosQSQfia6+9FteuXIv5uYX43l9+L371699G78BgdPX1xfiduzG/uCCZuJ5u5i2QD3h+WE9vV3S003WeBXQKBSvrKrSAt8w9m4/u/t5Y1jO1FFxvp+e5cYZ5DwbtgqW4y85yNJJ9zBl3yiETw6nuLbG2s/O+EctpjpeJRYqHk5BhZQa6N5zLaa5EDRN2IOluifY22cCKoavA8WxhOQYH+mIDKTnyio6OmEeiCinBlOJVjIq/ZP5lSq5hxyimKx9tck30N1w/+0g5xeZWPJqeiXaIXO3gExsxSBFvcztWmbe66s4wcseab/GijL3Vv1fMorVpsOOa3QL+eZIEqj0F/5lfly2xtKMLw1XELEC/5OMU/ypZej6erXh8Z+xdmMDOwko9xxcVKyoic47pYi0xkHMW52r+nSYBqQZTv2itmrF8fpX34PepmRb+WdnGssWWAvVeRQaXc8ie0Tzajg4pYUAM3r93n4pwKBDwHjzL1Y1VScOR41DoUv7aiKs9X0X3lGQ4rkezKLODnBst7NLETBd3eZkQ12lsKZVk8HPsQ3wZOS5EH9aOmB97q064LRN3RCZNv8G/6TJ0PrAZZ06f0axL/oY9bvlNOjAcZ0Iy0cqB14ARTs8o7pYt6+mVlBlfay2/kn76Q1vyq5/9Ma7ACBp+CWIWK1MAdgI+bvNOfW+Yr90E3MMymjg+QHwMP4m45ygYBBWDJBkNainP9maCRg3TJZDrZLAuusIAQ4MC2HAwONEyvrC9CEgITBSAjYwIOKJtUyBx6tNJ+5l2MCVgC7G57kMMUE5VlsCUABaWDcHvxNSU2qxKs5jABCYrRhKngbFiPUj6MVZi6xCIRZvYP/ybogvGEwNEwM/97j9wQEUMFWI0+Aud6lGS91/0AAAgAElEQVStMQERnRBDg7vEiuG9WT8HEAyZMuuaAFusR1VuqQwbpCJx4R40CHJjXbMWGNgFGIdRRgtTWv3JnNbgc5xwarQr8RQQ3xxoS+BuINoGu8kodJBsw2gnWcGiA3WGCrvtsiS+NNRRSS/dEhtKYPbv32tnAagtzcgVBYV0wHA/BEYEn8VElRNNSaQ6T9yv2NMKJjzQ1Jqqm26FTeCJdeR5GJBnQLeTb+m6b22pzR2GNc+YBB42mmY2pAQO+s0UMBhWyzQyK8RYU14a2N2AnE5AAVFxNFw3QwnRsEZfd2JyUu137B2zxV8MyFWA7QpCOexiiTeD+DoHf8i2VGHAkjyd2k88awARSzU1n7kcWXZOOLlrgpYqPvB/qWPJzyqYNaOz2oDr99yS6gDIXTwNNmoGqkqkUi8Z4MKsXsd2GcM6ASwGd8nTwCrLeRkVKFRAwx8id8HekbZv2poCdeuZGgQ3FgZ4w7N17cULLqAgwSol2tnlUXqlOkt0C2VizjqS+GOvGkWDLLQokIHdwQDsZKQX0FxB19ihwzov2KDZmRk9Iw+MJ0m1zVQxSGvk4LQA7BoGXh0++rwsJouNoqCyKT1gEM5BkENDM0Vq/oNBbycULsB5r+rrfBYESSUnwllGXoQ1YH35PjadllOd75xxw+cRvKmQDIM/B8VWl00xrWrotgp5VQhHaiqBEN6HAFU622hd54BtaZFrj9Jl4qIT+4uiZYHsXCMBKc8KcLjW3x0XzYHxPEPtIT3jHGCbBSPAWv6OjgrPrrGUkIt1LuI7IfCeF6tSxVANZhLYRTC9E9wvaYQCQAw8M2DXknwFXtPSyyA4kr+m7JTnCdh2FLszWUEMjtvccIEl6ARhcKQLWjqfPqJZVPTXzq/cjSG5rJaCTJMB5u6Ahh3Idar7atixHcWH1kJFqw1s/f7LbNrLEinFHOyP9SyqNBJl2H6WCeJvbSc88BSgsYaslqlTgiVWOrzRLA4DzvF8t7fj8J7BuHzxbGysLcfss8W4O/E4phfMcB5ARqK7V4Wdx2J3DYiBCEsXmUm6BthnmhWzsuKYYpMuu8Wc/UXHoYFEnjUJCAVvpJUKiOff/MxdRUOKufh7mFclP1hdPD6/PrvsLRIWioT4IjaAZhelBAw2s5i6+E1LeJpNia21Ld2SJANauDwrkw48a6uRUNLpkIwx9qzAcNjSCW5rT/AbEhO35Bxx0Mz00+cK3UhPCIxLIIPftsydpcxsu7z3uEcPwDagqg4lipvIOmRHqWJKCgSaE2TmLACbCxRrskmtQKGAnM3NeOftdxSz3X9wX3EUYL1tigf0cg979+zR2sJ2b84G8nr6LPtMlq0RE6+7K3q6O6O7t9ta3QxB3NiIGWTdXjKw82VnAoBs90B/jGguFkzqBelrS25nbS1WVtlzPZbB6+oW69j232BDsbS59k4GOGc8WzbB3YyWcc2EQMWuihd0nwB+GjxpmVD2DnGwwMMs9Ov5dVSMATjVGV3tbbF7V0+cObo/Bru3YmP5WZw5eVzAKjJKH356LY6cPhPzS+vx+a07Mbu4Ghdfe1X7kqGz7P8LF17RPX9xfTxGdw/HqdMnYvrxE4EUANmcP7qXJh5MCMgi7qOzjeHUP/7xT+Ls2VMxPLQrfvvbD+O9996J6SfTcfv2nbh0+XXZDbozXjn7SowMD8ff/8OP4603L8XwroH4yU9+GW+++Zo6uX/0k5/H9773ZypUXL95S/YTYALbiW3hGV+4cCGuf3FDvtLdQ+5EJLYiPn711VfjH3/600axDJCMYhYxw969e+L06TPx2WefqkCHTy1ghTOBTyK+9mcxsNN2TrKjGR8Tk4r9LunTkDQEz4tCG9+Adc85WFhYkqwc+dSdu3ct8yRZX3K45iBRfKykQDJIrfmF7sgB7DTwuWtgQAQGyS8ixcvA45yFc/zYceUoxAXqhOpiuPaS1kskI3V8mn3Ns8Z3IZPr/LDbbO+UhmGfAuZAGuPvsYnTM08bMmgiK6Q/o2Cj2B77m7NcAJrwc+h9l8yP8iF1ZK42gErZlhz2KpIH/5dybvZn7kLjRezId0qbnGfVYOjmXEZsUnVtVVEDX0Vcim1qLXYWqcN5CXvLoJ2LOyawkGPxb65FHRnt7dq//PfmrRu6LvJbYijyYv6es0mxmftR3ooM0tAukfPu3auh2u2y/dg9uhaKMOb42R0WmQ5mDO0YgmtiTxTwprkXxQYvH9vyX8WkGYfzX/mB9N3qnk2WeTGYNe8RktgqLGYIaO6qrtla/D7+qzGTsSWHMQjpgg/nDUwAv8A8Kdaw5okB5rNveR4QF/n3/QcP4/Kli3Hk8H51NW6tr8fZ06fVnTU58TDefuct2RLUDF67cFG2mGJk/2B/XLnyWTyefiJbzLm//sV1kS7/4i+/H7/85W9jeHRPrG5sxvzispB29hCEH2w5RWuY1ciqic29vibZsi0K6dGumZyQJplt4WHyXZIIZdi29u3mlkgL7rS2pKvskEhq7jAqOWDhNtr/dI2auCXijyQZTXxTHEHXIoVtycNuOMdM8oTyAs2MqTzR+6JiP2wCPsKgsGXCNFNncTF9CPNolqK3h0IFMy1QRvDQbZ4RsQXPVlhMdmNjMyFOEYul02rkBbw/hQr2Et1mKqi3t8XCPDnMpgsVdE6trMVaAuOeUWPyq85jznerfVzxTyOGrYLiDuC9fHhroaIReyZQXzm2pH0pVORsrbIpJpA6rlNRsyUwkEpCfqNxbZlRO+LKrvvq9Mh8oWYp6Ww1YYc8z1Y2EFkq54ZxjbZjjsP4fz3FqlokluBLS4JT5hxF1KicrHHBOQe19W+chtimehbWhmwpuSWyoexNziJKKZzjoV1Dep7IMi6o2EjHsgvPdDk6h3T8TJyrfa1CuosIvJ/msuHniIGFlXRpXhHdEJwLEbyKjMmeoEtsfd0DurNQVlJ3loTyM9TsoszLwZsUb5IDp8wXhf0q4Oo+Uwb61MmTcePmDQ+U70V2vlekZuyRfp9ids6rwjbRfWhiLB3Jnl+EDeBavipUvCyK/ur7f7QrMLpiLUkMJJU5VcrFsrScD/8uuQ0OeA02dNXQ7VmwriguGJjrMENToEENLjRziPeU/AjzJAig1gD1NuSEYR3t27dHeo93b9/V4CwCJnSGce6TjyY1qO3goUNywHfv3DF4L11L/pfJeoKyI7uGVQzQALFB2M8rYlbBhAZEQuKpZlZY+qddskAYQIBoihmsA3qfYktJsqRbwMHI0LBY8wQDGFDWiH/DbCTw1/yHZC7ytzUHQQyNBw+kkQljjS4P6bADiHZ5jgAzHQje11fWYg/D32CIrK5rnXv7++LB5JTY+xQ8uM7du/dYn29rKyYnJ7U2xUgWUFVOPFs2SbhJxM3CzqFxqa1n0M+FpBoGbYZBatASmDd0nG3gab+tYETtoiJSes7GsePH1L462N8HAp8M8Pa4c+9eLMHWEesc1qT1RQlgWGOKJyV7QsJJUQYjTKK3KrZejyV90D8meIUpT1KX7AT2FV4VlhItgdNPrVPPe8HYcueEGW1yXCnZwr3pb7MI11okYN/ghAiaYHHwuRTEBK6k7BXsbvZ+Db6twODFxqFZIGgFzhNP/NKfvKzgUYmSE7Lm0GJL9eQA4wx29Lylre/ZHvVcNUQzAfeaNVIBEtdDouokwkUbg0s5+I+uHwV1WahIRFTXq+wSEHZDBbZiejRubkdBqjUYK95Gc+xxgqz5xwZK0fk2I13XltIvBCtqZ84EijTYrFK0vJfU5i+JsWQCV8BeyXjjvzofHTrnFKk4F7AUNRslhzIXwMz1aogjmrqpxalBoswz2doS2xE5E4Ir1h4ZOg1PTFkCAAh+T4W1jfVYWUMT34UrtVhnwcvpjJNeGBWSYqLQKe3zkP0BOOQ8SQqtgr4MLtWZoM4lEhEXtrAFNajR7eAGPSl2DO6yxrs6UpY8e4VrrACZa+Y9eakzgGLN8rLA25KdUju4o9GGzdFezVb+6q7w73vWC7YXe4k9Zo0VxmZXiZLuZJqQ0IlZWp1LyVDBFmlGBYBtC8vRgwBdRKe4UUGsC7QGRXkuBIN8DgXyKlS4INMs/jQ6cLKtWAV4gbRtYqHXMO3qfigmWQXLVRgC0DHjhmeyorkFdNyURJUTRxc0xDoXEcBMGxJAMe80hI7iMIw8GGlcd6eLfY1ZOI3H0GCys94lQ6R26wzSfc+2kbwqOauEqgL/WrcCOF9kp4o52VqA+EP27IU/w3739Yot7Eqnu0N0dlVkB8R2h1/tx+3sJkHyoiTmyCEK2PfkISdf/u9WdG5vx4G9Q3Hy6OFYW1nSXr9xazyezK1EO8Azw0iZ6QHxQfIs2NLtGB4Zlj40LE3Z4gQP1HnKuSchF9MTORWGSduv7927TzEEUjT4K4pymreT+SDFD5J0YixJHm55Jgvvy7qyv9fW0YwHhOqOAwcPxNzsM8VMVcQQA1pJGeCaJfeI9aTNC9ANK7jXkmh8DnJTKvI9ndPeOjx2SIAN+x8wlbPzYGJSe4s5VHfG74oNTXHVQ+89eN6612tphztUjGkkkP3oSfu8tZIjqhDR09PsYnL3Fiw/uiMtxYfevM4F0hbqajQD1Xt2S8DyxYsXVAjie9euXRW5xbNwXFAw0OcEtGyTEj8xSX1WDJB2WBt4oD9u3rqV3Uy2Zbw3NrNi5ZKk4L/cA3KePX29Mb26Go/nF/5N8oRDI8MxQoyNj1P3DvGzh4BzBgB3WUcRALIQKkkBWKpd2ZmViXoVo9S929GlGzaDsk3rqmeTxb46407ILbeh2WBJyKAwAwOyp7dD/n51eTPWVzejczuit30jTh7eHQdGe2LPUE9srq/Fgf1j8fHHV+Px7HwcPnUylje24srnN+PpwmqcfeWcQKaJB/dFZmLfDfQPxvTsrPbByLDj7nQrulcksNhjCwsrcXjsoLT3v/7225KOfTo7E9987924fv26/Bh5BJ1FzBz5xje+oTkrd+7ej29969348MMP49ncQnz/e+/HL37+C8Xzf/3X/1P8/oMPJRuLhCjyT8BHHZq14j1H4f78hXNx48ZNSabhk9jfFJQgYnGmDh8+rO4o9kwn9gRZMfnYdtl8OrA0i0HknNIrd8FQnZVr65J3oHOdfVoSOwA1gB3YA6Ro6KjEMA4wr219VXnUvv0H4tq1a/osQGh8Dd1ExLbMvZDMB4OUs8PQXe+C6BWTuBPJA8BZezoGPQfN89oOHTygziSKRpwt7gd7BmDzxuVLAnM5a7C/kavg2vGz1ZWDnycvo4AA+YduFIAbxUOrSDExp2JVMrqzs8+0HhQW5ec2sY+eRYe0FDNOICWpQ1Vd5BC2fN28kOpQzqCZOgz0XXLuSiGvq1vgPl6hurxd5LV0SNkF5ITKXvC9VhCPXIQ8q0ApbKEl2yyj2lp84Flgu/C/yrUl0+QZZxXrVQcLcRPPnX3FtRZ5hucOK/3o0SMevt7eFh99+JFsL/acteT9KFiJEZ/xL/uNAt/nX1yXzeMaGVZfOT0drtwDvlfvoRzAcVARjQSNbuUQ2DScxIA7KVqthYlWQ8j3XUx1PkYOXLamBn1zvcSq7BcrMaw2ZFQ9b7ElTikpnW46e1Z0DmWnIdGtrepehoZH4uHDB9rTJVtN/s49QqaDXMj3mW108vjhOHPmeExNTQioP3/unGbdrC4vx4XzF+PG9S/kP167eDE++/RTAfl0Yew7sDeuXrmiWSms8/j4eMzNLcSfU6j41W9jZGSv5J+ezMzKxlAI4EwUsWBxaUGgJftdM97S30F0pBD6aPqJ/g6w3hK4NYw4yUmNbnUXHjgvkvuLNsUP7HERZzSseFCF6coJ2W/+XXfKVJENKT11uGTuon2f8lKceQAAfFIxYZzHOUdD0sn22rE3BUc6Sbg31BDomIJcSOwOLrS26kHyXGB/f4+lo7LQwfmBWQ9JdnXN3cj4Lj5H8qjJzWFuFgVn4sW6J2wle2BxaUWFCjpZlOOqWOoCJHPBimjmIpqB9IwKMmX3/Ti+be5oY+6iU+XdZzDXkocXYUrd5bmW1fXt3LbkJysQcQGi/F1G8o04pWzSywOMZkbdGtvU/dTfiWgB8UXgPF0yzB5ybqSfZdFP15gE2nqmrdiF85Ui0z2PatgOJBG2yJJaspIutgSnCthdnco9+fee0T3yo54DsSF8b+bJtGJnzYhDFmn/PtlofBOYEfk236/O25rXI7xJ92O5UXIqyUIJ7/C18zclWQ/Rlj0iSeg2y0v5/lEt6NRe5L3ppLB/hWxs1QEIJIrFkrRneVPHq5INb7N9ffjgvofEd1oiEdtFURWcifyBcwbxifeHGE2uz3MoOSxsJDN1vypU/JuE2V+9yf9IKzC0ZPY3SY+DH9g0BgEL6OO/HNACecpgFnO/hhfWfUnblGBMw5E6dKhxjhqOuLGuKqfAtFVAqDUZH77PXAhpmM4vyakTVJ08eULOGPYTxojEHid7985dd2/AhCQZyGqnBpRFm5zek+knKnacO39ejDmqkHv37xUQjrySmOYpd4Ax4+AT8HFttCiSREhWZpPhqsNyYLzvobGxmJuZERhAAoBxA2SgWEHLJi1c83Noo26qqwDDQuEDKQJJn6gNv19FEJIXQA5JFmxTtNmIZ7PPoo3Ar9danWp5o7tj/lk8nZsT+EvRArDekigbMmbFuibIFZNCwSMMQZjkHWqXX5ifV9UV5j9MkMFBJCBcmeVZcV0YXdZ2/hmBkpld1sW3trvA7gR56xlXINXbCQtxM9Y21+PYsaMxP/8sBnp6oieHTYt1+mQ6ni7MSyO1EwA5HUA5RIIjydpoIFG3ZVvyGu/ev6cEhCRT7a26sjbJavX3egiX9mUOndX1kvRtW3e2JFFKr5u9rf2vuQIeSMzzIkk2wwTG8pafHT8Ty9RM85JVoLiBMzWY5LZqBXepOfmi897otihAPzsPuO/SrKzzV8yKFwF4FUC0Fl3MxDdoU5r9JUtlRngGsi2DPDnv/I3AT7UEu6DB/jND1cM5i5qtgBAGT1eXgjqBkCk75mKHwzrWnXVkTxYTvtaj9X52JjUVgVWhosFiySsosJd9oIAoA0M/b2wATDfvZ8Dc6ioBQOHF9YgZwYUmAyKjSjE96z05YyRFFBZrqCvBuvYIQ+lg4STwJfk3hlq3dKSxFuz5gwcPKKFQEL69LcCAwIe9d+bMWdm98fHbce7cuXg6+1SAmAqQOU/Cw2I9mJf3IFAT00XAkluHWU9AAvYp9kCFYbGTbH+5ZgourC33vrSyFr3Iqmxhp/q1p/VMAJZyoB37oAqb3G8F5groAWM1X8EatQ7uKFovCaiqTokm69hJikBuGDMUBnK/14yQGrjOfWJzWVPLHQHwOpAtcNNBdbJJs1BXCS6/gw3H5juozhJPJm9iqOQgM71nsfuy4M2z5vuaGZIdFSUjUC3xPp8G8Ws/ks+wJnv27tNA9FqvYjAXa7DAHp3HlH3C5mKjkB3k+WnWkdbL4DsMVnUuJetZAbVko/Cp/XqO+BM+6xnPn3OZHVLPnZ+WrIrrATSDnVegCtdcYH6r7SpyAtdU52knyLDzbNfzqvcuO6XA/Q/ISH3JZqbeP+uwf/8B+U4BJi2zKVQ8S7DW5wS7ZPC9o4tOHAp/Xk8VTVsKFXpO25sa/Lt7qD/Onz0VW+sGtz6/cTMWVtZjZXM7BkdGo70Tm4Dc3Hp096K9jOZ3b2ysYucM7LDfmFkl1nGXB3dGR07fzaRnaXFZHZh9vf1x7949MQA9Y8mzVjjXzMCiyPD48XQOtjUh4+TJU2LMsr+HhgYFXBDDQHx4+tQzmGBQsleKUdvMpdusSa/Byx6EyfrADu/q6hA4QtcokiD8LYN479697/cfGZKtQBubz0QuEzAHkJKkSgNoZbNc4ObvZZPbiYvcYcQeZs8B/KlgnN1fPAPZtS38LeevKQsgm92Yq9UefX0DLqgi3cAMsIF+nSN1krH2g4MaUCjW5sJCTEw8TCDGhT3OhhNGd17xb8vEuMhSRTr7w04liPj46zdu6OesBfuNWIk9WcU4wBpiB37eP9AbSxBIkFjKLqx/q9ifZ3tiz54Y7urSuuKHiEtg4NGJxX1x38QtZqduqKOXc+4ZFT0qpGLfRa7RgFMXzllXSQ4xwFTzJpqzjrhPyXHmbCWx4BtDzZEfG4yOboocy7G92RHdyGsuLsSJQ3vj4O6+2Fiejm+/92bcuTUeB/YfiuWlzfj81ngcPXM6xh9MxMradvQPj8b8ItKlXdG+TdEYUo9nNmk+DL5hcFCAPOtMpwWFYcB2ZhLMPVuK1149HxMTloQ4c+Z03Lx5U/f+zjtvx42b47G+vhp//t3vxv/z334o3/z2m2/Gf/7P/yXef/9PJe/2f/+3H8Rbl19TDPvzX/xc3UHf+pNvK8/48IOPJemysr6pzk58JXkHICqSbBVPE2cTP4jQpbkHlp4kJlAHGDHn2ppIC9X5inTsXXU4mC0uX5OSYLw3nQbkRmV3ZbeSJY38D8/0wcMJFXcEOuZ5O3XmrAr/v//970Vu4nnT2UnMzwDvkkpBFpX8wgOoDQAT6xXxjPNR8yO4B0sYebgoBRy6NMiR9lHQVLdRm+ZgUDB5/fXXBCB1pN/Ft8OOBchl7wEqiVHa0yOwhmfOi8G3zBERQzrlJjX7I7ufSpYVn6nuYoBsGN8U75L1S5HOMluOb3kGnAF18NNpy1qxt+kQ0qw7s3pxMPhWXuShJvuk7rjI5k2iDHFmST2x7qyVCgzJYLZMk7swAbAqftB7r6w2OhIMqrmYLWA2O+HcjWlJsOfY0alO4OK9LYzJRZuxtLAoOWXOBwU6ziU/o4BKzAawhq24ceOWbBk33E9HxSZscySCPTQc6U/2zHab2dqVE5QPrviCZ07cSRdB3XfZvNYYhO+1/rvAQRFfUvZVxYvsmOWz+R3WUxJYUiuA8e8uYQPJfhUs6sL7evRRPE9CnGSB+brbhTQ+A8CT9xdhbnVVMTwFbr5PUfH40bE4c+qoOijw9RTRbt68IV/z+uuvx7UrVyQ7R9fEk8dPJE124OAeScxpSHRHu/w7xaCFxeX4s7/4y/jVr34fu4ZHI9o64+69ByqwLmuuR3tDJYKcF+lHnju2WwoWfQy7Rv66K+YW5kW8EulQkjLNznkRQsFEUk9fSgPhzgLIU5wzziLnyCS+3sZ50RpnfgvYyjmv50U8444XFz/woXyt+JbCXbvnYzSeRYL2KGmQJ7IWfCbPHnvJfjJJloKhnxxdD3RmIBfZ3UWRlFjdWFIbhM3eXu1JCtMQFiSLTY7J3kuyWoO0py6A7di/1zO0uNliqc8vLMcqObu6SbsleaiOhm2kEV0o1v5uyDV5Bl+9j9ek9lzznpXnajuWNHJzV+pMPDejrWSQUt2gMXuuhapXrJVc1BfhADvjipedtdbP9r01bqAhZVtFqeoyb3SCtTzXuvdG14h2V3MOR8VujgVbPidPqNPumpP3vEyrrhFZZoD/vh6RoNmPnN0DB/a7wMasB+zxdigG5t+r66vyP2OHDwuLo7PpwcOH6oSqTnbsLHaYAhYxnuWbOyVTyr6yBL6xJ75kX4owht3eprsdKd2c9dKe9qi7W3N1uR8K4MrxqgOjp1c2F4yPF59JzFJyq+B0nAnI09wHL4r73Cc5A2sHdijFlKdPVdzDDpL/SHUFST/IjekzVDz5Svpp53H46t9/7CtAR0WrHEYTPHBbsYZHp5PHqGEQlJgko9qMFVr7GSbrIcNuA8xBiRoog0F3NbZMtgxEDyw+BtSsKtnm0BGMLy/SIsyBdgDB4SRpEkNZTLxQRbECIYwlDH0cIRrRBKxIQBFsjR06pGFZtBNrcO7Guhz1w4eTAvMJRvEpu0dHZSxKeqDkjAhmSj+ev+W6Dh88lEChnSbOf2bW7ccURW6O34pNMduomsKq7lXbtlhtS8v6XEC00q0XNojU0Pamrn9tZS0OHjigYgVgHSwQgsjHMzMeNKaBvil1hdHLYYsEKySdvDcD1UhQ0SE+fvx4smXQplzy0CF1u5hVDdsbvVKun2Fi3DPPga4N6bCngzeI2fDUje6KkjnSTAP0u3mmWwZZ6EBBnmAACQbmjgwNCcxZIcBJ7XSuhwRXnSCwllbR5kRnc8vJNnI7OfwL3U9kxmB5yX9LsoNBkbtkuKsdruQkmBvC3/M+rHc5CzMeLIfDG7EfFVqk/rvYW7BvYJilFAX3T3JVbE6KPgREPg/uGFE3RTr0aqV8kY1Qq7s/sBHtFIhXxQcFEXmdLwtOdn6/ANlKiKoQ1+RjeIhwokDNroMcUu1ADVkdSwApAVBjRFPiqRgZui8NFsyh41nEcqHD4AbrI5aQ5LQsU+PbTnbIywxo3rfTjudf3o4GuUv2qmwBAAs/I1nS88iKiZJmyQwRAoeCHBjObqNtSXIkU2YrxRo22Bsk0LDWeR8NW7fkihKEbK0Xy5FkMrsMOF8E0Xv37VHbqs6dAP4tnU+KLKR9DMHETsBgPnf+XPz+ww8SYHcHi3U1tsVkKukF9iGfT5CiLiOGxqeMGWeodN1VSNAwRYO4BXJLTzMH0nIvBlOQNUNz3HISBHey0/wspSU02DlnlLBuAI6SI8jBniS3sFXEasrHVjrvxWZmX7tQYb/QKplSTCz8C8kZ7FJLI1jCplrNBW4mM0cBN10WyTTEh/FzbDqF5zrndd4K2BGI29K+Xox/1gmbwfsyQ6gYmyrWqVvQyVkVEaTtnAVOmDkwMgGDKFRUIlCFitr3LlS4q0l7NNvH2S+ACtgqANXqZrKtdqcY/1/MePaFfGUvhdJ1+TD2Gf6O9WnYmHwWzyUn+b0arFusxgKT61rrb1rtUxUgikne+jutp7VsWev3xCATYPPls/2H4qluZAG6usWuZvi0umqSzV1xi4rKdBtk0YJPYM9qCKNAteT4aRkdjxcx9U8AACAASURBVEi4R2ZuS9JPQ/1dce70ydgzOqwuxcczszE9txBrW23RO7jLHUXtngMkLWniI2TQtkPgYnWSci4B6PH/0zMzLraLzQqAQOcBg6sP6BoeTT1SwqJClC7R3X1HjozpHgt8BO/GfjB8j+etGSxt7igTOI5E2+Kyu/2SKGIgI/dr2hNa2HmV9NO6Bkqb+MF7APIz/BN7evjQmIZ28/09u/fE8uqK/ClgiGdDWIYNYMd2lkKk7WB1HCCvAFu6CnUqEqbkifdC6gDvkP/guRajszqzdPa3DVCxwVWkYThsd3bsrq+pUKNBvwBVff1u91enhPXq3Qlg2SlejoFTD157J7u/8ndIHCkmU6jgmlhrzgOfU2QU9rOLFJ7h9nR9LR7Nz/+hLf2v/tmh4aE4NNCvuJJuI7vrjob0HnaIPQy4CZmjBhAj70VsqK7Ejg6RLtS5lwAi36s4MUd7NWbcVPcdf2vgE4KTiR0UQTa3LVfK+CCArt7Ojjhz5GBsrczE3qHuOH18TMOg19eJp9bj3sRUnDx3LiafTMfC8ka0ddNViHRJtwhB3NepU8cVlz56PK1Y8OzZswIL2RM8qzNnAemf6nkQQ3PfdHc8efRY559ht//405/FiRPHY+zQwfjFL38dr144r3j0t7/5TfzV97+neHdiYlKs9L6e7vjss080wPm111+PH/zgb2L/gYNx+uyZGB+/K9DcsocMQ3XBjTgAQgPa8awl1+LC27ZAXwhZFI7o6sBmcF34YAH+zKDYt1dFlX/6+S/UKUpR1bGXC9XkBJwxii4ujLuIxjPj844fP6bnDthag8o9w6JDUqVc3+9+/6GuEeAEAAj5WJ3hJMpISifJA81YrUK8EssjXgDk93wwgBuHZJY/Q35w5smM5iQ4kgoPLd69W4XZqceP1KnImWXPSLaCwdWg7NvJZEXPXkWMZ+pa403cNWeQU/GDOmrbtc78THMUkF3t7YllSXBuqbMTWyQ5TgD/7GbgurDB7DGeEc+AThLel/1mUorjvCKFsMYq/is2Tdm8jJ1MvnDRVXGB8t2mzIeGeSfAW/am7FHNqahOAUt+dTcK3lwzxcHypQCorL8JaM6/WcPl5UVJ1EEOq85prkFg/OCApIQlt4tkWxZdWAP8GfYdaT46hESMKsazSGqhQrbio+ZYobwek5j0TIj1MxYWG7/ij5bYowxe+f4CTuvf/Jd9VXmccwnH4pIU3jD5Tzkdsi/ZIef3aQKfFdPrnGi+jqXZnM+42x57wjlh3gPvBf7AdfM35JPsKTrwL7xyKk4dOxK3x29qLU+fOhW379xRHPjaq6/F+O1bknJ999334vNr17T+77zztXgoIuJAjI0d0ro/ePAwbt+9G5cvvxm//+DTGBwaQWgg7t5/qLybq5dsTQ4jJ4I+eGC/O56lRtGu7orKZWbmZlPONkmEGsJuAoiJhC7KqXNpkOKTC/mWDfNeaObLkPAgyeWsQPYJBI8kgvG3mi2qmMadrNXhxNpaS9/BlIuBlgek67tISc6nHGPwrMitHUO1Z6EiZdS23SUIqNzNPCdJlXEe2qyi0OGZqGxHCkpIOQlTyJklSAyLdEd3JNLSSCAzV49ZkkPYpG0VNugkIi6hQEGchrmVfUiJKhcqnd9WJ3Ur/NHMTSvTaY1nW4dnt7r51rmO7mByjNNk8Qu7qIHOCQ/84eJEy+dmJ0nlCWmZ65+Zqif9D/tU+TXniGefqgw84zpD1fVRBXN33RgbUByV5EafQT9bv1qLMI4/qwu9/r5+t4qf9ff8Hp2odB1iD1Ec4LlBxON89HSacEcBm+t6Njen3Bz5eAhC7HPyR/Y5sSr+h5hYkqJZjJLseFeXMDx39mDbq5vDPlFkX0gpdEvPPYuBQTBJcmT23i7F2jobIgD6/CkXymKuZ025a5ilLmIe3cfcY5Ec8DeoxIDfSfEDAhH5bnbNYQMgGoiI29Ehu8T1cu3gfPgLbBl+9atCxb86rP7qDf5HW4H9m3bwaLSVbl4FneqsyDYojLxAPvSJs91bTHRplhvI4uBjIGowqoIrzacoHT6S6X4ZDbPYnOiur8FocYsuxgUHCUsPQwCAjqG6dWtcIPuFCxdlUAEqitmj4LqjQ8UJgkyMPA4JZ0aBAIYgySxMfJz00aNHlTQzI6JARQyF9OdhDK2uyAFybQ8fPHQLmoAwS2vA0MBQTU1O6XqpeN66PS5HuHvfHrFyuHd+T4BBAjK0N1YQK+b19rYCLn4fTUsAeAJtKsc2jp7toQGd21saAs214WQxTLx/aZUSUACqFSuaqqwYR6srcfzYMSWiT2fQiCaQ9oBeAoeTJ08qiWJtp2dmlUwVoK/fSV3zVg1CrltBc3ZglNSXMqbUe6S6ffDQAbGWlhcXxKjqJyimjQ+2DoBOAm4wAeUkNjYNdmw5sakCCNVtQB/WYvLxIz1HtW3TjaEBtO0y0rCiSdI0kDuLBgRQBGTcv+QQNGxwWY6lAif2rZgmGnBKUoPmp5n6OCqujUo5L9hfo6N74ukMQ3rt1CS3tf28TIqB/hcPni0n3gDIc3/Uur7QRjxXHXj+N3Z2I1RFn48v1oIYkDlHgcSmBgCTcDUAO5KN7JohuDfroXWAbjFFHL9VQkuwQ7AJ2Id9MNjm/YHNQBd2dc3FsXo9d80tvagGbR3U+Hdq6Pjz91yBnCDeDOokSwXbgWcGeJJDwwlGVHAFsFOH16oARQFfUpEpjdPc5VWo0LBkgovOZPjmbIC21MFvYYWx39hDBb5V0l4MLBIg3kwdGmtrMTkxoRsCuGAOz9yzZ8nuGtD+JsAu9qV+keBM2rDrskMGzV0oIQjHPmhWhYZ0WhaHuyGI0cD7FtmDYslaTsAtygUIFlO+ZBBKlkXzXgD+sO85jJbMqjopuF8SBc0HSt12EgZeDfnAxlyHYrRXwJsDtnOYuSUNNmT78ScUabVfW6SfnIj5Wat4kT5G+4dEO2dcyMYng4lrRQZAzHpktihmJ2iua6b4lfrc+AN8A0FuaeM6+HQRpBhBAuxbug9hpyOfUd0c1UnQyq5kTaqjQp2LCvYrId/UDCgKLCSFLgR5GKvPojVQC/DVOZC2d0/Q6UORAxtIwKpXdk3VAPFWQKDOGcE7z661c8s6/M1BnvV3xXysrqy6l9bf3Wm/fBa8FxoFhdYuphcavC9/U8W3xhA89r3btpTAalA6nUbMPOpSzKHuyuyQWURCjOeWQ19tWTKNMx4YHW1bKjaM7R+N0V39MTJEIrIYj57MxPTsfERXb7TRxaiCpbsY8SNcE9r2MGpVGCPJ6umJZwvzsXff/8vem/zYeWZpfiduzCMZAxmcJ0mkKA5KDVSmpMpMZdbkMmDAC6/cK6971ZuGvfHCG8OGgV4ZBgz/AW2gYAOFMsrV2eXsKmSXlCkpJaYGSpQ4j8EhGPM8GL/nOefeSyaVpaxG1gAwClmkghH3fvf73ve8Z3iGScVBWFLyfOnu0vnjwWCIIcoaF0uw5C+klcu+QRpqQp9vbtbGe/wOa6uYTuQozbWIIWZPt4xRQXVyy2WonWd4NTh4FryXG34bavzWfeL+0NCGBcbvM1QhH3GzzD4mQirnIIjCTIVaV7dMLGvYJ0QwqM40h+We3b4zZcZZDjhr8FXhv9Y0z8Z657mEEyUpFl9qD9NQqyE1sZUmJShhNYWXrZ1/5MhRsTx4HjSWQNwXKMcyA+kJlXR7blQV0mUgyZ/8LIMh8jeazPLtybhmdDKf240bN9EGYmppKR4tw4D63X9NDA3GXhCxmI0u8J4NMWdp3vB56nrJL8mHieV8JlCu3DP2Tpm7e+jUkglRrEngAvfe3j/ILgEwctPLA3LHf/Yc/9Y32Btry+sCrpw6/nxsLM3GsQMTMf/gbnQ31jU42NrsiHsPZuL67bvxwosnY3p+Ib68dC1WNyL27N2vxu6d2zcF3MFj4sbN2ynRsBHPPf9c3LhxXe/PtZOHC7LS0YivL12N4cEBNSCPHz8e7733izhx4nnl2ddv3IjXXntV5vAgLV977TUxbW7dvBknXzqpOua9X3wQP/7h91VjfPrJZ/FH/9mP48GDRzL2fuv33o5r18zqXV7bkMwJ5yfxgDzhpZMn4vMLFzQ4cszt0Ofg3jH0wE/jo/Pn0wzb55Bk2TpCRtlIQ33yyac6uzl3iGlq+AVyV8jZDmrPstZYy5xTfP4CisGooKHBl5iseEWkvwXx54sLXzT9iJCjIb5RCxnPYVQsZ5gnVol6T68Zo6j9WYTuVr1kVrrQx2pYrsuXRIOw+TkNG/gi5hE/OJ8OHDyoxjiDMmIZvhoaduUwsUxlCxDH/VvdWJMEiWKXWArEJhsMm9nvmoj9Sq0A80X3II2VzXam8WqABs/GDf5usbEsi7OsZjXNdl1DsjiVv+SQoqRynP+2WAE6/5KN5Lwz/XeSOajnnN4LzjXMnK4moBlKvo/1+XjNAndoPWQ+y5lTagCsB5goShG3NxWDufcMrOwjlg03zGZXlhXDuM6SVKI+6+vtFxMHJh5rmLwNBr4akukFWEAM7NY93K3s3DmcQAM5rOGZ0EAsQFENP3XmtoET6u91ZlSkpLlfgwfnRwbY+D18KPDMxYomF+4sVkteU75Hey2Clwn1PfUb9Rr7h31P7KKmFzNxxw79u3LP0VH93N07d+PF48fi+NGD8qXgWukfwLRgrcOo+PSTT9S8fPPNN+PTzz7Vun7j9VdjSiy+eQ0gj584rhzvwUMkaXrj5z//MEZHd8XK2kbcun03pmdmtf/oNZDXU8PyjDhPeIY1xGPNUyNHZ0P+DjY8N2sdCUrWjxmyK02WBOtN+WxJ65T3QP6e/C3ybPeeMbDB3qTOIdQ0zf1Zfxo8ZBCUPQwZZLVye9iZsJ0EktOeo+GPhKtrDnJW6k/yVfIinjvP1QCwEAOOfAFghth1MGcA73SQXzHkNHOwt6dP6gwGga5ZUjyBQ/Ze65KRt4BzG7xvVwwOD8bs3KIkvcUo7exWTkMglFKD8kTHlxqAPe0k9xyjNaio5d1iVDxendePthiJDrTV/K9mfuXJzUZ+vvDj0J7HTalbGW1Oh9ty3GYy1f4hUk1E3+JzyF/COXKtt9qzquczX7bfglVXzFxJk/amV4j7Bq7Ls5Zv1oLOu6ouqp6A3q85nPEAhGfKGWhzb/s/VDzj/VkrqlsYLAn4AosflrBjKP9jPdDLYcjPWUduiBw4MVr9MrygUqKR2M/vTONrmOyt1eVVfW5i6dSdu4qf8jxF6aS/P9bKzB1AQIf9E+m70b9Sr4t+GIM42NI5yFZ9i1fZwweOZV2duj5YEnzR++Oesj+IK3zBfuR+MoguXzB6fOw7AJL0EGDMqRf6jFHxu0+6n73DP+wdmNxqyVa4EDGDQgmUilB/rxoUbCCa3xSmoBIYDNBAk9a6DGVaE30FeiEyrOXKYUp+Q1EhI+J1dFaRJeHfO+LgoYOSVUIv9vLly0pqaaSDqkEWhUB26tRpXR/md6aqRvSTaCYCfGhgUMUpSa0S8EZHnDh+Iu7evRN3pu4KZQXaiiEDwwsSRk0puzrlUUHRS0FLAs1nhMJKIgBdFJ1ipqo2s5kRCgPGxujYmIYeUGwp+jGylBSTjEwtmcOhT8ICEsZFBEhl69mp6dbZITPs5cWl2CkdUTdbeS2QlzQuQQcpUFJYYsKWVHISMGicKkiGh9OYFXMqjPQ6RUsjGRmEmbJiYzWZ+i4uqhECitdSQej8Gp0E4grWiocFbjRZ3sC6xHyPgGzkj9HOQmBJj3471jbWYnLPbiEloO8ji4GusJB2HR2xuLIs2Qxs6jghnfysCe6OXBfXRgnYhcwGZpmdnWr+YG77aHYm5WCM3gAppPWYdNVC4YjR0AUNeVWDGIK6KOxChxttUoVC6VwX3ZPPwOvx/UJXCekjWl8IIVsJdCXPldjXRP3JxPzxnd3e9K8D3QMAIRWE/k0jWyHNEh39RHgoRkh7k6f1Iz7wedEmUyoRD+XpYjRU+ltkw7X9uqWd3yZHpYQlC2cVRzRdO4x6JXkwCi8Tr1xnHJ4wnpzUVomTV9nGrHDTNxkEqavf3s9sR5UUc4TGoqml1osUPZyCNT0HhP4PJwok9SQt/EmiwJcHNmZV6UvX4waoUOtqhDa0BkrSikSF5FfeJhSTgSnooqUSmtJUbiozmD14YJ/+nb3Gfro7heG6mQokUiQYNKdpBi7MLcSIaKItA3sXqx6EqSmuItuIfJovLm5susznpygTbR+/gWzAc2GsEYoy/iSGqpk654K2BsrClUumYlnNP0sAuelBoe3Ybw+bnu7eNGWlGEEzdr5pWE6xqya6Ckwns4oj7QV8rj0PNlzQGD1FMwSdeRBnmzortLfahlYaMhKbqtksSRI3JxSrkH6iMAVh0oZsrP3N6xoZbAS7hgAUiMkKZK+zpjh71JxhjajQ8vDRxZsbJ4X4k6a1fEkGVWBa89dIS7F8SiJN552lGQq5zHC/9mjpksrnQHJQK22mmyD5/Xpe2/6ThJvzjPMI2ScQQvoqRNhvYC9UnCuJEqF/ksZdQ8DW9mgVXjTIuGbWSnvMeBL91T6oeNqg49tmPOWfxM+3S2dVHMZoks979uWzyiEeTj9Uox0gBc8PrfgWDd3rSWg5LRp7VPDfzx3aG71dHTHY631x/cadmMVMu6Mz+mni79iheMawWuatjU7lKt2NTklKqnGw7mIJvW/WGoxL2JAgnFeWOWN7JF0wMT6h54k0SSGUaThVIx3TR9gPQl51dsXKiqUFa7DuRuF2zDx6FDBO+DnkJTwY9ZoTMjBRbmWYrRwgm1Cck5aOI171Ki4gO8lz5PwbHxuT9CbPGykcPt/V6zcCDxA8MWjmkJdQbEkehGFSyjkIaQ5gpbNTZ6ZReG4SOl90jlQIu4rJOltygFIoMj53FXvkTiUrQE4D4tL7y8bZNGvPnj1rr42ZR3Hx4lcxNXXXJsWKB5ZHrHyM2MX9rYKeOOEhuYd1yAkgq3XhwhfSA6+Yws8TD8mFkWPC0+f+6mpMc///Ab/GBgbi5N7dcefOPUnwsJ7J6wT6WF3VgIKYyFmjRkGaVJbOMrFKfmCwIpCc6bHUHI1egTrERLEZZX3VcKuJ3m50iomLnMfa2kp0YUy5sR5H9u2NWFuMXcMjMdC9GXsnd8TC3HyMTuyOG7fuxteXb8WR54+o8f/F11djfaszBodHYmLXRNy8djUWF1bi9OkTGubj/QCoav/BfVrjHg6BFibvdhPy4sUrcfDgnrh2/Va8ce71eIih7dKSWBiXYTtvbsZLJ19Sbg074YfvvBMf/OL9WFhajh/83lvx5//PX6hGeef7b8Zf/fufRndfZ/zxH/9J/OQnfxVnX345vvr6Unx9+aobzelvxt+RHn39tVfjo/O/itUVnj/ngRt0RM2xnTtj7949YrhIPquzEcM7RsSG44uzudYnwy+DB8r/ifOqW+dRybBSY1B3SPp1cSGOHjkqxgzNUUlB5PnB+79w/AXlInxe1sPswmKM7hiJg4cO63qQxmV9SIKl8o3MZYgLAjsIwWlGO3mHpYwK7GFwBLk6zXLW046RIYHJWIxmlC6budPVHadPnZGJd/MMXPaQS2sKLxrkNocG7c3X3xfTM8iUdYgZIpZnF034brFX8IOQ75g0xZEuGoy5bErZe8LSQGoaKY8wctxypwCNeiS1wT0kpvB+XIO8I9bdDK3YInYaDSnkYto8KjRUyDgmAF8yP4ihqqkxxU4kugcQLdNiDUwTPatGJZJ8nFXJlnBu78EHn4HXIl8UqA4lgR5fH7EdObSXTiI51ND5h99D01ejcgVkVIYGVGPxmjTEQAbPzIBKNutQdV75UQhQ5pqppZP/eAOW4Q45iLyzOhpioxfCukDb7QjrFvDN+WYm3/qdgUGbZVuCx55iksVccrOuhnQ8Vxp4Zi2liXMBlxKMIom+lKqs65HPnLwwPFiv/EeARiQ3QS/v3KnvI5F84rkjcfzoIfUQiPX4aF69ckX57uvnzkmKjdzr1OlTceXatbh35068+p0zqr+XlxbVgC8wyMuvvKaB0N/+7S9idHQi1ja3JV231QFos9f+AACMaGROP/TgN9nHDE+WYNpSw0aHpKB5XuXhptwqpbA9ZHMNwmvBXpAqWnm5JWiImFPrQDlcNqllpr5sHxvuIc+gQFB8llLN0BmZ570GWEqpfG7WsEPN5QQUKdfIHgHXu7nhASNntsBDfV0absp3L5+vJB2pK8mLNumL8HMDsbRsXyYGMyDRBaJYXQ+8PTi3WJOSYu2xhBg3p5jH9FO2thoBk5RBhfZ01lxmn/rc98CStdVMDX7tVG/D2TUHcfW9Vi7c2i+VUzsOWMpTQ2Bqj6Y8XKvJ736CWb+Vn9TAopioTsC/IeHI33/yX5vXRq0tWrHrzMrR698Vm9q9JBLQwc/zGQSGSV82Pg/PoQCx/Jv3pmsm/q4InHJtrv0M9tK/ZX0l4AfDqYaH8Txf7g89KcnA5QCJ2MU5WP0bGBXyZe3o0EBPwKSNDfUoT516SXm26hFAp7OzAjPAKhRQQ7FnUO/R7A81OmNmekbgHe8BS1hznhCHyJOot6kDBJjFP7WnV2sPyVd95pS/5pqJo8QKyTbpnJzXeUbORZ7KfpMJ98aGzkpYiNzP+owvvvii4g15AEoo9PvIbzS4UX639GxQ8Q+Ydz97q3+gO8CgQrId0vvdUFCo4MPBxOZkk7MRKmHg73XgGO3phlUh4NlsbGBo3/x7IX9VkDJ9TxSeaYQ0h9yUAzFEc5uCgyIJijIFJzqM6BrqZzEcY+POzxvAD8qm09roHHgcuhRBTOMJYvw+BQ/NnjJHIig8fDjdROcRPLh2NO2gg4qt0N9vnXAM64TSt/TGytKyEBUMaAh4IJ5Iogh2NPEYVpD0o9PKl9kloWuwdMuW0P/FWjACtCeWV5fV3FcCQBMLPd40WqIh6GbCtoKcaJuJQOKecO+Zwpbsik+sMq5Nv4A8aKuBy/uq8T83p+ZJ6aFqQp10Ue5BTdjVQEi9Rg7uoibLiFJIfSfTPdVI7ekMTI3HaLrSMF1ZjZFBqO8D0hmeW1rQ8CU6GFAYzUyhvLgwH/29yFux9mxyJU1WGpEb60I4k6BV05jgzzMo7VmegTUAt5Usc5gsLC75fqdZL+tZFOVEiHBIcShUsstZyeHC+uH+grSROZy0m0HEYmC2rCKVtSg5KFCFiSAQUigbg0U7Vh7RRF94vwnJ3pRUKmSGC5UnqZ9uIBeKybJKeiYqwtxEqOZJNTxB5Pp9nfwWAlXFVqJUi/WhPUBTK/UV6/eaYSgnDCU3wF4SiiwHFYVuZn8XalUUS8yq0Dtet3dDXXexSdoHBFxTIUtUpyiBe4JRkUyLZvJWqBFTK/Q7JB9qDmvYB4XZRpD6jAyf2McMTmgUw5Zq0mWLntrK+fw+DRUbHtJ06LM0G++wogZtTFfI3krqafBxr0vvn2fgtdLTjF2ihVIMg5hX89zICyf8bupVDJF+cjdanZbEY7+XXqx07btM8y6pJBL+en2SMq6L+OR760oQnx0QeDbeNiOON6ehpeFMDgit92w5JzVMc1hdcZB9wftaFmm7iWis9ekhpxPuQg2Z3ZDnCkiqroZMQBlU8DMeum7oWiTX1KbzXsMIxZ1sXLcjxmu4BFJOA7D0ZmFvS3ZnA0SwvTVgiohynM15kFoYU7JWaLi4SWEUYX0OyUElQobzU00QGglZONEUEqow/XzcGM6iPPV9rYdqRGINTLkuBjQ0asoLhXvPsygjae2rqkzSLJsYyPm0l0HFvLWLbSBtFGMxKp5MK6oYo7Bol2us4qOGDO2NgCquFPezydAchOYbVJHz5KCjPV49+Tt1bU8OOur7GqbJ9NdDKaRRADjwbMR8S2Nm/AQ0fOtA73jesgQM/SUVYUq7B4rJyBCrCm1lYuR2jO8ciqHenpgY26lnPD0zF1MP52Ibs9XegejREGre0lyJ7ATRBD2dZpcbuvhDDep9+gcH1TTCt6WhmIZ8xaAGFUgpsZZAtJIz0dyw+Z4H/sjG8ewosHit1RUK+97YuXNUqK37D+7H8PCgnjmSWGiJY9iJoWwxZLX2EmBQABSvYzeDYGPxdyOTN2Ln6I7YO7knrl69agbqgQNq2ADQQNaF+3n/wQOduzDCpqbuxejoDqG9/OyQ/0xTUL1JR2zLANDNRqPwzRByoepGIv9W51g1BpXnJPuDvVTSL4L/cW8H+t3Uk4SaVwo/IwBDPid+j0EGjS5JW4jSb+1krleDV5qcyWryum6dp+Qh+BgMjwzFl19+JcCFpaW6ddaUTMjm5lo8QuIqEc5P7rXf9X/vYVg00B/T08R6mKOWzatBEAhCniHLnvy6q8usVJqUAiMxdExmFQMefkbnfMZssUyFSnUzw3Hcz48X5TUY5oCaJfbF5lYMDfTE/l3jMdDYio2luTjz4nPx8N7d6B8YjO6+gbh1974Ywrsn98fi6lp8eelmjO3axa9a8hVPDaEbzYTraHRJ1gcWM/FRHnLr6/KtQT6NeHT9xm0xG27fuaO1s3fP3rh955b2O0yMr7++En293fGdl78Tf/bnfxGnX3ox9u7ZHT/96V/HG989p7Xz0S8/irfffkPDjMtXrsSePXvV1Cf/vHnzTly+di2l2szms1Z+p/xc2Mu1pmkQ2mTWeRioTb4K8UlMUkM4h3BsF5+j68oV2Edmf27ErnGzq27cuKmmSpkE1+Dt5MmTcefOHcljSQYt5Yd4LYzlzTb5Wt5/1DmWnuiX/0rJpsBeZn+7MWj5EtZSsbbcxPY+5d4rBsK+S7ABOYL3kw1DzfjyQJg8m/cln4JJxlrEn0PSkMrDbOLK/SQei23PvuzC8Mb1R/l2kAeRG6iRLRapBwI0mvsGBwXq4r4SG3h9Ic7VXGLdupHK9Sk/ywEnXh3UDLxusU3ll5dgjYpNhoVSDQAAIABJREFUWvvaFUYgK4YkaMJsyw7J3fJzHjYhI5syo3kel5ykagohk0uJoKSvDAjToCrPq7oOr6UW87j+jt8jZwE5D4NzDcrWViVTVrmkchTkkwb7My/uFAOUoSbST8Q1zkg+twERjo+cmKyNZv7eFsyUg2XTtX1Ao8FKSoZW/lQAnMoDKz+onJDYNDBgJLLzYUud1GCJ85jmOs+Ta3UeWM3QRHE3B8xeQ0J/dzR0j3kWxBHyPhr/HjxlXpZoetaDAHYND3tOHDsSp048Hxc+/0wx8tixYzLTJlay5y58cSFW1lbije99T8oKc7Mz8eYb5+LLz2FWLcb+fXuVXzMkfO6FF2JwaCTOf/ypBhUwKlBKWNugQPfn5HXpmxTLili6sbauPJXJM9eLNN4DtPlTZ1/necZh1ilxhxyQPebeDDWHQQEazvVgGA/7wLKq3FPqIvZSycZKhm0D37NBPQ/1chqcpdbd5wJrjyoHyzUBI4/95VrCeYX3gnV3CyyysQFw1VKM5HQllUvsYvgISMN7DDm2ZUlKi33cwcABtQh7uK1jpt3ZJYAq99mAJ+qGJfVvSjqKwQZnHpeB783CIoC1TQEiheVILyaz+h37pCSi77vZ7u9n9p2qx/4vr73HpwX+wSeHHFVrFCvBP+N9VpLqtS8K6Lqt4U5+Fbui3WPiWyYXlVu3hhR5jTyajNOVl1cs41lYacJ9CfYbP+Ohpns0zpk8eKnBq+JUDh58yY67Fb/Uc8zhsZhuWUO5jresOuwH1gu5TIH1AB3QK6Kup89H/kW9pPo3PdKI86xtgAusdRixMMoY8IqpqPrALDYNOxnMAUodGhKwlSEC5zDnjCXFAWy6V1pflk5jYO36UJ89wWr25jUD2Sbp9ptkSMorKL/XeyNNuKn+k+RSgyH9imp8zsrqwekzZt7Ma8Loqs8AqIL7y71QLvyMUfEtd8OzH/tncwfGVje0EavJJ2RG0kWNrLR+bwUvBaFEVqlhQZAtSZc88CsxFQKDxmceYZ7wu+FEEULD3sjQbaFaaPby+hxYMlElOd+1W815DJa4Dg5JCnpo2bAd1Njb3tQhSxH9CGql2BVuSDGRdKIWMmcjYSRoYV4FO6IkOWgEUfwQPDHiIQgQpKCKy8QpaY7Dg8NKcPjsNL/5k6RQBngbGzGxe5cCjE16fMjRWKC5BGOjvkBLELh9AIBw3pS+I4mgingZrKI7umyfBAziVp3sYkDNAcrPUASRZPIniMWaVuvgIIim9iFFFCiFohfzOZXwYEq0hrbuoP5O8ScE0Pq6DoN6dqyJ0oj2Z0L73kMXDgRTvzuiK4sYPDcYzgzQdAH1ubGpwgqjWIY6eFiIYo7h5tpGzD6ycR4HMs80UwUNptAR5gvcOw0ZGBU0dkXJyyEF18chSqOIqTj3m/tKsi0NS5KwbIpo3XKoZvOykGo1HODNZWqWe4HkRx4poHAG+uPhfZ6diwUSXstrGE1SQ4oqHrx2/H4u8PyndbzT1PoxxkrpjLZ0IN3gdRNUKJVE8jcRCNnQbm/8qUgAxSX0pAtJEgpLtRlhUmiMllSQm7XtX9XgbDVrQ/e+1m01/CSbk54QzSIqEzz2XJlpq2Bpyjo1O+ZNhLg+ayYDdfgrscvsUId8FtB6Xnmx1UDmAwtFletfz7oa3PnDGnAiZdJEjhvJUe+hxLrZtAJxlmh3Je42n5OWLAUBRlZqjPl5eV3ZMJPvUXToGWRSW4iVSnL4LEpqpDNpSQOzlrZUaPBEaBrxWLi+l8++rGIcxlkNmygaNNgTOqxbQ1m+GIwKDZWmncXEUONP8cSeGhq2Cmllk8iSBhjZMaK/8yeN0vrcMhcTQ8NJVTFa+NkyUZRXRxpZtiemXstOakuai2eh4U2idrnfxFK/v5M4rV3Qvtm0VHxL4zMZOKbBeHMgITPuEaFj6h4TYymImvIBnZ1C2ZOA0hDwfBG0OmaKg7onDDmtbd1q5lZx7ETbgx0ZK0sKEam5Hr0354hZGNa8V0Gd5nJ8nmr4uMhxkkujBOYNxSmITgpIkHsMPti70t7NuFXnLPJ3/G6x/lg3/I/34/q4NzwwAxASudSktJud4IaUGwNqUuUAqf3ZfdMAoX7maUlPnTPtw41qmlSc+LbJkpo6xczJwk7PIs+xen4g6QE7sC/YD8i08PxoCNS9q6KC3+dc5LmkD2uM7xiM4YHeGBno1xqduj8d03OLsckB3dVj9pMYhjQVi13lGMuXNZzNDirZyPsPvQ6RHQBMwXnL7/JcGVZcu35VyCzOL85s7g3n8t69uzUYZBjAAGN1jf3KNYyooXb/4X0hmGna2Oi6P2Zm5yQDJKQjqOqeLsvyZaFZTT3O7RqiauisQX6nEI2sXxq9fO3bs0eFEc0OmRmur6kRyIpVQ4TPg2wDKH013WzuWetbLIqODiF2a6juRrcH7UbEutDjf8V2aoFfcijRP6DBIblONxrFOaj3MNgDZzcOjVimaS7t+85GkwHrs8PFsots57bN16gTpZhIeT3ojNPcu3btmpohxD1Yp4OD/ULA9fb3xr25+bj60LnBP9bXsYnxaOCVBLJ0GSm+JYMhkA9YWYneHgNrLPXmxoriAjEkJdR4LiAYiTvW469Y6zPIMcSG22ILJPJaxTxa9sTZrga95Xjj1bOxf/dofPXJ+ZgcHY6u7U0NADu7e+Lew0exvt0RD6cfxclTZ2JpdSOu3bwbW40uGdazR5BPoZkFE2F2dk7yT2iKv/zK2fj88wsqznlUr776Wty8cVODo9u3bglcRe6PVwL1Arn9J59+KmklAFG/+uTz+P7vvanXvHzpUvzxH/9RfPbpp4oRp0+diumH9+P27Ttx6qUXde4h1fKdV76jBteVK9ek+9OHX9ymZd74ooHCsF0Sk5lPEMMZkFXDmngOSIr4rLyfPASmeUeHDKhp4J//1a+a3mnEYTUBt7fjyOFD+v7Vazcyp/C+UM3Q1SmZK3w2YEmKGaE8vUd5AJ+bs/DK1at6tgyKkKmjvgDMVRK+5Dfsv2In8tmRXtFZJ3amB1TkkKo12ph6Pue8tyzf6EYNa4GcBFaP/bI8cMQHh/tgDwmvQTV0knVV9dNGbMqnQkAv+XpsSu6l5OWIg+3gHsm7Zs5ZOYMkXlI6yuegpbMElsszhfDOXtae0Bq29I1ydrGE3YQrT6qqMZrNyWIHczbkYKokXrhmx1eftcUoqLPTjTozGfn8HuTaS6fOlJKHcrwyIKRkXFVLytOK/WfAofxiGLqoVjOb2dIprm8kEyRPHZhU63H//kMxlnjGTtNT5klSLRnPm8OrHOTWcDkDXisj912xV5kbj8Wa5V8s1RZWHlCt5jyJLwNHXJ+SP9Nsr9qtzpQC1hDH+KqBUcXdZqMXb4ruHhnGw2Su4UnlkdwvMxGcn9G8570Z4HH2s0defOFYvHXu1Zi6e0eDS/bwvakpfUDkBS9+fVGDitffeCO+uvS1kNFvvfFGXLl0SUOj5587qrwQzzL8DU+dPhPvvfdB7BxlMLYu6adHcwtqmjcZK7prHXHu3Gs632FwbDBwyAExfgqPAGSmz6aHF2azcF3sD2pWGq4yI5Y/h9cS65BGKIPrYu0CyuNeq4bL/5m9Y+Y1a6ZUF2TMzUCV6+myD59BOL76p+WJFf94oWq+a+9JQpHrzno38zn+W7Jc/X0eBGcBtbQwr/fDDHl5BcbgRkpebal/RB4iqSfVM9vKU6j/a4ZQQ03i+NISPoUbQr4vrxAHuj2QSMm1AhFVz6sa296z+v+/Nrh4clDheu5JiSav0hpgFFhQw8B2WkRzIJFsiqclFVWuZ23bnlPrObT9e8XmGtRV7OEZCIyQ4Dheg/2h/JBaOPe41kWTkfNkp6DVwK83bfYB8hqaYKnm/TBQpHUvHWdq/XgdUhvb3L7iI2dqMcj4XQ2jAR2Sd9tg0msqWWtcBz26vXv2NOMKa1egi6xlkafmLK7BCj0kgQm6euwRpeGbATjkOBoCJ2MRIHExTu3bZkllYm5di4CinZ06j/kif+Rskq/SyrLUWe7dmxI4lp9hOAhrgvNZg+6UuGRgwXUQ94iJGp6LjWkWmjxSnw0qnrZTnn3vn/MdGF9LwyAhZY2sL0d6Nq0Dfk1C0VCkuW1acTUfOITry80gN2cLkUNhq4CnwgbzWcydhnUIGZXj5AA2xYED++PmjevWC+0fENoHhsbNW7eVaCIPRcFMwUgSQbOc/6NxQIJDMotsAQexjZFMF+Z9aO5BtYYRAfoKSZFKWAgOUKkoyEFLktiTuCBrwBfBR/qeG0YMEbxoGGqaScNLRnqDQhpjsgcCQrRj/BWYhHYh/bRLCQuflWSmKKsqlmk+bW3ovgjRhKZqym7VgVH3mfvohHQzzVOXVTgx/Kgg6YPQhbhRtS5WSWILWeTDiMPeAa8MKHmufF/G3RkMZdqT6BMxbHK98NlEXdNwZVOo0rV1awWC8CQR7iBBApkxMChZqxlQZDQFpdVnSY6Z6UdpjGp93P6+gWyyk3wMWfsWxszycjycmbZ5aaMzetOPgs9CQSEKYBoBc58kxUFW12ZKLVRAMhEwWgcdKskDCoDNDa0hkDAUdEKQ0CBaXdMAanI3a+SOmpLViC2aazujooYAGkpk0erBhtdk+4Fce6eGF62EqFAahYB3MtCU1OGQbUM0e5hkNJzuh5K41uFLQsQz5FBrNpKbjRm/rhBTnj5kMlWsD19Dof/KyJTkxk0wD1FoqjWlsKQHvKEilftaTaj6vO0jkWqY1Xu7AeLUrRLn9jhbTcFmepSI+E4lF2Wkbd+MJoojZQUoByjk1zbXHQN6QF0ZiQsCA3ZSU+ZHH9r/RrMTRhCJLU0cJfDVYJNHw6piWv0sDXdTvs3GUWNCNFSaCNZCJcnhq4z8ilLNeqfxwWcfHRuVzBvNSf6bdUhTk/hSSV1Hl00lXehyndZ7NRIStty6jWUH+vW77BOh/BLNSdygACNOqvE4OKh9VybaQsYhE4CEljTgOxXHlUjBLsjPZskCN82VCOfar4GpWVKWdyhUHd8ro3Ajm+09sWt8XOuHBqd0vGuI2yY/ooJavhC9LW1ZNT2QYRlOz4CWeTyyOs0hYiGpheayoSlfPD/5ADQ61OjzkM7/1jIc9KBPCMXUa6cprqFxT8ujwsWOt5SRpvZt8tnohg6a2py7tX9psPGMtT7SEJh7XHtWhYb0c/06aIJzHawFNRgXF/SaQs+lOWANKCruCb2aDVs+eyGbfG4YkabP26Rit6QVnpbvfNPQoRoG/I5ixGM6tC0ZmW+XQ7nRY1R3aulqMMm6xVzejIBTJ0/qXiGDUoNaGmKglyueaF/kucBaMfXe93PPrp0xggRST6eGlFev3oyFlfXY7OiOkdFRNcF4HgzNeX5uFllqDAlGzigKHO7h6Pi4YsDN27ezqWcUGgUKcXF055hYCUZIdfucK/O92NIZyvq+dw8ZRhBcZvXt3btPhQyF0/q6B1rIv/G69x881GtrSJItMfIW9h33h2Ed5zmNCQow9qoGPvmsZUKYcp96jYzvxW4QQKPLDClyslqnLHIzuNZ1zX4PhkXIj2zpLGZ/k2vxp4edZhXxs9VsUqNIrJJC6FnyCRaKf4/4DYjC2vd8udFX7LVQoXfmzFmvibW1+Pj8x/YNyDXfGgy7aaiBXg4ry2fIzTmfmQwqMAe+cfO691x3l4pKnhV54cTu8Xjvq8tmif4jfvFsX9g5GusrqxqyLi5YGoV8nWuDBeIhGJ5DvWokbsJoTU1ms3BCyD/OFwBAyuWzucD9LC83Nw9txM25UDUBg4Ut5BE7O+KVsydi/+6xeHT7Zgx0dkTH+nqcePF4fH3pSoxOTsaXly7HzMxcvPLa67GythX/4WfvxdpmRxw59pzWwMfnP9XA43vffSWm7j2I6zfvyDDzBz/8Qbz77s810GVdv/3223Ht6tWmlj1SaKxj8rtf/vJ8vHz2tHLz69dvx9tvfTd+9QnyTGvx+uuvxcUvv1TOf+7117UPkUL6oz/8w/j0s8/j7u0b8c6PfxQfvP9xTN2bije+90Y8uI/pN2yTTf1d2ucybe2KAwf3C0RFIwIcin2RGjJtxcQb5tXnX3wRvTT6dYauRkN7ZlO/y7+fP/8rMSJ0bifamLW4Z+9e5W4ArNgDPAfOcw3SpUOPabzRomqISNYOduSS9L4vfH5BAC1iKPkG58zNW7e0z5T/djn+KKdI40/leSTr2XSWBGkyqsUWrkFFdt28nz1QriYUjXI2K/uT3GpxwTKsfDFc4dxliKI6KH0yCvTBa6xtrAb5jdCpCbBAAoZ4Re0xNEjzpo0phfQQ+Y5yYQa2NgE3g5JhvL0sCrC0seX4J5mp3l6xTlWnZW6nvG3dQ3wNi1cxo4Z5bvlYs8Gch9TrygMoz7zS7yfSVK7keGsZ1RoQc328lwdfrrOruVyDFeVUNOdUc/s8rLOcc8yMM+cpxCUa29TfYiu3SSY6RNnge8fIDp2NszNzejZL1KudIPArB3duL09BrceWL5IWSg4qdW1tjdY6e7jn9bkN2JtQLOcc0QAsQS2sGZ2dDFZSZ17DpbwOSVMm2IwPKdPZ/G/uAzkt94yzi/OvcjZqUHJehg/EC1hR5I1CSCdojBxCzXaklBj0DJhNjET066+ciecOH4jxsZ2Skb129YoGFcTGU6dfii++/ELguR/86J345LNPtT/feuO7ce3adQ08kUtkfz6afqiz/uhzL4hRMTAwIv8+GFDTgCaTcU7dBoOM+HT48IE4e+aM9s21K1diaZ7nNKta+O7DR0Kac7/4HNQfnEliSeTgi3yA84x8FvS2B5L4OlBLLyWYEdUCDxYlhZgDN3JwniExnn3Ev+ksEbAofWI2ATr63BXYUuBLn4EGP/mM91DNyHsxvRL4CUNCISaNi9mTPBcugRgohn5XpxuxUv1Yi/m5hRgeGojVVXxnXG9wrHMWa7jZwfncLdkzDV1RBoE5QT2cQ1CMmmESwmhpiLnl4aXzZdZFMSdcDJth2XKSb89ja6BRe7OO/3bmRfu+UFUrsw7LXLSH0Gat2g6YyJq/CnPe24CPHEx54+nLf7gWKBaI4AhtTIBW3tUaorjst7Qtz4m9RS3XZHG15YcCqqkpbqBy+3Cm6k3fi8cHNKUIoTyzzfS7CbBsniFW01C92dsjtoS8vwbMTK7hBUBk1jVqAfIJxa9h3UMMebf29Smek5/wfiXNRF0rmWZ5pfU2fU1Zx4Br+Uzu3XXGyOBIqiAYGLvvwH71t1jr7C2eIXEAlLEBbWabst7Yl8Q4sSIS/LW2YhbTkSOHBVhiHzy4f191NB4VWsMpOU4Oa2Z+S+2DHiKMTfJ93sesi16BAK5eu6r+4bNBxT9iAv7srX83d2CX+hElN9OSp6hEsor4mmaa/tpCYSrhajMOLmohRXVRtWQipmQY0z4Qvg5EBGWKWqMLV6RvS1OOfgEUZQ51jKBJXvCEIDCCOJLGqqSVHFiZcNIwlemO9J4XhSJQQ6CvPyb37FEgAEHApJTD7OEDSz+VWZgGFXsm5WtR9NIaPCiZosEEwmNpKSbGxtUYQQIIw1cCMMngzNxsHDp0OK7duC4k19j4aFPPnWSQ35e2PUY+8wtKFNSA02EOtdaFv5JVCnUo15lMob1YAw8CMMF9ZWVJ/hgkRqK9gZDOYYIzZx/YRjFkw7fZOPd6Eup2fT2DrWnHZmJAQ3TDqpDbbnIPCHHJwU1iREO/TOkkDUPzRyj+DiGiKdJ60J4FeQZaE60/kNgkOCCEaWj0D8bXFy+qWUHjYXxsQp9VGr7DO9Sso6nC5+aePUqdXpkoJaNCBqqSapnX9Uq7NQ1N1zFUAuGeiZOa+20GryUDo9RdeqiNNPW2pj8FLol1aaTSOJVxaw4ESiaiDmb/6cO4mAxO3FKjMRMNI7RSBqqympKxEbLDyZ1R7mYjlWm9WEOJrC6KphuOHlQUXduo83zWak5acqp03UuT38WENTJrWGCuk/+7tISdtLYlojQfDKPRz7VwFU4waYQIPVDmx09r5IjBYpZHOxqnBhVGShfjofT9uSeWJ6jrVFIrFtO2WQKSEqhiriWBRWKhAR50SRBZnmbovU01N2MEtLDRO9Za3r9vn2IIhnggd4QI6mAYYN1V5FjQpCW2MQxlbzDoBG1FA6meDRrbLgAakmEgmeG9bALfGTNzMzLBJFaoKQfiDWO9/gHLMXU04tbt20rCNGxcX4ulZRC+IypKiNliTICQ6uyUJw+DFRI97aUlDyNqkEoRyTov/wpWC/eh9J0rTjjWN7RvKYi4F6LctlF/GV7w3k3T4+agwkWHNM+r8Z8SSH4/hqarTT8LjF4nJzEa3tRQl+YsibPWffrLqCjKNUPCKVk71nA2sUkQiQeF4rbsk4sXnkU172sQQWOj5PaIU3yBMKwiu5JvJ+ped8UmoWCSRm4OKkgYkeVREp7xl+crhGcbw4HfYW9ULCCJxcuI5+NYbukJvjzEsTyAGB6sdFGS7R3EuldBCmNtEy1Vb+Ua6vH8nmRU1Jov9LrPd17P+6FiYjWy2/dne0byTYMK7eG22Fb30E2sdhTWt8lvLO/RLmFnds+29oausaNDAyqzEC1Bw/2VD8SydeN1DQyqN9IUMItGFc+bG3H04J4Y7O2KjdWV2DE8Elev34qF5bXYQvqpb1D7aGGJ/UMB4fjC92gm6PzpsDHszPyszjLO8qn79yUxgBEkyD9uyfLSSoyOjml9kg8YyGHtcyG3dP5ZipM9z/kICpDzV5q40gPGFHRWBV3tTySlMO92U7HkyszE48yS8XVfnwYtkm5Iz5N61kjBjY/7DFaTs8uyYhq8jI6J+YkUlLwZenqUf3DWI4+0MDeXzKFN/S7xSl46eAjMLijP4xnU8LmKVKM/7QHF3myXAOQ13MzyOcFe86ChxzEhpVv4rDaj7VFsPHjoUKLPliVxx/MqLXjnny645fuTjcMmkjxHPDXYA7iyf9+e+PTTT9T8toQmxubDQq1OUWhOP/o2i/h3/jOTw8Mxoecyr2YM0hg15HQscQ5ArsnZUveWz0QDW00ONezMSuUMJy/wfjWKm/vspqzZYhpQZUxVswhpncZmnH7xWLx47ED0xmbM3bsXPSlhObRzNKKnNy58dTEePpqNM2deju2Orvizv/ib6BvsiX0HDsnz5Bc/fy/6errjxZMnJJV24+atWFpej3PnXo0rV68p14cFwKACJgVnO3tofn4x7t57ED/8wVtx69Ydrd/jx58XC4OGPnJQNAg4y2Bg/dVPfqLa4uTJF+Mn/99fx/7JCSGh3/v5h3Hg4J44fvxE/Ie//o/x49//Ubz38/fj5u07kp1jtm3JOSP+T750In71q8+iq8uIy2pQca8YdsHGQgJGgwDuGXIQyX5A8k+a2YuLTVkH4hjXq/yXgd/6ms4wgQFK5qK7W8htmhw0LmnE2pNtUzGO2H7m7Fnl+Re/uijfEp7tsaPHJJVBjqLXwyNOyVabtFAOEmu/8p+Wskq/qWQcFYq2UMKuaSwvS0wkNsgQFMQ8IIvFJTc/u3vEltGZJWZ2NXoM1HL+uxE9fTC3nbfRvAHIJWZEgsIKDMSahoGNdwcMIjcoeR3/vpkbXfrcTRasGuFmv/H5iSk8C3K7YhnSoLaPj89hvsilNEgRMy0NjzN53s5zqc45xfYEQXBmlHSu62qYeXh72GuR37HmOrmO851qABbLghhXwAb5PMonzueHG2WW9yE2VR1Ow14oX8XRzujqbujfqZuIj8QJfB9nMZlWTpf5v4SunCOLSSX2mq9JuXd5lTxlUAHt0GeZkcZqsGGCS33XoBFpABy5qnIheXnYg4k6EeQ8X4Bw1MRDyqW7u6lJz7/VOikfiBpIK99JtiQ/Nzw8pOHcg4cP9fssRvYo51j5bXGvi2XM9cBQYlAx2EujckuemVvrm3Hn9i0N144eOxo3bt2Iew/ux/fefiu++PJL9Sr+4Me/H7/66GPl2qdPvxSPHj3UABOJumPPvRC/+MWHMTIyKpDe7Tv34h4yTgw1M7aSNnJNnP+DfX3x4onj8s14eP9+fHnhQnT29Ma9RzOqSwrYRu5tWRtqIOoN5+nUr2LyJIjJoD4Pp3mmxMDyyeGeSBYwn3Gd1bWe2AMMyQpEUGdu5cKqq5kC5ZRK53maUvusJ+dqAfXI3xhIsG7J+WsWwDrrx6tOPnuAcToEFAAgUGwirlMvlzlYs8bW+3nYzr1BlYH9KBlDgK3c594eeXkxdGRSsrXVEdspD2a5J34u2/ApRVT5arEkBA5qZ0E0zaPziG+bVGQ75vGz/ymDihquOU9+/Mfr38ozUrFSqiZ5yrT9PN+Rlkl6QvBidb2lalBx3o+qHVCZs6pk2ObcWvdS+UACwexZ8+R1thgR7UyJ+nsx8FrMVr+mWW6WB+P9+NOsCcA5ro/Gxse0NquRDwBQ/URJunWrd9SA0Zl+ghq+ZX5o8G1KQZVcd4/VOlS3cfapPt2I4R3DiguLC4s6M/ft2691xvrjXJmYnNAdZ1/ZB8rs+AaAMYbnSI433D8jv2b4BfOSfJPv37h5Q/kRTC+8m8hLkagFTMUgDvAB78O5SbwqFgbXL0WSxUWBKWBXAOSGiaH6OfP1Z4OK33mK/ewN/qHvAIyKKsZEv0caozmxdSGipp76kGnwqyjqLkipPddhQYMGiaUKavzp5q/lKdjMBA8OA/tYmIZOcQxaRcOBlUUlsHwJXbG+YYQMJlcgGleZqs+lYex2bDU8KOC9ZAy1DdJuRUkyEgb7DxzQgcdGJ+GnIJ6RGTY0QntrgE7itQulo2ZzoyGTykIC6A5smjZJciM04eaGggnalDQPjp84oQRGenNtDRqSDprdRn2uKSEkOVVSmbI80mvPpoEOcLwokipMIb8mylu3PpfR6esyEq9mDY0HrqmaQVVUVqNXCWY2SPkeSXLRO2X9maVeAAAgAElEQVSgnk0wDTjSMNcFvJERFLk2TrfMjKj+un5rRFqz2411tG4YPFFkBg1laMadXULvgAaZW5xXYkBjUYOo6UcxNDigpIPhErdOuq+JCmbBsRbm5m2oqIMM08ek2Qmx3WhoXdAYIvkSogpzzWX7I/BVbATug4r3lN1ywtSjQ4VEGJkHDiFPwzdU+OI5gNF6Ia1kpJzJSt3zGixp/WQSX6iEkn4R46AtkatmkhpFmQRUg6+FaHaDXol5GUWnjE41FGroVUNGP3fL+dSX1q00fa3trwI0pYYUB1Lz3giEZHBwyOcArO43a1VrUJ4WNOAcJ4zsTg1G/i7013qi9x+bZDxBc03KcDubQ/HIeqd8KQal5Av/rUZuob7LVDuZMjIPBQ1L8p4aw94YqZuZcYmGLgWskI+SKaChbvYR945GQdGfX3j+hbh2/Zqky6pILEYSLC5enCEXN5Z1DsMJRLG9eDyMtDaxG0CwKUimq9lJ4kEhd/XqFTWKKdZkxMeeSx1mvsfPIz8nFHBJi3V4YMz3WLOgM/giVnGtPCuZxSZiniaikLC9LeQy719sHOIwP6PhIQW/DMcdF2pNUpAJqZvyUXx+Pq8KXDE5WmZxRkM6WaxGM/9ehoY82/JUIfYT4xkCu+mEoXWXhiL1Os0Bn+SqrO9a+4I/S/IC6jfP0tJNUHeJVaa3S6dXshtG20j+RXrbZqRwfSTGQmAmbV77iQZdSrcZWdOn9V1SVj29yMEMxd2pKcUSP/ccNsCoSSmxYhjABuSL/ybJ3c0wPrWy1UhNySiKe+nEJ31fKEeS+JTZ4fd9PtqDRbumzmlp7ObgM6+nzicV5ymfU9fK1ufeVKPlaQPV9lzlNw0dakjefh4Wyu63y3cYSPSb3oxeOUylTSPHVIijuZ5sP+5JZ7eR4BQA/PvSCvsWea4WCk/XVgNqeXpsxeTEzhhA431rS2cYKOyZhRUehDwqRtB4n5ttSnKxj2js98ucfk5SKd4voSEhiGlQUDRe8MBQg5z1vrElaUvWDo2a2gOcc9Z4p5HU7zWkhhjnWEO5k3yW1tZiaQkfFMswgCCkmEPCg3vtRr4HGvpvDdLMbuU+TSNTJF8Vs2rrWTPswm8CbX7u26EDB8RgBTgCw2N2fk5DDu+jTg1ad++aaBpxeiC/qeLORoLr0d3TG9PTM0YRa9DYiiMaNIktYRaM1vCK5XIUJ2W2SZOxZWJPPkSsJN/hXvA5PTg260tm4hnDQYKWFA1nFL8rJtPaqrZHyR6ZlWEgjotn7xdi4u7J3bFv72TMzExLumcQJHunzaMbPV3x4bUbv91Sjn3xo//iTPRd/8v4i/Pf9Ksn4k/+q/G486d/Gx//lq9+ds+eWJpfiEXpcG9krmoUJp9vYHBAA3dikYEN3Yot7A/ve5+vMuLNHMJIdGvHk+eQm9IwLq8P/pscSUPTrY1YXZqJ8R39cezArjhx+GBswzJYXo1rV6/HMfLkubmYXliI6zfuxpnTp2LXnv3xf/3Zv4uhnSNkF/H6G+fiF+++K03yifExNfkYENDcQ0aVPfbg/gMNzM+cPq3h2dTduxpQsdYZ5lPAs5bvTt3XZwVA8OXFr/T8Tpw4EX/zNz+LkydPxGD/gEywv/fdc/HwwYO4dOlKvP3WOb0er3PixMno6evTEGDq7v24fO26maPqrHmANjI8qP2BlBVNQ3JISUGIcWWjTQZD/nKzjgWoJktbbCo9cJ+llnAlnsvweWFR9YX9pJAC9MCd4ehLL70Yly5fipmZeeUbamLpENiO06dP67VopEpGVHrYIZN44hfPWwN04Zs8LNSAm+vrNGOM11lZYd/1q74ibze4xe/B/yQzlvIdrv38PtQGMFzYV6Dd6yyqswGmss96s9T4JecLqxqMwuCq4aARQM53xCJYXdeglEYVcYRrn52fVyOpiVymscSZKGCDY5CZazSaOj3Yz3PY0nsN1SGV6/C5lH82vW0SUZxGza6tDA5TbZTPpX5f96KZx7aG9Ab9lEG0wSxl8u1cyzm4PBtSflLrLWuyVq7v95bPnO65EeFCIvf361nB9mU/SzZYksxbMTSMZ0qHmIA0iu1Lw/P3dbkEaEn6mCmYprLUaHmN9gp7XLpGuXlqtVfcJwetmlZxhLpBMqqW3BFQSrNU30dJyiKZImQ1aGRM1oe0FshzyBU5L11Xe4BEPsYgzMMIr5XKX/g3oa+zQW9ZNvvL8CXWTJpFF7L61ZdPR39vQ0OCPbt3e8C3sqyYyntcv3kjFpcX48x3Xo7PLnyuocoPf++H8fmnn2tf4w8z82hazUUk6A4cPBzvv/9hHDp0NB5Oz+o83UIOLaU3iVmra2bCkVMszs8J3PD8sWNx7OgRKTlc/PpSXL89pXvkQZljAJ9LHpbpe1LsRSHIs6bjZ8iL+ZzGmHmgYyBMrUFyJ8sT24ci2UliOhCvQJEX+I5nhbSzhyGWEvfrajCQXmz1PZ4ta1wMTwF7zAgpGRvVpimZJPYWTVjl7VaSGNkxpHsv1ihDL+oC1nR5kGxzRuFL5j2ruIsxc5qNO+cnL1yOtfVN+Wd1dHQpX+ZaAbgVeFfspGTiO655bZqh4OS6bR7R/LuAb7Uf2igTTWmvZsxM+bwchtRwxLlL69AX4ChBWaqf2oCW9VOKP8WsyF+u4UZ7fq4415SkygKhTiU13F1H+njKwXX7IIN4RQM+Y3udZ83ryGtovy/NC0sORuuTOcbU4JO4U6x6hhB9PR7IWkq9R7FBZ1P2c6pe5XwRI7ZBrWemJ+uLNUI8Lzk95XvJdlNkkySdBy6SxM7PxvUM9A/q36k7FUOiQ0BqKJ6sKQ3RxfyoWtLSe1wHfUhuoPoHOezXuoYlCdBmZcVm2aNjGgcDsqg+A4x4ZCWJybUn6U+yl6lLOSNL+onnqhg/OKDzTzXwM+mn3zJbfvbj/+TvwNiap7JGsqWWXyZOTfmHMs5TgyYns4USTc1LTVrTeJvJHkGGpMJG2m4yEtg21ykAQwWeGtGiuCIFhQb3hpA383Oz0lIlqTh5EjTCtGQDKDBBthH0pqbuilWhhkBHRP+QUTZqrqHxNjisCShBiU0+MzujjU86dejgYUk/QRnji8K2UMV8DhIKKFZGxd5TUq5hTTYI0cykIUFBI7PuiYm4ffeO0FJE3ZIAYVIqs7eUVUJaSoVH3iuuqTR+aRxQ3JB4UESqqdgRmbjbmJygxc8omaI5xvS1r0f/TQFDYUPyV0FcDZyU7tLASdrZ9ipQwzk194yIMYKuEmBRqfU9J4ugbkgW+Xf5ZkCr6+uLO3zu4eHU0SVoG5VP4k/RxvBhi2bJ5maMSO7Lkg3TM4+iC2ZIZ6fMESki74O4436RPCBfA41NiWyXkks+PwkWxaIajd3d+nk3r7ulY8u1qfihOTQ9rfuNWrIQTtnULjaCWBfd3THXZrTN/esfNIKdhg2fhYSOYnVy924hjzILa2vuOCnzcMt0bv09EYhKwhIVq0QoG0dGSpX2raneloXJhnrR4CUT5CS+fsdIlsc9LvRaGpzQBKOBkMjhfG9+3mgbN6VKt7YounzfdNFk4Oj6s5DIRnkVXlrHOewgsdP3lZi6CedfTS8OCm2ZGbY0WJtU2GZS87ieplkcoIstS+NE3NrBGq5kQs16FHsLllYWkfyMBmIUbWmqTbNMxUqYNUESIdkymRyasi+UowpONx9ootPkAjEMkookgQEAe6IaDUiZse+QZmJ/IyNGfDhw4EB8iaTE3LzQOTaK9t7lAVejzUbc1lgubx7kOebmGPZaK7xksFgfGH0NotuqIr1TRRqvJb1sIf68l7lmF6Os3z41kFysulFC/II2akYGEgPbsXfPZBPJyXvVoEIFiRgPblLwJ4gPEOF179mfJGwUZnpOOVDzkNva98SdGlQI2Y9UXH+fWWSJytMZQmMSJssw3hzb6VFRRVOa26XMgptoaP+jwet4p0ZByl+Vj5DLbWtNVyPSw14jYviqoXX9rtBli8hckZSXVrS1eG3KaR8C0ZOTpSO0ZLcH7mgiq7BPtpLXnxtIdQ7wGpZ+MuKQ96aY5fm4WWCaOEm3G6zIbHmt67NyZud+5bOwBnluxLQymXQsstRTMSrcBC59+SzMUo7DRb2b/zVIr6FF+/5vT26+aVDx5KCjGgY1pHlagvTNr7Wldcw1kZTDQnCjBBSkGzCsW8k/4u0hvwevbw2gtO9oZri41IBVcctSWhomdWzF2MhA7IB23d0Zg/2Dcfnq9VheRzqnEd39/dHXO6BYQfx0ccF+bMT2xrb2I/FfcSsllfCLeDQzawZEF3HHawqG6eTkHq0dEFVC88I4knShafcYSpJBUdTgT8HgkcHLgf0HdQ8ePnoYO0aGNcDns6JzT/Fd5nycj0KxsoYErli3R8aATVe5bxtCE3sPsIYYWJL/EOvYL+Ojo/Kr4LxneEgsAEGqBkDmeeRYFQtgj2kvIYW2umYkOK87NOIByfTD2Lt3v6Q4yeeQ2+F1WLdTU1MCfgDiYB2ULIjQcD1uMGnYgKl45gTsPxeMNcR3Ifn8c883GQK8F8MiDffQ6BZLw9IqdZZSYFazkj/NbvFgH5bTjh2YdXZJDoTCkM9HjvpgdTWuP3Cu8e2+9sW/+rf/R/zPPxyPmP4g/vv/+l/G//hrw4q34n//6f8U/82LPbFy5afxr//Ffxv/25Vv9+r81IHRnTHM4HhpVZ47GoTRrMXTAabO0JC839gH0hgvSTatgS3F3vIw0jCrkO65piu/4U9Lnxk57TN3M3q7keXcjt1jgzHSG3H6+WMx0tsbCzPzOjd6BoeEIl6N7bh3/0EcOnQkzrzyevz5X/wkthrd0gz/3pvfi3d/9rPApHxibCz27T8Q5z/5VE2rY0ePao1duXJFcfPM6TNx+/atuHfvntYUAzti9IULF6K3bzAO7NsbP3//ozj+wlF95suXrsYPvv9W3Lp9J+7euRP/+Z/8Sbz33ns6/zDcvnXjRizMz6r5v7K2Lk35H//onZhbXIi7d6diHZQvsUdSuY6VrAXuAch4ewB4SMd11vnA92xkvdkE0yjOd4RM64m716/faKLUidv8Pmv22LGjeo4w9Tj7BZJIzXe8b148cSI+u/CFpFN4HtK17qUx26PmKjGIc0VsyuVlDR7JB9H/rtxPTe5k0IhprAGg2Uz8LHUG723ZI8sVit3Q1vQpCR3yz5KvZW+bIdCIAYzaMW1OHzViEfsNdCixGGCCB62wJEE8G/hSsV5s6w5Yz4AJMNo1gMED4zH5jNDE5ixQX1HNXOTokkmUXhsyXFVz20CB3r4eNT0lQ8d92LS8ls7KlIVs5grZFK+GmM4sctZk73EmFxK2YgoDYZka5yDIjTwn+9X8Zd3wM2ZJtLOtH5dAdZ5n9mPllNSMfFbuA3mVAYebYuAR56mLNZxNFhSDtN6+btdjeARud8Tc3IINiPElyfvSUqPfjs7ws6+GbfM6mqjuZFjz0bIGYFDKe0q6iYFLSh96AO3PyWdgbZOXc+81cCa+46+WPhTEe/I81jDPiCG+/i6PDYzEXS+yv1grzsGmmt6MBqYgS0xjETCa14/Zq1ZMYI0AmpSsZwNfpZk499p3orMB4G1JzXhiERnTc8eeE+DxwpcXYnr2kQarn37+udbe29/7fnz80ceBp8LZl8/G4uK8PHQm9+yNfXv3xUcf/yp2TeyJ23enohcmoeRSc0C4vak9wO0DfCBpJNX+q3Fg/974ztmXY3V9M9794EMZn9NI1eA4QVCsUdYx/zOo0EOuNZlXG4BVDVCevWScYK0sLOgZFeOXe0IMIIaUtKuBAJbsrppP7O0CIOXQo2QTvcJtmlz1sPZD1vXEDkkxq57x2cznpiawCTGSeuR31ICWSWOwQc5lmXFLPiMh5eY6ewYEO8BLGz6TPxEfWS9C4G9ZdeDRzLzktlynwt5gSOY1YAZEyrum/0bz+vN39NmaJtutwUJrX9cmqHO7XU6qlJ88sC5VAEse1c+3JhXag/pP9xWytdAGQvTPPv67fj//Wuu1ajThXkUV4OVpSm/IYOKSp5YyQRX1KU+m2qK8JlvzkeZws0CFFVtrGFu5VhNEmb0wx0jHONWbxEHyMQH60l9F/Y1UqshnQw5nMJ3lx2E5qv5Mhgbr3OwhewByH4gTrHXiC3tq795JMSvEEiZ/b3SlB1MjpdRWJWnO2ScwR7eZXRWjGY4Ts9k7/IwYH5yvQ8MC3BHD6CWS47OffW8bAncSfxiWIiVHHNJgrJth3A7n/Ak6K4WDI0eONPszxD4DcmDSDyuvl/n4s0HFt0+Un/3kP487sHPZdMEKWJUc+c800apErZqbIFwSgaqgIk07+zTUBF/UKNzrGSAkY6Am/9CgSlObBNAT+/U4ePCACihQggwLCKSnT50WC+LyZdB93fKo4PVu3rxluhaI7c3NGJ8Y00CBpnmha6cfWt7pyNEjCmQUyPhHgLDCENnFrxtcfF706ZCEQiJi9+5dOUSxtEDRZUEzYcbHvXk0Mx2Tu3YpWSDp1fQWKYaFBQUeEEQMRygISH4owMtngvfm30DqkbQzjIHSzOeXWaVYAw0FTjTPhXRBQ7KXCXN3ypyAHjF1n8Yh11VFiNEM5SNi9E/d83bfEQKsG3dO1rmumnCr4EiWjdGGLVQDP03g5TmT8CGFxTAD8AT6jzQaSJZ3opNK8rmyKhQ4TX/uF40VMhOmzQvzCzpk5FeSyAlu8J7JvUaZiv5pBA1rjULEjSU0xI2WJJkiaJMw0Tjm4Ll3/77XdSJquNaSpJFhVqJwfD/Ckja9vUKxr66hHz7q+940ucOcG/NDo6+KgunhQOqvJ0OhNahIUE8TxWwtTbFZGNyRgOX11wBLPhapfy90QDaZoGZz3dznOow9TPQBb9mWNL3jWWH6lL4S0riXcaDpvkIDZOHmgsZDkMcHFaZ3m+VRtEw3wjUkMdykKf3E/TB60K8nBE0yH5ah3SdCL9MtB8hCgLSgIE0ZJg13UmpKBmnZiFTMKbQtnhSJFC6kdPnFcC0k4dxLhoZN1BsvkEi1lbXV4H88k3oWnR0uYFlTFKoMIV4/d06I4Q8//EAX7cIY0+JFF0X9A9no7pHcDMMOCl/2tBuTDRVVrPOhQSPCSHaE5kAGZnkpJsYnjJh8eF9SUcROxZ006GK/lQQHw1HknCQHhxRDIjtpMGG8W/RX9iCvQfPWDCUnccSYBw8fRXeXDdL47CQ7onVv23jSA003gmlmoP9JTEdWwsmkdYGFxkyquKj7bbrLao5SqCa6Tqi3RH0VnZzveTC7bdosa3MDE+9hrX0QszVcQ8KNgWQBc3hvDweIiWWA6VhGoTo3N6uhpVCkxAz+jjSVWEmWc5DXyOZWys35XhADWC+grry3LFXIeqzGg5Z/Ikj5DGJkbWxaRqt/MG7evimqb+1hronn72Tc7Br2HowKNaNSUophAzrEJSvlYYplPSRtlYWnzqU0p6/BHZIm3C9kCNUISPZAxf56/q1zPg1CZehu9H1JdtRwooaEXH8NR5/Mbr5puMD3q/godJcLvF+XhGqWZ+1QsvY3Agne36/nBdKQIZT8Usg9OMs1BPSXm4duqnhghyTUoNgGNZjl+zofkgFmdtJ2jAwNxnBfrwpkGfpO3Y9Hs0vRSREvKZZhmVW3I8F4z/7ePp3DNiPdUpMPbXj2DkNz7f8uF33lB4PXBHuNJnoNEmTIq7O2ISQ5hTWMQwYQNFiILQwSODdBcsrTRUyqvugfwD8qC7pt9oClfDzAs9wPkjecjyCzZKBJ7EtvAj4TscXMA+TmPNhkrdEcYO+L1dMJo7FbEipQ2A0wdGwRmjARhTYCn8rnYVCBEK/4H2A0nA3Teg/e00AIGAvOIWttsV85e2lMufEJAw5d6h7HrJQ95PMzWHj9tdd1XylmkdspDx9+j5jcREom8lvDGocO7XWde8Sy2I4D+/dr/dy9ezsOHzwov4KBoQHlN5/cvR8r2bh8cl889b//xb+JG//LW7Gn/vHXhhWtIUX9yBf/9rtx5l99q1fXD/V2dcULO3fE8uJqzC0gLbCgdSGZBJmH0uy1/JCZsWYuFpqS4ptzzDj5bCDlvoT5rNiZPjk8I9aGcpFE5iObBrnwyL7hGOjaijMvPBcHd0+STMTdu/fjwaOZ6GJYBkPh/v04duxYHH/pTPzp//3nsby2GQPDI3HmzJl472/fjY2NVfkVTe7ZJ3+H7Y6OOHTgoJC21nXuEpAAs1rW3q7du7W/+LeRHaNqGJ59+UxcvHgxujp74uzLp+P8+fNCMz733HPx8/fej0MH92lPXbp8WXHlD//g9+Pd934RpFBvvvVW/L9/+ROd5WfOnpb8FI0Hmqw0whaXl9RsWFldFmPjypXLyQDalpwOW4MmJMwkBv0wOjQAZo1J+okm2ZakJWlQfHHhiwSSEJ9SX3w74vDhQ8pLGJQBGGNvyUspUek0+gEo8PkNFkOj2yh6hic/+49/qxyA/9GApYlC7BBoKY23JY+WTXku3HWhB+zUVgyHvVed53FWav9pz7TyVjURkeRNQE01+Au9ymvQzHF+tKKhBO91+NBh1V8yveWMJO/sAoxgJo9rSUugaiCmM9d+EpJsyWYe5x8xWsx2DStg27mhTR3lAUoxC5zTFlsRhkarkbatRr/kvRLxXo0+y5c4b1ZOkGbCHn6mJBg5OfG3jUVp1oTBNiXLZACBARDF8pDEY0reia0pFjjSvFx7b4Lnkm2cZ7OeJ/WB5KRWNbTCo3EVLx/Qt8oD7a9ErrhjdERyx0gcMUgmLpBnwoAr0EsxmhUXU56ID2h/iALAafJvQEQGUeVcMNR7e5pgFCGns29KXcx7WJqoYcYszzONcEuil/xakm4aUsNM8hCG7wng1yYZxn9TG7CHWQ8oKqBrz+9qcJU+SgX0QMaPMxEAmliZ8sxwnc16hz33/e+/GcuLMzHzcFpydOQegBSPHTlsYAj+l1cvx/PPPx+//PgjsY7e+cGP4r1339Ng5DuvvKxhKOfg3n37YmJid3zyyWcaVBCbyRnuTz+KDlifS4uKuOSM1MoA/ZA9Yn0CSJifnYuxnTviwOGj8fmXX7mZn2bCque2/Dnd0Pegp/oueHkK6JgMFAZA9hxMH8Y8a2uPMkTwIINn4oE+N1Ay0yW9mP5qxU5UOpX1djErXFsaqa96ElAZ75vNWjWSqXc7O5SHM0hnLwm4hTKGch6DFvCqWV1j+Ga0OzkItY3WgJiD62IzGRyUa5FhPB5djQ79XsVeZBGBAqn1IRaBewJRfhRJCSAPd48owXhpAF3N+CfT1W87qGA/VX5cQKKKvY8NHJLhKZ+ZrFudP7fygQx7+Y0aSrSa/5VDVe3CD7YGJA6bBfbgOZG7ul7Msz8ZbgX00J81Zm3NQJosk8rxW/JZZk3U4EyN+lQT0X3I3kyxyMTsZqgNAC/ZZPwcz1ngPtU1XkuWNLNEMjljvTfrir2gwfO682P+G3Aha2d8YiKZN+yZTTEmHY89YOdM5/XF8CVPHRhU7Vl+jc6DyqPIPmvkTbxG+XWJ8ZZKApzFNXBgTy0tLMbAQJ/ObHqB7G16NIMjQ4qJ7DP6eyjUUMvxM6+99mp8+OEvFQMBtJXZNmcvZ4PqxmeDim+fKD/7yX8ed2DnitGcfNGkKl30QjRrgpmNBZJ/DgAKXBpgJYFDslieABU9a5BBkwizx0IgUyxXk8LUKU/F+XmKcprZC/NzsbxqTVYScevIu8nMNJ9AwjVwOCrBk3HQtpJz/tFGWhSum2IngLCS8ayaF25msPllspNyMgSZXbutie5GsQsBUIdKbkkOE/FKslJsESXyaoQuxdzcfOzbty8ePHiYhrcYZi4LFc294zWFIE7dVF4bejHXgS6dUWkbKhAtsWS0LsmGmAwrNGWgLDO9RSfYyTaficY/99B0Zwdrfl9UfVHOTKfkAztJpogwwtZIQherkshCYiSTNg6QugZetYm2SLQVz1IHmoZZNK8bagwSOHeNT1haACQHSXhnZ4yOIvHVHw+mbZ6HQsT2NrTXdaNpJGfTFQ0OxkQD0OwR8qnRiKXVZSV33A8ZmT7mj2I6J9fOmuGZCDWQ6O76TE4GTOUjKeV+0ATk2YjunTTu2hesNZ4h6HiZQ/Me8sYwmtsySN7vGhTksKLZsE9jMSOZSsYoaRNNsEOa7opWmsbnuVeEYMq/+12coRjkkM9azzdNgzP08Gx0PW2U0F+LSm3Jjl85kaRC2FZJ5lTCUgUtI2AlCBRqpTmeiKQa/Om6M5kANe7hxm+Ki3xOMxsqqSkqcRWtzddou+4W4ssJD8aHQryCcpCcQYeSAvYKxRB7vZgVNBBBFMsMPtH1mKpr3+QAEwSgzbf88f1vjhEk7GoGprqW0EzLNpAVQpt1jPcM5th8H/105GtgXmHcuHOnYgxrlcIRlpgbwyFfFaHyNBQDOQUq1sNJYh/rdm7BHgw0sPk9NMZpJpbec2kX06hoxpIcVoHMVI7e8DBhZMRIR1Nn3ZwHAUJ84JqFsE0Jviq2iU2OgY8jdrwZnNir0SVTUZ8zherir1WsK56JcWNJOfa2PDMUz9MwN+UnSsaN12+XdNOgqTZiYKhrJh33hmelRkOvpZj83ln8IC+Xw8da3xSpJIoYvaJxq2Z30oT9d38QoxnLKNoxkFhOMg3bTJIZuVbtHWIWlWJRIrPKMNMI722dVxTOksxJryAX0C4WvZ5cSGjgwuAMevQaw+Ax3S9YaiqwsrgX8yJ1VNXskZ6qz1SjuYox4rjiz+gLbx9CtBc637STv2lo4ZjVGlD8pp/7ptemEU9eMLpjR3NItjDHHnABoeFDpxkNLD/us+UmOmN8bDxu3rqpwt5DTVu3GoTQQonuHB4SAq+nsyt27hyJWzdvxQJ6yJyVPf3RNzCkhg5nDA0WiguGEcQB0NZ1Zi4sLUmihjegGeGBt/dvyb6mDWYAACAASURBVFSw/7kPNNRLdqf8vfhZ3h+WB/uStUnzhfiGt43lWZLV0QfbkcYQ+7Ez5REb2nPymkl2AnuKs5TYwzkP083oaw/puS4GFaxfkGceCJhtQXwxkCGbmykhQUzje9Yidxyl4aSGCewuZDqX8aawNBcgAEs6OIfR66o56GfA56p7UHG2BoTeK5YDKcNeGerC6oSmv2p5F+5xrS+K1JIPKCNPNawUv0HY+tzw4MJnaDWy3BzrVBN7167x+OzTz9T0npl9JPPkzsH+OH/j1m861J7ybyfiv/vT/zX+h7eHW//WHFb8+pAi7n0Q//q//Jfxb34LRgUvfGL3RKzOL+re83xpUqnZkzGyingKXA8qjNL2PYIdZ/1zDaAyT9bwGmmezEI4Z/R6zaYt/7YVDfLCxla8eGxfjA52R+823i/71DhnjXx0/tPoHxqJpbV1DX1Awp978634P//0z2JhZSsGR4bj9Okz8dFHv1TjCUDP6NhEXPz6a8XIgwf2CUXLcIK4iv8D8ZRGP/kaz/eLL7+ON944F198+VX09Har0X/hwhcCIQEiunLpsrymDh08FO+//34cPnxENcjf/OzdeOXs6ejr64lf/vLjeOONVwWu+fDDj+JHP3onfvnxr9TALFAHmSQMQIbbDFwufvVVni/OK3X2bGzGgf0H1PyU/BJDgK5qKpuZx++yEtHQp8kmg/MuwAI9RmDm2WF5I8tMGIji58azEQAopYLUmN2ybBQgMM4UWCdI5zCAxFjbz9zNRzV9miayLVasGo+NhjTyqW24lpJTa0mllYF2sYs9IFYunxIcNHZYg3xR1yGfR75taUwjXok7bv4u6WfNAChvN4OvxM5sNDyUlfxQt3JzXRf3qrMhc2OG13w2N0rNBJfsXb+97LjHfAEUoC51EzBBP2IzZj6P5xnMtPRBEtJa8jYt9K7OnRxYFKirwAOukRjmYpoOEMSeQwLyJCNGZ3Gy1+UbmKbmMjNP1YGKw9qjbazsGijQ4BX4IesFxUoGw5lnolRg0FOnwDej42OK+V9fvqR4yb/B1qO+4TPItFZrqIYxmyHx4DYjXKOUnK8D4rLXGOC+zPXwb1NH1z9jto1lncyoYEjlhqj6D+SBNJVTprQGORXLWdPyaUsfQnIgyUKJmeGgJIBSmmvzOcys8R6zX4JlhIlvvA/3oMx1K182s9Hs53Ovvxqri3PK0/ft3at18/DBfZ33x184HutrK+pbzM3PxoUvLojh8/23fxAffvihQCPnzr0eX371lYYnR44cjbGxCTHDRkfH5SF0+9bteDQ/3xxc8kGqPuF1NVxOuUYBErjetfWYnplprlvWn/LmbgPQSo65JJ2obReXVvK89TrxvXUDXowWcsYOy1+1SxDVa7GWDPzwMzcwzhKBqtuT7Vt1Z7F3K25pDTxxGpYvnHLoBP85rnk/llRrARglp9SJP0xvrCyRf3ULWOKcFt8xDzOJEwIuZD1Z18RgmTqLmAKglKE3xbtiQA5oHYkeN7lWZdz0aWr5MPCeJelW+S1/toNzmnV4G0OqgELVY6imfYF5WuCM31gwP5ajq9bPOqxevxnDijH5DQAh/V4ywkqazXHL66R54Lc9v5KdM/PCQ0zHrhwgtyk+tN+/Vg2R97FksjSsyl5HvhZgBJtUm2nSlKZNv0Mup1icxBPWhVRFtpEYXG72yHhO5J6sVdY3e/7EieOxubEaCwuzqlVhOJO3MmgsBRPySvY9tSTnKPX1BuwhpNGVV/boZ1nZYoql0gj/Rr2t/Lrbvje93fjm0StcFringHXIy1v6FT/GGQH21vFTESANmc1QvkK+znDlypWrGsihFcKwlwEMTS5ej3Pz2aDit0zHn/34P/07sIukIU2lZcSlqbclbNTcyAalmuxMHFOzTWZg2YgTuqK0PkUbtba/zBiXl0y7atPUA6GGhAEJM4k4oXhzDXqUE2gMZWggEoBgOXCAQNGmob//4P4YgDY+dU8TRhmgadK6rqEE70kxTYLMJBRZp+GhYSFraSzwGdn0FP7WjSaoImGArMFYsxFdGnQ3bt5UsOjvw/B7NQYG+9RcJJEsTeSJXbuku0vyTkELfZbOpRAnafZljdnJ5oCHz8L7875KMlIehftIYmDT1y0FVhI5ihZRM3t704zW0j3Sq+7tUYJJsKthh/T2UtrDDQbLHLQ3nKW3moWokreS+gAxv0HB6szPSWvLDJifJTEsyaxCEJkO6AYX1wxzRYjijTUVmzt2jJiihj7+MtrvFEfkJB2xzoAEGQohkCQqHzuGhvVsZOAFBbyrM2j+LCwveZ3SsEjpAQ5UrothESgtpCk42VgLvSnfwM846be3gQ457tPmlpDsGOiZoQKahYbKqtZJrSFM0s3csMHuY1mXLtqJQtFeqxHoAVlLm7V96OC8wlfjg7j8JGpwofSnRT14WsaQGvx+pZb/RQ0uatj4d0UjnpuYBak3W4OYStraE6FCc5TJnqQjikKRiFSt6UycKRppoj0GA/Gnbl6WG1U5DVBMsRZld4+fdQ3DKhlrR241XySHNyWLpEY/KKNEsblpZV8YCh4h78Rs4Rk1hJ7jmUuBS0MG+3CoaSBq57wKFArjYiioUNy08TrXyzAEJIh12EuGYVmfjfVMYVWJvhrP2ThirfLVpP4jCSB5PCP3SVTEWkp0GBdJTCO2NCR/taHmIv+uZk1J23R0OLaRpCU6CQNSvF4oREvGyPR7xDg84DJTAaprt+4LMcZ61lmcpkxIc4CVD+HJkUWdE2pSJ7OI1zdLx8UxA00aslWAE0d4PqwPKK2syWq668xIxp+Ki5Q1Fp09v8/5BcOMBrEBU2YErdPITf1S1hPrgddyUy5U4LI2Stpubn7RuqJNw2sXaL7ONhmnTOo1kJGcxrD0zYuNp7jbZKWZpcL65vkS22qdcM9h1pAcU4zWs1EiXMMDisON8sRw06MGFRNj4xrygzbkd0A0WmrOwxWZcQvk4yYN+0r7Yct7DUQSCTPosvahRHPPtcO4viGgPDmAePJ3v82w46kv3YEhJoI2Ed85eza++uprna86j5A6WFu1jBmN8j6Yh3yuzcA/hrVDk1Cfe3tbjUZpQCcaj9dQc3ubQecahAE1ZGk+zs48itnZeSEeO7vxgdgdUxhyLiNZ6AEROQFnHmd6Na04R8hBaKhzvhjNngjgvI9uujAQe9Q0eq/mCs9jbGyH4l9ppCvPYhiQ5wRnPkAQPsfG5rrXeSdN5hWd+aAiGTZKQkbxo9e3NiU2KKhAkyk25aCCJiKxgDypCmgPyuy7pQHpXMmz9Og8d/GHeWVDg1I+E01ghipIcLFnbABerByMQz0gleeLhvtoBPtEIOZY/smX22T8pf4wuSLAjWp8MkgFMerX8bADT4NiEtEkkgxcSqARN3pSvs05U8of0XhIDyjHDGLEeozvmojRnTvizh1LQAqNvb0Ri41GXLn/8O86Wp/y708bVnwSP713In70os8Hff09hxT86qGxndG/FTGHiXl63kjiBLBLSuXwDIw4N4OE/LtkQThbPMRMCZpkMhYTTWywYlam1A3SA+S+Pd2dMffwnvwphrs7Ys/4iAxp90zukh743XsPY2FpNVbXt2Pq3t3oH+iNk2fOxk9++rPYQOun0R3Pv3A8Ln39lfYNDYMdO0bjQUpvDg72yrPh5vXrGtYhi0STmvMJ+aeRkZ1x5dqNGB4ZjqGhET23HTt3aAh36dLV2L9/j2Tdfv6LX8Sbb35XQIYLX34Vr73ycty+czce3H8YP/zBm/HBBx8qdsLuuPfgofbE5StXZdDNwHh9w/sB9D6IZxDT+FhpAK/43tv0vhrow99mRHuHPcZwuBsvnAZ5qfcXA1DilL2/nJfaB4a8g/2EvC3DJ5i+1n+vwR4DF5oYxH6YkjSO+QLMc+rUS2IU3bhxQ/GIz0EOz57gnPHP28y2agJ5BmRTksYMTVN8qZSTJcO1zkIPKu0RUOwchxniEfUH8kyWSGRL81n4HYHQ8ho1ROtoqEagIcP7w4pu1khbG/IxJI4NijlmiVPlemJJrSp3HxoZjqn793TficfILyKb11rbePpwPcRuWMacj853Wk1FN9Y5n6uJTXOJHI8veQIluKzkZpuN2fJLSCnWkjCiQd/eiBRCuw0L5AGEfd5gvLopbO+85jAihxt8NufHWcNpPEi+beAE90W+M5JCacTuiQn590nWK70Fd09OKoZeu35d95jr9ADO8jt11BdoRxKvQliXV6VrDcuWkseYBSipVtXlBjI1axwD8vN1GXZbCpS8m6KPRqGb2m6GV76jmJ7Dqno+nNXkVrAZuAYxh8hlk33Ou1Mrm6G3lNJ11Gxm5xik4iZ9AU9k3CvJS3IkA1P4PH/0Bz+Ou7duKKf2QHQz7ty6FS+88Lz2FsM/JOKGBwcly3b50qX43htvxrvvviup4nd+/E589vln8Wh6Jg4fPaYBxcfnz4tZsbS0Etdv3BT4Tr4zW1vqEchzs9EpKWxKSzfeAUt2xdDAkNbv3XvUuGZLF/NQDf2sb4rBQMynHiFlaPkVWt5TeXUyS8vInX1ZigUleWZpyHwmGly61q0hhdaccpLWHtIz09luYIGHVa2jjd/nM5XEkPL4HMay9wE0FnjHgCdB4zSc6ekxkp3P29fbo1yC/IPnr1ylAFU615zbSuptjRjSp3sEmEfgFq4617HydP6jea01sPBGrVy2YoU+TX6m9vq4fV8266X88PXf7bWfFQ5+Ped+Mpf+pkSj/efae23tP1/f/8b8OwFV/hz+zSdfqz39NzDFkr4+v1wXyeOHPkvGg2avIIe5WkfpXeJ+SQskpFox4yavjWQ3e4G8v1g8BgIiqes9WvuW1yE+syaJKwCSLKXtvJDfqaEZjMh9+/ZER4NhG/Wdz7qlxZWmMggPVgyIZSsIVM1EDlmydSwcecNkrc41ckbRM/K5tRHzy4sxvGOnapSeLnI7D8R53lzP/Xv3xWIbhiUU24rJDDg5M3kODPSpRYgLANE4t6Uesgr4cSWGR4bUSzVoJJ4NKr5pkzz7/j/fOzCO8SODBRpr2TzRJBXkHl3kNiMqodoyWCsp6DbtjkOkqb2pSWKvCgbQrLxO30CfkgoFQJpr0m8Dvbuo91aDbmsr9kzuEWKBCSNoVJJZkikOWjwrOLTOnD2rAxzNYRI1DDI5VNBGJ6ggaUASzjVV45rkgoP8xo2bLlwwpJmbbxbYOiBiO/bv26+mEbq3JP18H71LSQ+tb8XevZD1ja4hQN65e1uNCA5UayV66IOG7tzMjAoKDn/uEYk3hymSVmpOdDZUOFDUE4CglVnayLTmCso8CxItG0Zaa9uGbkmjS/QiQdEGYm6I8r7lF1ANVe5fJZ0t1IObqRw21WAxndSIkko0ioliDducYtPgTU1FJ5Oms4vlkUZ3sCqWlxZic31dyRKDHA4e7jPXsiLpsV5ROu/em9LaALnUQZNmx07dOxqZNP+6+/ri0dyMhhxusak1rveS0VIHRTm6k15TQvtz2AmhmYZd+jfkZ5wU6HBNtCnNJnsGcE3dWkMcGEj1cOgiz8VByIHTNLXN5ML7wllLDSpYf6WDq/vtkz/1oLNRmL/TnsA5kbC/A1/tvg+tRKFFKSgKugcKqcGfKKZCiyYR4tcCVfv7VsEh+mzKhXhv5N1OVEb7a0lUJZEyeu/8/Bq4bbtpKzNIpJ+K9fHYVTgjcsHroWM7GoX7zkCrOlhVZPFzTxtU0FRmLbDGrEnqfcO7aCAo02wkyozoejQ3K6ox64UGAd4WamqM2PhRQ9xEN/IzvK70UJNtUMPEGkCArF5mXy/b/6QSeoox4gTNNw3PemkYmmlRCW410CmISNLK6Hp9hZ93kSydTGJErk1JmaVkB8NfCpHFBejjHm5UMTK5e5fQRxReoL6XVlZjaMiyLpL4aUNMcw9Z3+0NZpr+SEUgIaLCQg+gDWX0NEZFJmMa8gg9jUeRZQ80ZMxGIM0KBgTIwIl0weByc0MeQ+wXYrVml1CzJW3AcNvNM5gBZvVEPudEo3V2Rb8GURj4ppG1tErTwFRMMjdKi1Wnplsih2mWiJm1vKrXL9k70XpBrkkKwrJr3g8UQjSQaT5ZcoCGmeLElq8pb1miK92k4fOY6ZUyZxsbgRyBE1EXAi56sqDmPO6kKDSTwh4sJTOxIdaA2GTp1VPsGH6I6ybOyyxe8lyZwGu/wBjysK7oz62h6a8XLL8p43lacdW+lv6+gwruoc16O2ITE0aAE9KwXtVe516zlmEVyuCd57BzR8zMzMbhQ4eEvmaPcG/E/hOTwjkNa56mBvkOedDo6IhkfzDNXF5ZkmY+Nx7oxvAO0JPWeYe6jak3YAjOZhdJZunxbGVsCchgEYTwqvSoxT5NyUlyFfb9w4cP3OyRoSWvw9CyI8bHd8ba2orAD/53Nz+hffOzSFBQqDOcYo+CHF9cQp7FSGJYIZLGWwVJZr8F7hP3h3VCkS4kazJNWecMAYibNFO5TiR0iEncd66X9VGUczVpadr1DzRR1sQ+vk9u5JxkNZZWlvL8KzNE3tPX5iEB+UyoSCzUHAMY3SfOD3Tpm1Ipjt32cPEzlDXstk2hWfOc2a+++qr2Ka9//uPzYtFWIUtzc13NShuxqhmZgBHttxxoVUMQRHpPD9rNG7G0vBgD/b2SG70xvxBT8iH6+3w9ZVjR/jL/CUMKXmZ8cCAmZfC+qIY0SEHlIVnQk6Pbl8yNwBoS8bwYxgvYI8S9B0c8/xqmaz9nMsIzM7oW88heN/uQJtpai4OTYzE+3BtH9++OuzeuywdpdXUj+gaHY2EFxPxWjI2PKkccn9wb733wcSysbER370Ace+65uHdvKlaWlmIAObahHTGT8oeY0pcuM7klbCI+D+viwYPp2L1njwZfIJxHdu7Ufvn4/Gfx6iunY2YWvfjr8aN3fiiZJdby7//4x/GTf/9X8pY6fvyF+Mm/+8s4KmmX3TLHvnTlevzhH/xYe+HiV19nfOlRLaKzv7/PuQ/SNH3O54lJxaZjX83OFNvBTKO1jVV54HEbQVY/99wx/fyFLy56XacptfKjre04e+ZUIGfLuSIjecBSNVRrdMaLJ47HJ59+ruYIr0lcKG34U6dOxc2bN/S8+R51ByAw4iCm6jRCeP408nSeegKcuUlD+4j35DrFFG1rZPN3xxY3BKupbBaU5aNALHsvOq6xXogz5Nx37tzRmpRx8NKS9iMSuIePHpVMHWuXuEbPiZgqxrdYGksGnS0sKc5y9t2+fSfGJsbiwTSSbxuSBcbzrqenT+tZKFadEwyZGTbap2k7ZeX4LDWMEJMzpVN7iCtZ+5An9icojjNaDbAEIRRLvSYQfH5yNwBU5EEyJhcYwGdOsU25fnJU3cPs5tOUraF1K2d0HmG/Be9nnWG5r2twJeZInz0+iJ+7AdDNzspjqFioAPswp+dzSbkAJuYyg2/n/2omJntUTP5CN1O7JRPTgwryZMsVcS2W/Ckjdc5TD0vc3E0pSGqGlLHZ3KQW5HOTx/BzyWRpL06aNUJL4pZ7wHVrEA6LTua7vYrzvFh5VhCXqOMYLomtQJxPRr19RIzc1zPJwYoHcV6vf/yHfxC3rl+Tz4SMtNdW4/q1a3H08EFLzN24rn34g+//npHOFETbHfHB++8rRzz3xrn47PMLAlYePHgodu2ejIsXv46x8V3y3iQ/2W50SaaT/gRIf56tgKEMJ3p6BORZX11zL0Dyk8gQ3m16SMr7UPvLHjP1jHmO3FvVHimbw5qlDoGZVQCZqr8MZujOXkN5ZZltx30z4AtWDL5Wzk2JJz7H8dgsj0LXwdWMfXJQUfkg19IE9uXzlh8c3pDZW/JrZO+pERrmyvMEabkcpAI25B4Rd8VyYOhHjdDBzwNosF8qfRzuJ/sXGbtV9ocUEZxD8AVYRb+Y4EHXZ66l2r8MnjNr+UkmRLEQCnhVv9eq9ar+dywsQEjVKn7v38ymePJnnsyrn5Zn1xp/MlvRz2Y9ZRlrS8JWT6j1861rqufbXgNVDe+601K8Zt+7tq/+E+tFTIiUFKvX8mDEn5380PUI8ohm+3K/zUxuecGWVw8xtPJqADyW6rPkNXm/aoKuLq178j1i4eragurgycm9imEoGmxsbotVxj6TlHGjIcBS9cTEyE6AjeTrtiIWFpc0LOVnuY6lxQXFxck9kzEwPCSJ1s0NzsCu9F4y48dswLm4eeOG+oWYdQ/hzSiW9X3VCu4ZUIduxb59+7Xv9+zZq5yeeE0ewHpG2p465Bmj4u+Tiz/7nX/SdwBGBQeYtR2trSxd3jzsNCFNQ2aCGRuXw5RJdiVP1oG3DEoVhqYwWeagEpIKvLPzczpUmNLT1JO2fadNrzGUW1yYFx1c3g6j6MltS9JHBdTwkP0M0I+TDqoHKkoUE03gaarRQgQukgO05PkdEmO+SBoIZgQCgiaDGgYlIFkJziRABEZJRimIk2xvyegbHdrZuRklMtCuSKx4bZoRaE6j+SkzrDT/VaLR2yuzODMlNjUl5Xdq8u4g3EgTtIYOVw8/ko6mgGTpCA4BF9BmrtSXEwVrREsmxF23praqdE71rRZSqlD3arzlgVKoGBkLJVyg6Ma8l4ojH+P6jFW4OFlCGgB0Q08szs/rngbatSqCVoVI4YCChi4kNgka8mN9vUrQlCAi1bIVMn9bWVx2w54ElkR+eytmCs3JYScEElN8o5Rn5+aFqpVcVxplckQKQZHa17yHTY5tolpIDp6Pnhn3KGWzmKbTcKGY8iHTY8PutiJS67rJqKgku8UiaqEGnOg4KSnTrFZC5CGG955+LjU9pQ/aZFr4abcPLJqDihyC8FyUkGQy3h6AnpRJauVCrQTEGrG+p4WoqaSt4CPVpyCfEz4gkwsbiduQU5JY2dAVDT8N2p8aEHPuUoUue0FrMxG8YtqkdEw1F5vJXxPSEvI2YFDB+1HsUowRY2SwnMOQkmSSTNP6msyMlRQzzKBRx2CqaZbYEd14GKQBNTFgbcUyYawHkgTpZarx3uXByMqaC43+/pRmYwjoe6qkO+OpEClKqoVptVQb2qoMCKVP7CEajRCjG82wkpxNd1fMwppIBBMXSIJD01aSNOz1lHRwAupGg4aDq0Yx8q5GX3Y1Y7SQtWpoV2FpWQS0ctn3xFVTvL1GlVimXErrefhvargmClvSAtJNXtNnYj/KMK8F3UnDaptH81mRA+G+0nRo91CqgZj1M1Jei8JY7Aj7P/AzxHBJYaRuMmcXzWueGUummqAqwDRAKb8CDBVH9Lxoanm/+TVdgDhJrnhcz9VJNgWWJQtBgxajQuyLMoTXGrCcjvdRShKEZYRgv5CA6jmkIaBf22sgATn6g+dhZpwjNQ05M9aQvcthRKLMau2BaFbzKNGYHrqk705n+gxUDCn2TBsj8qn7t+2b36bA+vsMK1jrgwP9kllin7KmaQxwr6FTC0SQBpycNcQx9ouGy8l64C4J8ZWxVgURKNQ0ceV85t7cm7qrs5qGNPGewcTy6nrAnuxodEnzmN+VBBc+CSl/6bhpyYhiIHhQYWM8GA3VhCD34HnxnB88uK+znPVVzXv+zh5gL97Hb0lMoG6tcxqqFFUgrWmgk8tQrPT32wyz/AO4T6C4fE53xuzcnJtc6+tik7E+YVSYaePhPfermoj83rVr1/RzktkQq2xB1yRkfV5vmaJqz815qIHsldbi0qLRj8SPlHnZ3AIsYMktcrL+PpqgINdsZunmlxl49RxrkMu1VzyooX4XyHQ1IpwjIe8A+ozPpGtYWFT859wWEAF5sIzHnC0yXE80ZwEK2hsIyAbR2CQPGB8fVe46NDwQF6cfxWLK2fxd++Lp//4Nw4r/xCEF79Xf0x0HBwZiZQl5g4VsMneqIVZAngJwmNVlcAv3QwO9Jec58pTLQYbP45R1yQ9UCN5qdhh2vR49jY44ODkSE8P9sX9iZ/R2MfhjiNUZE5N74/bUdPz/7L3Zj6VZluV1bLw2z2ZuPs9TRHh4eGRU5JxZWbSqEYiWeOIB8Q+0BKiQEGrxgIQQQvBQT0iINx4QiOatJZquronKqXKKjIzR59Hc3WYzt3m4ZoZ+a+393ese7lkZmRSdJbmlUh5ubnbvd7/vnH32XnuttXfqB+X0mVNSBfX2D5Z7U9Pl8exC2T9otfIwABTWQmetu+yg8kYBs0M+zPnZUmrMWNhHEdSpJrwBEuqLjtI/OFg+u36zvPXmG+XOnVtaszQiPvr4s3Li2GHNIbt77245zsyLzs7y6OFDKRwuX75QfvXhLxWLL19+o/zZn/+FLPlYq7Cka1gWYefA/Dgan0l84Xzd2pSagWYA69EEof0yOTGpa2N4vJo7MH0PrN7j/mtA+O5eeXD/vvaaSDaRR0ESuHjhgvY79QW3BQKH2aSA612qL/C75lqoyQT4DwwIpBsaGi4ffvihcvCBgUG9DnECoJ9cmNdnT+iMCra0BtxqCKlZyuSZNOqID8QuFN45R8kx377psmUVQGTGfwJPZqq7huTz80UDQOS1yFkELoWtBnUm5LG1tZUYoBxDVYnzUWMA3EJsQrkl8KuNQewbUl8TM4n/bW2dAl4hkHFtqWJI6zj59BPLY/YTgLfqBzWN/dlzn6jmDVWaVdzON1K1nLbBylGx4AlFBLFN87EiP9Y9UQJgBa389YP4oLy/lQaycy2+eN9siKTiqSKWBcFQ+YnstkxycY2+pRqOtct+UT5PrtjXq+d59/597TOaa1L0YJei4e62Phapi0ZU5Hyqi8JKWJ+l8sxvKC3URI6mjvRYkeNZncN5ayszrj9tn3gWUj5ozlAjt8zcS+S7Jmst5erkURpib/cG9hn1IGxp1rwUxNT28qavK+6x/lUDYXGGwiBswWBFewAzGAg5XjLwd8r3vvvtsrwwpzOcZiJEStYkQCdqzcdTU6WruyYb9YexTAAAIABJREFUqCePp8rpM6dLf19v+eSTT9Vo+8Y3v1F+8csPVO+fPX++tLV2lNt375XRkTE1KYgVBy1tZTNmJIowoRkcbhpB1pP9ms7GPcUEeeiTI2oY+IY+Y4K+tmrLJqOVQqiJsCvL5n7ef7shuPjK+oL8ykN63Tgjn3U95PxXVt946JOPSKVA7DDh0ed2WJQGmdL1mtxpKsW/1wSse+8x/S3Z9aFsyiYH60yKferK0sA1dne9TpjhoRJcKu1WPZPEWbJxlHsm7VPJE8GUaGRyYdwbg/hWgbkEb5ABs1mR8+GsTg7rt6ZGRZKvct2+eOZnIyKVaI2mbtrbJR7wfJPi78qX899f9XN/1+9HKKrUEY7ZnjeS8ooXsQIRRwKTsirNzdfEgfSaNBZUszonZi3yOnmfGusxZuIKf3Eeyvqq1bAld+7o3BJczYoGnkUOkudavHcbc35yBiK1DeuC36ExcOTokfJseVk57sWLZ0pnd0fZXN8sDx480tnIU19dNYkaggTnHAs0idtcu1R6spuL8zGwlrxvxFQ1ZVBvdbQrz2eP8H/2K9dhtWoR2WhmZlq2TzRqUV0fmpzUZ2fdclbTxADTIA/9CNvM7i4ps2imgDWi4GC/QHh63aj47TLx17/1e3wHRhjQW0oF1CnwhCdp1f2tkquGt2QWcSnL5SAhGUCWxUFLgsVhAQNZoI6aCbbLIcklSSaZJqliw2PzA0Aohmlbm8G0aHQQ3CgOGAA2OjZaOmtdYhYB9stPL4oUCgcCGgkaRUtK2QlwvBizH0jESOiXl5Z1HSgmSLwJYpIjt7bYl1n+1EPl1u3wm20BbNzTgFvY1gzKFXOjFKkEnj6ZVsFA4ePBesjm/UXSnnKxyiaptUVgPc0ADzq2bUMW0wYZg/FbzPb00Eh7N5rJvaNrz8F2BH2xYTSfo2Fxwn3RwRmAYoI02cVuBh2VyPunA8zxp1CiEclFg53rw0neqsEMFuhDkdxVK9uyxuhQ0kaBSjMIAIG1w+dp1WBRvCI31HUGRFESDJOnXi+jQ8NKPAUOAkJgO7a7K4CGL1lPhX2MJXUMOF92EodtgfwOYyBhC53uTq1zhg0rUWiahcA9OXHiRDS3DCaJcbq3r6Seooc1TVJsQMUAo5IoMcyCbSFVgWXjLhyw6iCh8zwWNyhi3oNeJWSWTewJs0Sen1VRSQqakifnly4g45WiKHDClSBOFmb+6YZtjxhzzyWPKd+1Yqa6jlcwO/S2Uq/HSifpD0aELijmdoipx1A3WKtN198cFpW4anC6lSeNostSUM0fCPD8ucuJz5DJFGuHooq4Q0Ep6WY0G0kOskmhZgGScZgW0QiSioEkfBOLOCc88j1HyRRsbQPv9vFOaauKVQEHWCdRGNpfmnvBn6w7MzvcQHOik2C/m4pmpFIYWMHBfdIeZlg9AGYMhRT4iSpEiZDtkPisNHrV3JFipCOGy1mKm9YvJDdq5OkaWmX/QqJDIYQ1ntZmWP6JKQeTVnZuB2K0wGQSUBUDipV05zpryqur9RDPEfUJccDzO/CV9TwNAFcx3GL9VjMGYmA1VmwoJhgunoWCioNE6jVjwetZDZ8XZlQAMuFVnU0nzasJ6xnuL/tSxX40J1muyWxyXG0vSwwnq1g+qSxgf5iprfcOv99UVnCfAYjmpKgwCK7t0GRrIBVX5UPq/a733t8TwEuMSeZQMoYcd11kcws0d6gaXuxrGxsZkcqQ81LnSVovpBe5JPieleEiJM+FBBTMMDWD7NUDr5v37ov/3dyo+E0KpF/3Ws3/xrpjL7AWuX/aQzrz8aPdUJ6Bh6xyk/Z2sXBpxLGnKUwgPliRAwBa9H2ePwSIXJ/saZ7fjOaLeBOwLgFtmebR29cvUKGlrV1ApJh+WJLgvR/DMMk/sgkEq5O9T56hvAfVTbAFec2xMSsjONNy7pQtmNxkGRxE2eNZKQbJugT0AsJz/lNE8efQ0KCtIDsYPmvwjPkUFHKpYOK95dMe4AKNTjUMZfPVYLGmmiKZxQwB5YvrIUfiT1hexBnWCo0OFhL7jS8AFNYAVjHcTwAeYkvacFDEifUd9h4AIeQ2ADhpc2KFF5ZZq3o+Bkptc8Z+4LNUwAy2VbCH9fld2GYzg9fLhjIFMwAFz57rV3xumtfgpnEMWFeR7TOcLxQVlJWoKnmPgcH+MjY2Un7ywCz13+3rhWbF/wdNCq6H2H1xaEgNChQ5+VxybQpEVtxxbkIsFkgcLP0cvOqZal4jrE2RZAAiBcSaTGAVRVhAII3BLrWjtVw6zYyKztKyu1FOHTuqBuDK6kY5fPR4+eTGQwHLV6+9WTY21kprR63ML62VueVVNZchCOClDyucZzs2PlmWVuwVT8MScH5+blaMRAhOxHOaYsQuhmbj4X7+woVy5+79MjQ8IJXb48ePy+TkpGLt40dTqicAcf/iz/+6XHvnip73L375Ufna++/KjuHW7Tvl29/+Vnk6PVOeTk+Xt9++Um7fYeD2ujzffdZiOYftYl85wRyM6zcqv3ipoGms1Pc0hJ11e+feXZFwzMal/jJDGRCUfcJ+s+Wpm94JxDIjgi+UyUlskvI9WJ80o6ihuAecCyJs7TqvOHr0SHn85EmZn5uvmviwzNlPAK6plJFCUzHPlmxmC/tM0GyBUCTk2WAlvWdkNFjEJg8532zYtglsxqZPRBgTO8iXOCs5a8lBPJTdBA3ee3xsTJaszC30vue1qSFtN0e9Sezl2liPqazb3oOUUJM9IPdctjk0ibfNhs25OiIFiYBgtq4Y7Kw7yChY6kg1h3rFCsbM+bg3sqepddmqp7LtdPOiQSqL+R9hr+x7ZDKGm71mCGc9zTXy76rjAvC1zYkHtIr8E+p1k2P8XgbyDbbnF/kVA81RGbBvOSPSHhj1yfWbN8pGxHF+x04IVrQQP722co6Br5N8TDlbANvC/LOxpXVeV53HutesqBiam/kbMQIgTnX/DjUtQ9lbpZIFZAOIzBysWdGptVTNCPBZpSZOkF4SpN6B9Aaruckui2vNxp/sfNkfAjTN6LaCz7OVzH0xccOh/6B851vfKLNPn8gS8tLly4ph1PisS2Ks5r709paLFy+WTz/5pIyMDBUUTDu7W5o/ATDKvAri6aVLb4h9/WjqSRkbn5ClJHZb25BSIGBubYt8Qk3C9RCfVC+GQtruAR0iA3B+82+slZyzkYQV8rqsozw4nnrB68rzSFpUb6th3+5noHxWZylWUpv6nhsVPE9cBpzz8nedvQHOkn9kM+9FMlpaO+n5qySMOQpRL0hFnbMeQ3WVsYM9lcQ3K7LJ62yXxvoifZUqimZLKGG1ZlSLmTSm9dWGVbXnc+TAe/YZhEfVD6R5Uga5lnU990U1Q3M+XNlZ5Y3WGBbPYvG3QkWdyqGo1dNRQT+WCpKwJU7Saq715pzid2lAvPh6zaqN5/LrmE2V+JJnTrhG4suX27DC8r02GVH1esw84Vo5v9xwME7iGGxrONdL5O2uTzVbJOqUnEVmhTnnuNclv4+aem5+3r8D8XRjo7JcznvuZrD3RMagnD0pF4ODA9lEclZit9pZI2dYKR3tNV1fd3evcnwwwo31TT1T9o7INvoc7VJzcz0mt7khbfIuBLZONbyxaEsSMEtJTX818DvK8NCIznkpkbu6y6NHD2UZV1la0YgMK2qISsxi4l6TR/MnDY249cI6IXObOGvC3etGxe+Wjb/+7d/DO3AItkwwK5Mpr+K7GsRrUhNJRw4DNfODxMYsZMG0+KkynDqGknEQ0CAgIMFYzgGLgGoqIiWn6tMQU4HwDLXq7BRTEMYCMmWGMr9x+Q2BDQyoI4E+feaMDsqHDx8qqcFCSsPBovkhAAIgo80dVD4bP0MQQkXBh6G7CZOBwEBHn+SJz0sBA6iZxTxNh0dTj2KYGAko3qo9lil31xToXMQel6ctrCXJqvGN3tmpus1u3LSVw4cP6zqQHHLw0ujIBCFZxEraInlLFlMykDm0CVKAMZwZav60twu44QCB/Z+JqFj4wQQScItftWZUeOiOgIzqfdJ6x7C1WEDRcEiGfw6+5DBKRmagGxUTMZPdvO/4RZIgDA14aCT3j2KOxH9hccEMiPbOsrS8UvqGBpSwsT6QXuIfPTY86iKIQllsCk3ArMBDsZyCwQXYSvCnmUWzoqe3V5Jg2YPARqp1KlHkd1CrOCn14crz5/vMEOH3WT+SauNb3tOjwpifBWgSUykGh7HmnVyYXZEfsrlRYRaQiyErAvyzmXhUoF4kLealmcngvlA0igKQ9ZsY+cxGhZIBsbr8/JK5EJytKuq8mOzke2cSmYPxMnGVn3CTv2gqdKr31hx52/g0QNO8vsyUzRhj/gj2IdV9qq4qPl9I11X4xDA5zcgJto3WcgCL6SHefP2NRoWLWT8X268ky9ZDtwxmEXuIH+0ABiT/yJ0pzhgsrcQfS5etwiB3sSnqdQ2u5jWZDyBLFyVM7QLSsBdosHr8Plx7svbM6rIMX0zJSP60h0PJliwS4iVgo/cpTeSaQH0xyClqY/i3mwmxBgVMGWRS8crPR7OMtS9gI2ZKSFoK4KEZENhOrKuBgcw2FTTeGwznwyIFy6RIKIN1rXkRwfaH1Zr336lsfIXvP3GW+0ThK//6pjkuFKWyvAufUll9yb7FQ+/4b+TxaoBFs9QsxvCVDTWP2D0UMtFU5/qJ+0vE6GpIG2vCjd5cO4pnHR3y019aXAomj88O1gtzPDKx5j0ru6iIkyp4m+yZ2Hvcb84+GhVmYppLZgDCsmUzqcymFdMxbGe459iNrMHoCfWGlEAxiLxqPDBwDW9xGlRRuLE/PaNiOxoVDXWWgJ+w5aBgzUZE3jfw2rwmN02+6JnbDBRU2/cl//Fio+Jlv/ebvlbj5R3zenu7bQ14UMT6JtmHLc9nlz1QS6sSdxVbMcuF2Uisa+IZuUIqQOkt2/rAw+s5M4kdNKaxlsyhwfwejGOInqzj3r4B/R07u1o033jemksyMxOWB7aBBMzg9TlDBAoI2AREs187ZAizQa24yuHVJgDs6d9zbpABsD2xkDXHBmZyNLdsqQKrvKPsHXgQH01bgDQVkHrmVjJxlMjmAyuUtO2IuStcA2uSHIm1y7qkSU+MIGYCyGA9k7ZW6TXPmcH5CDDKvs0vPquH4vrs3dre1E7Y2fWebz5/KRL5ea8NW7BwZvhn2jwoULHDjU6RYDhbovlLzNRr7+yIPHL+/Hn9LnH09q2bWieAign45eworpXfyXkNCR6mFSrPjEYFgPT0zGwZHR7UZ+ystZeP5haqs/zX7Ykv/Nsf/+flZ3/6j0vXX/4P5d/7j/9VuV8uln/2v/535T87f7/8t//Bn2hw9ql/+qflX/+nF8u9/+lPyh//6Y0v9fKKwy0t5erkRFmYX/L6lc3qriz2TCyyOs/kCxfi7C3bcnr2QYLVaS/TDKYkoJh5hYChAOB3d7dKd3tLGR/oLkfGB0t/Z6sUFZOHDpUbN2+Xrt6B8uDRTJmeWymHJ0fK4GBf6ezuLTPzy2V2aaVs7+6pgfBs+VlZWsBys7McOXa83H8wpX1HAw+AHdsVYv7E+JgsXQ3Ytgvog5AC6ICV3sOHD/TMyNU/+eSz8sYbl0We+eijT8sf/dEflo8++kjNhvff+0r5/g9+IMD/m9/4avmzP//rcuL4YdUdN27elBXtrVt3ytzcgs5oAHK+uKcobWA53r9/zw2CGHRFbsHagkHNfiQ/pY4QSamjTTmqrQwBL6wA07m4ua38kzOTXNY2lsz9MxmMtU7j343P7jI2PlqmHk153lIMomWNQ6p66623yvXr11VjAYZyPYAxNC94HccPzwqQ93fkoMkQ1YdUIwvA0ENT01rSdYZn77CeuHaaYsQa15Jeum6utCiXVyzY2raPt5TxtsSAHcpr8N8GQEsZGR4q46MjqpdoZrB2e3pQDHj9SuXZZrYsANShw4fKxg5NJDdRsIMCYLf1mUHEZO3T4NSML3KmPednKDkAqYj/We9wv9knfC6IJ9QkSZoQEIeCRZ/VLH8G/UqRDqmDgyNnOyiH8KBqx3iT6/IMkhI5QDoTFJwrcE+l9Eiyi3IaNwZ9ZnSoDsyGhnJTMeit9rXlk61YOKcePngo0hcM9cHBIQ8gV55lFaxjn2vIZOgLnNuh+dFRzYbkuj2HjpkCDHVtkf0I61X5bACbjRzIGSKfC+KSmhqhZlt+tiTCQZ59mSMkQMzvpIoklSbpae8mfqfmztC8Z43kz6RrQmdXlwBsrG1gMe9jQxV5kdnOkUPK6tWzrCAlff1r75fFubmytLiguEHdQOMMGxbm44BF0KTHLeDmjZvKo7/9nW+XW7dvlNOnTunM/OEPfqC6//Ibb6nJyYybvv5BzaiYevqkrK5vKl/hOqgJ2IPUGFjB7Gjod1vp67H9DPkL6wASDV8muOx7HwDoBzGR/Wq1rK2FyAGSXKPZjBDD2LPx3zlzwOvNSh6eR85tZN3ToKEO4/VYn6m4YZ3pe6FOSvVw1h16ltVaCLKRZq1h0dlQ2Mi2CgVfPGtTeIrmf9A8EVgsS+pQghC8VCs3cCyuu1Jgt5bS3+e5MryQCELUVVgFbqC0N3WO+G0SqJsUJhraHSC/sllvAlraMjd+z3lvY79YXcAzfd4qT7VVYDHCN2KGZa7vFw/65gbJr0sCXsy7MwfI36kwvZcQD40BuAmhuIESEPVMEOJebFLwmq5LcqaMLb+sNLflUuZyfH4rdk1o0T0KfLE57rmBG4O5o76EAEoMhrzF9WBfRw6XzQg/a2K3rzXrM6v5Yt3jQBLnEucOzW/ZXqpGdyM2Da4h9mAxzLo4e/as1oWJdVi1r+n85txRjrhri1DOYKuMrSpC0UceRWzjnCfH5vr6+waCkNRZRkbGVL+BC6CwhHSNNS0xtKV4jiC1qmYU1TqEHfJ8OB8hahNDyKv5nOSlxAk+E3n760bFl06VX//C7/sdYEaFDhj5UXpj50BtgglgHQHbgIsLdb4oWtXJRxa4vSN1AMkCxQDDQDNJECDdSlAzWCuZ/c62EkUFa5JcDufdunw0J8Ynyvb2poa+AficPXNWh/L9Bw8UWE6dOa2EGoYim5uAQWKvjnvYqgDYkdSSGBA4T546ZTBu2UEOgAO5cwYrEjc+C8EgrQrwOtTZVsn6DDjTKJg8fKhsbqxLNYEtkAAyMX8XBXaj9pifn9dwPakZZKfQq2SRZFCWOrDRYmi2gnZI1/RvwWiV5DM8SDlA8aajcCeY8XMA7nx+FCkkCpbcmu3tgG/7H35W53lKKmWp4zMjAcIEBzKJTEmvkwCzTKrXbLKecrecDjmJKn7ctsMhacZbmNfv7e6S/z8MrhMnjtuGC/BSDJyD0k5RArASUkESyz4K5s0G4wbwrdbbLbCYQksAG8qZ8LSmSOUaaEbBfOVQIaHh88PI82HmggBmjBoye8jYe+WjzfwRwBRdE53yULeoobSyUvmKmz2YTYFQLYQti0CvmM2hg1w/F7KCpkCQeYI8xLn+kDrqtYMRryQyEgHbLTS845XMBaDPZ1IxExJ0N0Jy+JwTgmZQMBshyZLg2WWzLGy5o9gPkD1SCzP+ncDnAGL9N9cr33sPNnPx6oRDDPZI/rFY4gGryVlJjZ0kZsFHcqD1GDZIVvyY8ZIepWlLZPWFGR22K/D94YRnTViCb2ZxNicYPtXTDSPZ90cJI0UhSgsKM4DfYMBn40INKgbyMQtHn8mNCn6eL7GNgv2cagMA0GTV2QO3oYIi4WG/phxdhQY+76EA4b3aSfYAGxnqTuISBQX3gDUqhVb4sOKnyQBksZ8AwePe2nogBk1Hk4Hin/jsoXke0kXs5E/NQ4i1X+39L2TMLz/Nkh2Ua8vFtdek7IfkZ+wvkjwntJ1iUvEMie8UX1yu17NjLcCOB9oDRDeKDzFtYOhg1RDdP+IvhThqllQEEOvVeAzpOmdXCylpyNNzDcgGKYBsfL15nqwhfm/5maXGfs1mr9ocbm3mj88K92skyx0ZDoAkiz5Ysx6W2EjG3eRk/wOKAG5xzcQys2d8z9QwisG/YmrG4D81b8RIM0DLvhPwvburz222PMl4alx8/VbAOZ7nhSNRzuLT7+X401wkNRdCL66EPBvy+/mzL/5+8/dflRsl8Pn8+xntAvhnP2P3Ymag1z3nN4PTufZh5ljEEHs/MzdU1bAHsI3mtIcrmjnJHZJ8WoM2W8XuZNFVFoL7DDjdVeOyo6NL+jn2Jx4B7B388gEWIECYpenYNDI6ogbi9My0h8yqmWCGFM+G/AHwC5an8wIroqyM3K+GdJs1W8rOtplbmqWE6i+UJBRwkCdgX4E3AqDAasOqkuIKAEpFHfG1hSLdVlRmUPv7Aoywi+nv15+ALwlM8/5cF8Npyb34wjaGM5/v07xIBRB/Hx7GvmwzXtNsSBYpuZ9txwDBvb7Yy73dPQLeiKc0Ng2eOHehOKtirPIYr1WdsdGo5RznNfPs4f68cfmy7i2vh2UT98pKQa9/9jTxFJVOc4MoZ4Alo5D7cvHiBbG4Z2dmxUym+dXT21V+NvXkyzcqTv8n5Wd/9R+WdzTXfKdc/z//m2hWNHbEqX/6P5bv/7P3yqTS7dXyV//VPyp//D+/ase8/Pus/WuHJwWqSzVTiuYkaI5Craa8xg2nsD0knspqyGcSeZhtJZuGnMbZnnlxEjfc5ASsH42ca6e01LfKYHd7OTI+VM4fP1IW52bKxMR4mZp6UvqHRstH1x+WtdWtcvjISKl1MVOov9x9+KTMLa5oFowUrqtrZU3rba+88daVcufuAzdUenvK6Miw2IioK1A5MxCaGQuok2go8JmpG8YmJjSv4datW+Xq1bfLk6cz2m9/8O675YMPfilg+r2vvFf+r3/5f5c3Ll1Uo/gHP/rbcvHCWd2n+/fvayD3ufPn1Kh68PCRLJZ0JrW5NmIfmf3Yo/VG80HgCIpfKTVh6Rtw9FDpzdJR61DTgi/2CvuJZhr2VTw7D9JOr/BSLpw/Jx9qCD3ey47f5BS1WrcUGTQjkp2frH7OvcuXLpWHjx4KaCRW8RrEHq6dmiSZ5ZpPp7zDDcBsrLLPZdEKIz6Ueg0wyvvJ9kRuZCQhx015nzWpJq/H0HsDpczds6UqcYCYvrgwr0aFlF/bANAorSASjYvERl1I/cX7U5/QoBCAjX1PWCN29wLqY51kdSl2Wfr3aMDRzIKnrji8D8hFIwOlv1n2qcISNyptYaK+5JnkdWn+WYutIPUsQoms/XDgXFRKJtnc2mYwGxCaN1RDScYacU4KwMX70ywnRtOc0BpobVFspGnF+iBPpEmbZ7QGukY9rbgZ4DWNbK6DZ406jeYUa4w5bKiENU8FIt/enpRJqF9VR+7uep4Rlsz9/Z7pxhwNT1uvVFg69yE2UI9ubJQ+uRdEU4p/C1tmGnr8ruYk9PTpmVhBjMIFlj4WJs9U36a9Dq/TnC806k/XF5rhFvluzqdqb2kL27p1E4kgoXV2KJ/a2tmJBrzXKtiGCRmcybb7MvnI9k/8N2TE7/3hd8r044eqE2Fjc400Q8ALuNdYtU0ePqza//PPPtV+/IOvfqX85CfEkAtqzrK27ty+Ww4fOVJWV9bK1OOnZWBwWPnlo8ePyy4OCaiCsLlhPYY9I8oXAbxiqXcKxAdHYP+urK6VWneXZ2ulKhkiE3lwPKfK2z8Aej4razDnVWWMqKySwurJ+Z9Vc6p7UvmchLIA5JW/x/xBncmRUmZuLSvZyP81wyfnVuQck0hyiZWuFa1UkqsCtVk0tViD1PTGSlwP5vrwTEn/Xb8b6nb2wzbDtjs9Iw/MSqp+6u5aTXhN2rGxNtifPvtCddxgXEWabCttKUkCYzHo3kj+MybnvtQ1BTnR/+08tnJBiHub9ysbSc0neu6BrNnzZzM3a86T8/Wbc+j8d9fwDZJW3r+sX7JR0ayasErcV9Pc36gUIy9JPVxfuPZ+2TXmrzRe11iVrzMa//W61btaWwf6b/J+7g81Oxgee5p1jsVyNk1Yg5k7m5jlc4dXHugf0FrFnp35ueyNnTrz4uxcQv1FvANf0swJzvDODg20J1ek8QDmxHqzGtggGtcO6YfYzeft64NAta0cheYf7gfk4LTq5mbmNNeK2oPfHRoeFhGI5if2r8Y5mL/iRj3nCmRfYkqe14NDw8IyiflgjcQqiHa8hhqD7ZPvxyP7cgnj659+fQd+X+/AxEEMlwq/RzaKbEaiEyzf9JSFd3QosSEJElukBV/JTTFHCTIECQoGCl02H69BIgb45EQu5IYxEJrXIgqK4bK7qwbH5MQhzX9IhiHsXxImEhz+7BvoNzC/V1exkDYksg3RtdY160CyXNg6+wflypUrAuPkvxuMXYAc7CAM5jN4rqZEIyXPunaG7TKzghkZaxs6oPBq57PzJ79Hl39sbKw8fPBIjJ1Tp06KjU/QAMTQALX2NgUx7o+ZGi5MuD6AKQG84RHtIqdmGS8MOIHqZksTmPk7910glPwp180E1+AhB1wf1OmfGkPLQsKdnfFk3QvQDT/5Rte84fmYLH2ByYFkN3fD0wsbwIfkmgSAhFUXIWk0zCdbU2jINozV3mSzY0WBHVBr6eiqlTV5We/rfgACDfcPWL4qIHe39A8PlrmFBX1mda81vBFGlsEdEstZmDL7BiB0P5S02VInkwiBVbJkarDnKXpZE6xdyfIY1L6x4WHe6+vhtWjJehbuzU0Aut8qygIUTpWDDvjI3jJhyMPfoFQMKqtOFr9OqimaCB3VZ3AS4oQjmRkqXENRkddlL2lnGinDzPdGUqnGoayEUCtg52ArG+3lAPJzsGmyu7N5UFlZRTHGa0iJEMPp0o4A2IPfZX+SrCeIraQt2fcCXJ3wiXEXDTU1A0JNK+ZGDGfWR4qf0eeu1ibJtfdCrlEl/uFnz3XAcOA+WWIPkwaYcackAAAgAElEQVRQsTEMksKQ2MEazEHgJCGoHJTo6b45aTMr2jMCnCQHIwfgLxKmLHwE7EQcbTSSDFqzdlVsBEsFMLTOsGSK3WApal6NhlUyoNwxVXM3YqaE1kkWbTFbJJl4nqXTXSkyrJJp1wBeYglzHHTtshGw2uqlXy+RQ/s5JlvKRasTXq9NAxT+nNgAKJblELVo1Gn+hp6TLScAHrh29iL7PguxvG+O9XseoBtMVP2O3sNMRX6W8wVmX85q4BpIfNPrWfNFIk4IoKNpHjE0BzEuLi95YHd8hmRH8TkaIEFTM7LFwzMBnQBv3ajy0GviPzZi2Vzz4wr7FTXaYOgUWZRgC6SZTzTOomFh32cXjnxyNYICVKwaFYNDUi9ZIdNm9U1IrWWJos/XaLR6mC6FudmwGngeDDzvLX+2tJf4TfOYFxsXuR9/10YFigqeMTJwgAPNz6LxVYM9S/OSZpDnvLih64LCQJabZy5mGOIIyAjYEwWQQDOGkDrmsx8EdAPY0nxsN8iIBzb+xjpTYAeHpZwBSM9/kUozYh97z9ZP27ouzmuBQfW6codULSRYoGZCFG6AinwOSBf2923VzAmuAYCHgXtikW5wdvXp/8RxgFmBOWI679ktLBQbAFMzWOasroutxZrM/ENgWU9P1fTyPTLQw7ogbwEwYOHRUJPdJOCIGhkGfRiYquGw0bDkHnZ0OtfjvrPvsGPQ2R6qxp4uGGh9lWKR79Mseu+9r5Q7d+7qfQGWtBajOa/GOXt6r677DTudLxFomtR3rGueDQ0PBo4Ts/n3nH0hVnawetmSudczjhAjzp87V7Z3tpTrArZz37AB/Wh61j7XX+bru/9l+fh/+Sflko+gLzQrnm9S8O+r5a/++39U/vhPv8yb2PrpjbHR8mx5TcQc59AmDGleTyhqNfxcFiA+YwR0sk7DzkZBKUAHrsDFtDGpBJfUcJWFSnjPw5BvOSgXTx+W7dOR8ZHS09leVpafle6+fsYEl+m5pTJ66IhIDsvLC6W7b6A8fDpXnq1tlbaOToGKAhPLgQp/gaAC4IIwUbeiZmtzw+q0zppiLmdJX7/tXktrmxojFy+cKzdv3ioDA6gqjpVPP7teTp04puGrn3/+efnKu++qMQAZCEUWYOBnn31erlx5S/Hgr/76b8rVq++YrLSyIoKLAG3uU8yS2toB9DDAL1AlBlPTNORn+rp7tbYgb0F80PrC/lS+/wflwoULApGnph5XgBb5p9fpnkDSZ8tLWsdJSDLI36H1PD4+IQUh54gZpMz5qCmHZf0zmJz7A+jD3xkSPnlovGqK0LDRUHkN795XHu+5VhlHbfOWA+lp9mCnx30g7rF++Dtg+ANmfURTvAGecb61ld1oKGrPyr4HK7ZtXQcqdl5PFl78T4N7aSTURPyigcI9XBHQ5NgG4cHzVQ5Ug5DXwJEFzFLNEoqp+fkFgUzkfiiM2lHPpoKhPYfa+hzGYoZ5Z9lgYW2ntZnylSAPeAaDiQxWy2I7VNN9z/ghRvDEuNxk+EzUcIBmzWcqtl4QDNLdwNZqtrpN9ZMA9c5OqTwX5hcCVKUZ5lz+IFRxkDu4BteKHnBvdYdrdOy/eG/yIzzY+SK+mwziBqUbj56bxvOkEZBWLQ1lppv6jXjSqc/NaytGy9KM9ULz2fmtYks7z9CxwvWIgc2Z2Wm9d+ZYUg9HbM1GaDMo69wqt7nVJQcQL/GjF5FvS2sdQiH5mAflQk6jMWsVkghPoVxlLZissxONoxbtgW98/avl0YN7qm8uXbooBjSNijNnz6pGnJud0z2ieX3nzh2pkt59793y05/8uPBcr779tgdR79T13LGGm51dKCOjY2Vh+Vl58vSpmhRcqyyLgzQANuCB0m4aQEiRzTWDtev1Mre4YK/7sCwjV84molRSodLk98VCh8EQM58yR/FMCc+kS/eEbBYQR7OxRlON810E01CL++bHPMxwDZB7QOSN2WStZmYEuc5nLfaZEFfdmPA8nCBTRD3IGcW1cw0QHU3ewWKOOogzql2xTes1CIGyntLeNKEW8gKxkDNfmI1sbLsU30RUhTjHfQ17Hq3xmKbhtdVUgQdJUZ/P8vmorUP3UTUkgiTaNCcyG5eqM2Kehl++MUuE/87GUZ70zes985LmRsWLGYFzrgZRNfePCMjRcM2Gx4tNi6oj0WTv9MXXb/rOK8pENZgi7uZMCu/9SlDx3Ms6d7ADgteO1Z5WEHo2j1wF9vZNAiC31FBt16q8l4iyalz6+atZl+TFcA+R9VJbq/aZm5OdUh9zjtHsaGsBU/Mg+rUNq3fJjdo7yIm71Shgf1F10dhUXaW6whZpzn+9l9Y3UEDWZO2KnR7Ea87nR4+eVAomYvTg0FBlIc91PZ1+UrY2wRTCjrDF1vHZgOH1sIE9euSI5lmxP1bXae4yi81Y4OtGxZfLk1//9D+AOzCiLmIOWXbyoAMrLT5i0CDBHnsD7Jj44vBAXQBLKCX0DKIhGompR3IJ4IZPZqfZKmbotJvF1tOtxoQCqTNjBSTYbST2C4uLCgJHjhzRwbS4/Ey/Pzo2poOcRggJFwGGhCwHD6etFEkq1iYc6vIl1oCcVW1kSb/W1sOmAWkuHUlbEhHoSAJJ2g9NHJL1E6wZCjypA/oYWNmtA5DPT3AZGx0VY4cEmOSHALa2zhBWDvFdD+XpxefUPq6VxQCzHDRs3AkIgBif0ZJ8AybZFQZYhBWoTi3XGUxkFTHhW8/rOGiapdQ8PDsZ+F9YksFITjZwdXiFVVEyx/P7AuDDmsFJvBMsd38tPdawWrEoGATcWXYBRFtbyskTJ3TA8Jynp5G+9kt+S27T2tFRnsxOi/FAwck9GxsajpkH0myWWk+PBoByiNifHBuMdnWfuSeAGQywTQBX7CYBp6UaTs5aEcu4Aq1aVRwlsCa2FJ7hKysqlD1oMFmgDUaCwKQYHCUANfKZZl9rNfvCVqTJEKc6jAWeJUAZzN9UpKgZohkbVrTw97QJyvxJiU3MV7AywQOl+PL+tbTZhA9nFfk8bXPSHomr5z84yfTBnwWeGonBpklmnAqsOPwBiRh8rgZODHxTMgkbq9OKFl1vGz7ry9HQbFaZGNxWkafkJpnqVkq4B2BlipuSlkM2GBiNRNLzJ8JyIRa6Pnc0EPycnBiS7KihE/fHRRUMODfaAKrNRrd9GbJx7j8xhBhGLGSf0qgEgHTz0PcTGygxE2NAc94/qTVChcE6VxEQihfuvTyBSZzVSIhByPFMKcZ1J7QeWuQtrPtczSnwM1d84b7vH2iYeA4JTyWDmiJ4asMEjDkaFFtqBgJMVYypFyLF30HREOz4BfZNYwAigA6fANVKqvJ4r0qaHjZSHnhtH3nFTBgsUmFYHcJ9MTC6V9pi9pEabTEHiGRTwxAPHFuZ16AYypDokBPnvuMTasBxFDUCdAOQo7Blvct2KlhgfMAsog2wGsDJpDz3JfcYwJgzgWSYJSjv0JiJYy9ps+5Rw2h9qPHgOU+w8GlUEM9swZeKDTYDe9OxQHsirkmNwnpdDHz+jUaFmYG+NxSXssyRfVhD1cE1SFmwa6CIhqsLVzd8/Jkazab83qtSm8a+fPlP5F74dT/X/L6NV3EDbGio32eDmIYUJbYiZN2Qi2j2FQBGS3GjuYfGI0Cncw/WRxa6aWfI8+PnUB8AdvM+AH7pbU6MAwRjHQ7gE39QZBnHnxRSnPlZqCgWtKJy9Jwu7jlrAJBEw1E7OlUgsy8FYI2P6z7Llx5ZOXZOMWeBz46ChH0+O8uMJMcPCjpyJ95reWkxGFxmX5FXYUlku8cdKRVy5o6atsGqIwejMS8P+njNbHArJ2lpEQORNcjriG0axS731c3hRkGeKs4GyO91k+ebGdKehUDMTEs89oTuE0WiyARt+myyopECw2xJbNm4L7xeemLnvRCIo2ZEu/YDZzz3l4afLSwONJMsrWl0LkezSjE1z7homFZrnp9DUbezU86dOaM98vTpdDl6ZFLrhBkVHz2dLmvM7vmSX6f+/f+6/Is//cdfaFb8R5//k/IvKiUFL7pTrv/v/0W58ic/+pLvUEp3R0c51d9X1teYUbEisIb4kdZO1aygODO492Yj+jl4plSocOKckkc6Q65D6ZWzk/h75W1NXG85KH219nL2xOEyOdJX2vZ3ysTIcJmdmSs18ueDtnL/0dPS1Tcgi647d2+Vjq6esoUzXjsAAuBDXbadkA8YmEpGCdtxZW1NwCNfPA80mKdPn1T8tKULxX2nWMdvXrlSbt68LZB7bGy43L//QIoJ1hKDs9l/gIcff/J5eeuNi1rvN2/dle3Trdt3lQfy3599fl0x+e13rqqBQZze3KLZ6ZhNQxiyC3now0dTYTOaw67tHX36xCntmTt371bKUc64JDucFMlpTZ8hm6isaxGcWlul2JA6WIpCA0/yB29SS7OWiX/sMfaTc10sV/v12dl3G5tbuh/EM/YyOY9AIZ49ysFo0CZZLHMy22ju6zNSp2GdkuqA3IvEOgCZGzduCqipFBVJTNFzNDicoFJ+BsULWRxZSU6ewhf1FK+7FTN9sP1CQYaqQspXcgr2ubhRvr76PvN0TA7TGRcgEjXj/PySGlEAxzSQZE3ZaWsSxUj8wWN+hM9C54asfXJamqpqmOxZ8SqFu/YFinKfmzSCsMQkvtry1Kxu8jXsq1RDimDloeOKYbIgpcFbZHPH8+BZ8/pYBJkEhY0gbgFY1AK423qEL+4Fz5eYye+RO8EW1rD7fZo4PbpvxH4afAIDe6zYwLaZ2oDrpt4R+SaJEG3tAuE1Xylmpfm+ml3Os9QQb+xeNJTdVilKVII0J0VFKk/Dbod7xhrkh/h51EKOK74XZjnbCjBBx6xDnbd4RoUJaM7pif+sfakuURD39Ys9zWsAChor8CB6mmbsaciVtlABHMV+bFX/zrOZX1gq/9YffafMPJ5Sg/DixUuac8MzvHTpkggENABhaXNW02SEKHD12tvlRz/6YRkdHi5Xr7xdPv7wV+XUyVPl5KnT5Wc/+3lZXFwu3Zyv2LeALQCm73jWA/9nthqKRhRlfJacBYrtI5+dvbcu6+qYP0l9KBslk54S9CeF496y3ngGuR/Shse5lokciQGo9mwaapxnZANDcK6Zez5Jj671Gjmj69FoogWgy9q2msYz8vy8GxZnbn5b7ah6UwQvyFnYPZmImiQ+zx6ghmrMR0qyil45FMeQCnjWvBZ7gtrN+RhWdG7Qcx9FGQpruMZh62tsKAuyEDKZ0PfKH7uqdaMWStWBGwNZp5po9KKiItd1NhZedthnXtzciMjaI3OYBk7TeA7Nv9ec72QTRP9ezaNrfN7nrtl3oboXfp2XpyTZeMz34k+rD5r7Ps0UTP1k1Ry1pfCezpjdXc8nI16Ro6cjCcRf4pQGZgcpx69vImmq+zwXzpgI8UDN0VLKqPJnXBKwIXUO7+uE9ESTd1fnAue6cDxwo716GR4cKpOHJo1xajae82M5pCg2enYshKocfn1Batyd8uTxY9lwup51g48vsEbWA4pf1mZ9d6+sLK+WjU3P0mHNU7/yrA9PHi737t6TcpOh98y7IO4+W+U83PBeeq2oePnCfP3df7h3YJw5xcGCSiYliWEGPDYiwABqAw43/j46PqbCEZsdNSN26ipqeR2A3Ry4J5k9HfuDfQ2mk+xTxa9lVbbiCJ/V3b0yNjpSTpw4WVZXliVvJTCdOXNGaoj7Dx7ptQ4dPixPzXv37imhgD1KAEqW4sDgQCS6ZomQ8J07d05JJRJuGIwezrivZkUqQySHDJXI/MJ8OXL4SDW8hmtdW9tQIkKC4mtvLY8fTwnMJuhxiJL0cN8Wl5YlX8YChCCmwaxt7WV8wpZY8u6Lwdb8DMEIxQZApZs8+FPat5EDlevC/oTX5p7xPDicCXj8PiwMDYrs9GwOFRhhU0KQtUWOO7MK5GJihy1QxYD2QaTnHlYhAsKqeQqNg9aJv0GTHGCXUl4xEsMTEEsguhCyWjo4ECticGhAh876JgOpAZAopvalqKAIgC2OvK6bYUy79bK+avZmK4NtV5+JBYRiRiCvGDAeTMy1AjwxbAlgQYeALD8MLtoX3D7aWucCoPE6HhLziv/GroX7babFXhkbG5dvoKWMPgCfA81j2KA8+uMrB8v55piRUp3QFShtsDmbULIsSymrAH8rRNICxHJQM9Sz0RAvWlnSCMAPNksy2j26rCEzVeIYhVsC5VpPMeAvk1OBUNGcyE6+QFp5Dpvta+/NNt3rVooR9rKaPwZwzTaEcRCWXm32aRcwFdeQiY4Sucq+ytdrlY8bE/mVrBmxCWUtZKlxNlX1PZE/zerJ33VyEsPNKNg04JYhxwDY7WIzCkDTEO19ye2zSOe1u3t71IwjUSE5AlzIwXLcA/tW1mWtIPBahUfY7uSAMlQcGiK7H56vdcVJ7pNYfjWabd26Znkls2+YnwNbOweVhXe0CjgSa+JGxIW8X9wPNbt2sbmiUDeDRAwreWvaB5/CVA3SmFljL1I3edK/+blT7e9qVISaR+l6kwUSYAOAAMMS2Z+eF2Lv3PzBimEeigGun3gCGMUeT/apgX0DD/odWTq5YGJ4mda9CjaaIR16TsR/7d8ofvK1E0TV64gJ7zNBQ31jvhGvC5jrdehiI8G4RoHQYA/lngTEEGt9ZlZJciqqIiRUsRdACTBlY5OByBTnBr2wQKQA5jzxfAIX8mkdlICzFUduhmro8/6emq6si7R1ge3NWgce4iMYwIhrDl9aCnKSYr68h8xQbS6ashBKNtarMp6/z0YFi3V0dEifh/lHYoVKsYcc240BDcqO84s4UcXfAKRzBotAvvDp557Q4JmfZ/aCgXMrUliH3msAPZwhE4cmtPZUbFTFvZmhsKxpxgrQAyTc41lO6MzAMimZ6GylXMeAEdxnFBesSV47bZ2suBiRTzZDN1Odwx4GhFceo3Xp8wISA2ccjTo1HcNKj/tG7NS/qxniQZjkY/j9mzEfKigxYA3wAW6yL7CxzHwwVTesVTU9Iq7C1kzgLZlxGZc9DNbkFuV78oR3nPbvuLGKHQuACmoRwFpyrBxUD1uOOCAP4arB77kefOXnhyzDwOtjx46LyUos4D79/Oc/s4We4nuwMMkNQkGVtpnEzVS+ZUODZ33m9Cmx+yFCHD16WEDW6NhIubOwWGaerfxWBcAXmxV0ckFm8+V++yYFrzDa21uO9PbI7gmVr8/lGB4cnuYCK8LL3IQXEyN8P3eCZd0gOyT4lOAkzz+bt1JXQMrp7ir7AOr7B+X8ifFybHy4bK0tlZHBAQGHC0vPSn2/tdx58KisrG2Vi5cvFWb0lraOMrv4THMqcLeXVerifNlcX1OONj45WR49mrKior21nDh+XNZP9W1burDPNDCZIZU9vbJpYn8xp+LRwwdlfHxUexp247Vr15RbPnjwQPMbGHbb3zdYLl48V376059q3tzVd94u3//+DzQkt6u7R1Z+44cmyvXrN5UnCthSE5y8qEUkKuZU3LhxSw3fXTysA7pjdszYyJjOl4dTj6R0gvVPvMrBr1YQ1qVUcn7oeXv8n5kJLS0GQURIwNZka8s1Dg3Z7h7VYFNTU/HvMMZtK8Q+f/ONy2qQsM5Z/3wdOjSpGKXBxts75dbtW7YIa+FzcRYY+OnodIwlJyE3chO2Q3GK9/cZhapiW4oKvsfZTa1IDiqQmZoDcDMaFewx9h4WfnyPHEgEuVAKAthw3cQsqchCqcK1jowM6oxEHQI4NDLs2YDUTzwPwGYALp4BMYO8itfBGhCSGsqK6Zm5slf3uSpSWHeX6g+r7iCJdeq58pr8DvfBqi0IYOS6B7JSSsKBzgNmANR3Vd+yznku/J1zgWflGWsQ+XJ+xr5yUf6N66eWM5ktfPs72lQ3y76KYe3Uzlvbqlth1fJsUbiwJngPZpFgeazzURYmKAkG9IwF3HV0lNW1Fc+RwV4k1hb3CI91zkaIf+Sz/DxrgsZFrkEBdgwxRikb1rvkHHz2JINo79V8L2mk8F5uzHf7+biEsqIi7Cyz7vA5E0SpIOZInRHKigZhyvmYYr8a3TSA7AwAkK91RD4fJBTWIs9ejgjYXO1CEoJA0K3PnYQEA7otpburpnyIdUPN8u/+O/92qW9vlc8++7ScPXtOSj+IBe+8c00WWtT7x4+f0NlLjOCeHztxpHzwwQdqXn77698sf/PXf63c7t1r7yo+8DzbazUpKTw3yMpE6iiulTjKtYpAsbqm+KKGFASe7m7l78+wQoq8Juu0zImcy4UdbuQbqVo3EcIgK3vLbHXvX+XSkLiUY9tBgPtjYNUkCn7HNWkDtJeiKAiMznNd42o/Rf7MmhTRSPPyZMLq/xND4+dMlELRT9OOZqAtMhPIts0TQ5bbPIsn1onWdFh88jlNVjQQDGbANZAjcr7LAkrr27ZtWKDxPDK3zTqT320WVBiob9Q3/F05gvJN/3ejAdEg+CR+kPWDGijh5OH3aKgqXsyvn2smNP1sVROHeqI5AcnGRNY4IvTE/0XWi5wpn1P189WLPN9E+OI9+PXpzvONCje9hANEXZh10vOv67rVNarfnxwXkgJ2hcRiFA00M7le8jwUBKxhKQSZnxPrk/VEDFYOQwzrbJdyUk3V3d0yMjIqssLjx09MtqExvG6HE0ivxA2ekeJeF8rDeSv+WlsU245MHi6fffqpYq/UGVLCu26y6oj1ars9lIFY449PTPgcI7bSnNzhLHRODj6K9TjnheJaS1tpb+0s8wuzapagCOMzSDGyf6BGtd+XM2ijnDh5XNgV57PcbV43Kn6rfPz1L/0e34FJGIZRVCtoBwCQiWHOAOAwI8BzNFF0p40LhSVBQmy2kCxKVo8lAMkbw76qIYitSp7M+LWCghfkACHBIFHHzxHW0Owcthk1AQgEDcBpBQ/ZJXXLKzh9jDlkxTIiEQufNl4b2RaH3MVLF8Uo0/A1LIJaPOOCw4p/50+CFOwqMTmk8jgQ2PTk8ZNgDcFKsVoABYUOzjYP7OL9CR4kHDQ4ABWWlhbEYKFxQ/NE3dwEhTncgillW5r0ZjRIYksZGNMGgzNx5Z4nO0csmZCeE7A5BEi4ObwNzuScAA9zS6ZGJjDJBhCDKoa7JlMhE4z0lMyDLIG2ZGHkfIMEtKQmCMYjCQmNCWTtG+trpTtAWQo5NahC3tfWiqftgWw1kGxzIMCQAn7o6+pREYLFF16cm3VLchkiJn/r/QOBsZYI2l97fnFR60ksMD0jimf7urtJAxBsf2zWkQazyk5iTwcBBwvXQ0OLZJQ1nIAXh4pZybbByiF5ZlHZk9xJhxNoAUTB9slDOZOZZkstnnMCajrQQ82U4FHaHqUSpJm1kkyY6hnJCldPzpLWnFERaWX190giG4luNiCyGeJkKiW0aaNSKW+iYaF7A9OXzn/YqrFOxHyRSsMNMeA0xYGwGUtVhmzfoujIZC+bZUpgxSBPlUWyO1Ne3JibkkkpkEoystyoMKM8raIACiYPT+p+U7ihqIBVx7OSTHxjoxrQevr0KSUrgB0PHj1SInDp8uUyMztTHgj4GPfArd16+Zv/52/KjRs3tC7Mcre/ciaDxDySJSkLornC881ZGMlItmrEw97UWgmQUQ2/sC+TiiJqhMXlxQr4VuNF3sgHAiOwWCO2qIGVM03qdSVx2L1ksylZ0MQvrdcXM8goLl91jOkaQ62SiTo/S0HBc+b15UENi1lNGcf9bDxk/E5royy6SPTEHls3gzsl6qwPQHwlhWHpY+/5JvUPjPD+fttaRVEgdkqTusbFV13PW2uUYjeUTBToZhpSJNrn2fuxWaYcRVZTE5NrA/QAVJjR0GE3yTx/wMx+NWpCxWEeltUVChkHpYyPj6kQpTBVYwH1iLzNGVQHa8cRQE3DYKrpDKnXS//AgK0xNNytVY18N0FdhFtx5yFwtlKzsoq5Ky4QGjOJuCe8f96nChz4NflMFqgJKuSPvur7L3up5kKr8e8uZin8aarxnMgPsGAgRnMuArCz7sXcZHaVfMpRNLrxLwunAOJZc1hHcXbwGfnd9bXVQv+MeLakxgGe2vbqBkgQO7TTtl5z8wuVNzw5AaAMQBMqGq6f9+MZog4gdgIU8zy8/sw45VmSU3mN249eQI+YZLwvCpmB0tZuxiiFSao0suHC58HOjFyE97FfL7Yznh+GhaIIc6FwdJ7UKfJHFmTEP1aH16gZyXyGHI5Mvqe9E8xHM9Q8y4AXlxJJllpWkal4b8MGJuxxAmhTbAomNeQFN3TMnmVvUyTCEoPhToPTy9EqEH6WfC6HrbrhaGCF9+Z+y25Qz2y7DPYPCGhKkJC8MJlstgBoK9u7MesqGlq5zg3CeMdI8cVstFMn9d4MUeU8IP9SflcOyr05M4F/m6+XNiv0Qr9bk4JXODY0WHr2D8TS99pHFQT7nzXDfTdxoTnu5z7VwFYINU2DLxNpSAa/GxThAS07xU7FPf3cfr0cnRgrtZZ6qbXWy1sXzpX5mafKsZZX1kprR3e5efdhoV6fmJwobR2tpdbdU6Zm5svMwnJp76hpntns9NNSp5iv75YTp06XqcdPpAggp9Z8peUlAQZHDk/47JNdal0AH2pdmhIM4cYrn6G371y7Wh49BMzfK2fPnCkffPCrcuHC2TIyNFT+9qc/L9euXtFenHrytFy+fLFMT89pNgkDuQHhOd8Ypo3STkORK1JXaxkZGdLZhqUszTbuOZ+X+yK1JOr1UP5xfQAQab2S+cvaqi3nAIn5fSlpUUWUlnL06JHy5OkTATT5RdzncwMuHp48pPkZmbcTg7HOJe/gZyBZkc+kMksqd81xaBcYT41FHLX9xb4BEhGCnEe7jjAIyf+l7MaOIxjc3A+u22cWVhi2PeTLAJyJIfLcjvkdzYoM9psU2GEzI9ISwL1ydqt+yYn4zAHcKmQAACAASURBVCho2Jso3zbXN8rgwJBJSJC49g0U8X4on7B88Wwug734gnOdIi91dBpoJ3aGksNno++7SGPMOFhbNznrwMAyzWP+T55tn3urLngdahie/yaMWA0CdtPCVoFWBstiOYBURfew/g1Kt1UxdStfWUMbm45Vsuzc2JRayOeIm78mMtm+kWvR/MOuLs/ZWl4OdVTkODFjAvtE6nHA+qxdlJuIUBLkqDrOCF2K5QP9fVIhVfExFLEiu6BsBPCGJBdzMah5ycH4UjNg1+eMB3LbstGqIMcQ1p7Bc4PbrL1s6GcemedF5iZ8eCvlwupR54gbNVxTzhuSmu9gX2ukrxcViTIdq1zqtovhWnOYezL/+anvfPubpbe7psYm8ZBmKddKg5P9yLM4cvSonhNqC0DDw0cny4cfflg629rL195/v/zyF7/QPvrq+18tn12/UTY3ttWoQFGB9RNrhrOfz6F65+BAQOe1a++U6SdP9Qy5t6zv3u7usgVGAvkhbAsT3M1cOxUPvjce8ru7Y0cHag5+PlWfOcsvrcua7TBzT9iSy9aXOWuGe8P1pJLA6vDwKW2yUFQ9GvUB5EXNrIiaTjauoXRONVJ+ltyDqi/jRJbbRDSosI1ib0p5JOJJgPBhDaxaOt6b50ncoAnH/kkbYWZfSjmkLofjlOtn76n8ckn0YqMiGjLRQHA61FAyZNxTk1OkXc/X0k801VjZqHgxf8j74B9/UYHgn87GRvO/N+M1L3uNZiwor7lBbvxiFlM9j+oSGqTVV+U8zv/9MbNR9TJVhXEo37MkkbmRYqcO6l6TYFuUFxMf+HHwSP50o5Gmo5vvSbomztvdIvAQxTzb8kGAIBZD5hKRrLVdpGvW0NDgsGKx1IAxQ0eNeA2Ox9Jxt5w4drw8fTJdkdeoO1O1IfIBaqx2yF9cmwl6mk+lJqrjM0wdPqdszKWm2lLuABGAeNRd6xZhkdcl7+ScY3/QwJ+Zngnr87A6pcbraJf9nNTQrxsVr1qWr7//D/UOjO6a2aKAFcz7BK4EhKtQ29OMATYKDFPLTj1EkWRVQT+HKockUPMV2Nh4wAeIq4RmH5Zjpw5LNiUbEaAPux9eDw9hClAAY36OkEjxTSNA/pK9vWJnwHSYY+BldKNzgJ2GN4UigYR3dGxUr0sCnGz5QxMTujb8aDMp4lpg4JJs8HMcvgAS2C35gCHqmq1Dgid7jWewJ1tlTzU3Oy/Ac2R4RMHTVkhWP+RgZgIyBZZnUgBamJFIkSH5MQNhYSaE3Y1tgOyhBzDHNSVjnYJHoARzKrBiCKCA56gBmRW4lYO7La/Uc055ZjCEE4DzYW0WRHXAvWD11HxY81piS+IrT2EbjSkzOcwAIsmgUQGwRGLP54dt5NkFdXWOKTxhwM3OzwlkEEN9Z6cMD1jtoKYYACoF3M6ODhgNFiPRbRpAx/rCEozkXgloJE3A5MnMzuaKLTsAFPsNEgZrnc/P2iBpheHTzERISWyqJtRJl8qluVFhFUomOTnYrPl7VRMp7rfYZQx1C39FeR0K+OeZNXs/N2ygtG5VPDbsf5T0h2xSahN80qNZ4kGD9WjWmX3iBCElrC4+XdxZ6aRheny2DG4vJGF8G8a2fBuDxaQEJe2qePVQa6nQENhuC5osdtLj2qwqMxRVbIn5vSurltw/2dCQdDbmH9iOyvfITTerOYgvmQCRHPNMiVmnTp4sb771luTexC68lH/y058oeZXvaRTbDN389je/pWKd5OhvfvAD/Xns2LEytzAnoOLY0WPlD7/7XQ3s/PN//edixnlIq4tprpd1SsGdyRrgKntcNi+w+Wtm89uiJIAxlAXsEOwGxArZ1n1Lb2g+uwCBNgPpAM+yJ4rGEj9PQiMGRljq8fmRukpZAGBOwyKKj0yEBXpHo+ML59mvUVRUjYpk6kSGyn5XPArvZlnRBYPadnf8u1nkntVi1YfPo2S/oWKx/3V60WqYJvFSDD0D/Kwf2QzGHuA9iTUJKAG+KBkPQIB9XTULgoGVoCTfF4AM0x1GowDmhvdufl7H6rRRiv0TgzVp0s4vLFg5ouacbW8aQ95zgJzuULQRfK9IpIn3NJ2zIc36kCIl1HRqVKSnbQIGB8WWZPW61oX90/G4dvNLnv5xHQxiy2YqDHw+i4t9PzMBLznNu4kh11wENa+RFxsTzX9vLt6qMyg7bS9JnF7VqKBBDFsR32czcAliVk6ybtnffJlBic0coDw+5HU1D92Msqcs5xbgUVokwGIGkITRyd5kyC3xAC9znr2s8lRkM7B8UH72AsqxGtvfE8OL1yQ30hkrtVarGFi8vwbjylYThjPMY+wSsXRw3kM+Y4KCAam8T3iud3S2iYChGSYtDAX30FnuAaxeYgyFDq/Jz3M9GvIaajoUisQlMYEBLGIOATmWHoPsDp2TcN0qEEOlAFHElpMuFp0vpa93zL+SKotYRS7n9cNrwfLO5no9bCf4N653ZXW5UhrpfTUU15ZCNCoYDriza7JGNk1oLK2srVYN9FRBZcOzmsUSxIskz3iOwZaLQSmmYvCmGPF+tsRr9guvRRyXJVZa06lRcUoNIXI+YtfgQJ9sQFu7a+XTp7MvWcW/+bdeagP1W9o9Nb/r+dHhsrvB+bUlxqCtbkzaaFYtVg1geZ17Zo6sw4L5qrwzbVtC7ZjbV/uLtQMpYQ+1IHale+XE0cNlbLCvLDx5VC6dOVZG+nvL2sqyzqNtcuL27jKvodlt5dDhCZ2pzK64++hpWd9isGm7cnesn/Y1d6qtMESS4bPEcPvtc07YkpU4AIt+aXHZw6sB5DuwIt3XMPHTp0+Uzz+/rpkMKKCv37hVrr19ReA8A5ppRPEn7Ogzp09rb3OuM98OktONm7fEoKbBx3warkG5ioZHM0PBakkDdVbL0oxLNazUBj29ulfMqGANbsiWwo1j1iGDdqkdiAWy6JPNiUFtnhfg/CLszi2Y7p7DlTlL7iENAW6zuko5M3ncLqx0M/s3BARHPdMUg2mcnDh+omxubUiVLNY0AAiNhXg/1xU+7wRS7hG/sMxwXICZrwGlEB5iRleqEGzZaTsXkYwyqxQxwGeRBriHMo7Xk8pBuZutMtxEs60Hqh2a0uRj9+/eVRMpZ0U4+7Yy9WC/LvUNM0pokBjoct5LveX5LCYiiJzXZCOc1hycM3rPGJSe9q7Ud37mVgDnvCf2WJ6fVuW5eSOFTHuHPiPrglo2LT+lrA0/dudAzPJw/p9nD7MdZNe1vqEa1ffdZwp7jvXCPVP9gnKgvhf2ITRPyBd9XlJv5mBh1iUgWqqok0SRqrjMz1B+6t6Rw+w5p0j1rvJ6DQb3AFjVZdhOavZAu54R18IZyH1ZXFyqZp/09nTrjOaLNcvaz/yDe8c+yVxCsbmyVHSTVY2P3Z1wAUBRa7IKc6ySWGF7JDft3OhoUfOKvaAzMRpFXOPY+LjWNrFes5RaWsqbb1wq87PT2h+cS59++qnUPNeuvSuXBog0eMeT5z998kTKqrFDY+X2rZta0++9+5Xy0x//ROfd17729XL9xk2t6VpXj/LL+w8e6nNwf2moqdkfA8pPnzpZLl64qPOfpusqczmpsVpbyuzioixg+ExyvggbzAaphya0G5FqVGwT+wHNuaeu0UWSg0BZ5YfOFfV8QynADapyMuFEgUDTtJPCy0OLlfcEQTJzLeUCUedyPtgKyqA0DXM32PynrNKqAcg5H2O/dCgWus7M+SEiFeyiqPWsL9UT8exttxyWwiIptahxTaOJZ4OdFjdcpEjWg9aqI5Jim+pIrcLqOPVHcA7Z/JVxyUqshqWxZpFq5mDMoEt7deJFWMA2vfwXGhGvakxkbpmfNf+e15Q5WuIWmYvx8xWh9CVNEv1eEKVezFzy7H++V+Iz4GVf2ZBwM9HqmOYZmRXeZPaobadi1g/XmE4SPFvZw+3YykwWr7Jb3laewbrmvGQtcd7bsrKZWBVzKJKoKtvlWhD42uxEgpIobN+4bvYe8Yh6wKQvn+0Qubiu7a3NUuvokg2hmp+aXeTXohECOYYZbtgTUm8rfu9agcZ1ijy2SzM9zrOYFwmpyupGWxjyO8QgMwxNoiQeaf6tciBqOc8g5TPvctZpXmjtdaPiN0+9X//kP5Q7MFK3zyabimRGhWgMnJTlkWSHFAmDYq6wmQgKzUOTxTzr6BCIQOdfktRQK4hVLf9s2Fn2ieOgtBenJb9ifyAx7eqSBGp7d0sJwMjQsGSOvV09KpbFNmhrU6Hx4NHDMs8wKQDrOByzqcJ1kIhxGFPIc5hzzQ/uP1CgGh8bV4CTdJc5ByGFTQYvYDdNixwKJ3/E8OQn8PQEC/Px1BMBBsePH5e83oGqR0D6/MKcmi6LC0sKqmnpwH1KP3WB4wBmMWRbCa0YgTwHDvi2YJngQWrvWYoGAmn6cotBCNAZMymctFleSfOn+QDT0dtkU+Qz196haT3kJDEP6TjcwiLEvtQGUVz8uEFBIM+mlAjZYR0E4xyAiHtN8e8EqaVMTlrmJklmS3tZXd+Q+oIiEHADmyuUDgKvw4ecAwUAisJyZW0lAHkGjJlpLOuGel2yWZIDDRYLazF5MmtuggcQc7/5kwQNxitMf3nK0r3e2FCiTVE39fixpOkqRMPD17cmpJqVrVIjUZMEsMXgua10zFyu0p7IfSg801pLDGAGjcJ+icS8SkBiP9qn0IPu09M3h6flTI4qUQoWAe8BS5XilcGAZrxQ/JhhbUC9TYUczLBk4TQAKTNUXgQsG7HNr5GKDxXpAR5W/x2MV5gIsJP18zxXsXGiYSe/fjcJzDyxHz0FHU0rsWjSJg7Pcq7JEoHnkkeB9eVA+53mnofPMcfEzxAl1Pvvv1+OHj1qq7bNzfLDH/5Aw/FgyZJ0o4DiPrH33712zYNz1zfKRx9/pMYCv4MF3KHJyXL50qUyOXm4/PN//n+o6YlfJPcCIJFEB9CYL5o5qLM+++wzFWupKOO5W55qcFJNwmj6imEZRQUxcmNtXcm2rKAYiru1oWKHZ8Nny2Sdeyu/9lBvSTGAjZqaGyR8yKYZMu+93VyAOBp8+a/nuD7NSXCsfM9Dsb98Mvv9LgmI1a3IyQIpcmDuGV8w3amNrEIyyKCvVgM1fAbbv7WIUes451gs4BhgNVQoYpMGQ1NNubZ2g2xK5N28ADRSIb8LELwWCWlzo6Kh3MhYwr1MZRWNDdSBmm+RsUJxs1UAciaXDfDFHrEGgfndAc3WsKLCxbj+FBsrnhDFVMQNwHMAItsFAEY5wRUxICzCMoH30GR70FsFRkxvSPUddxoWW1UcCvD9VY2K5p97WZGlWBOxLdfdq4qxVzUqeI/RkSHlELJNC0CIJiPPi/1Pg4diwSx/3yuRI9ppiNOIcGxXnOf5AxxtbsraEtZSV3dNDaHppzOljd/B97Xy17UaQSxmFaJ6MtpXAAwCKMM+LeXgLg5bxNTMxgnX2JwT8GwAaMxEtgVIDjQlhnDNgKVeHwZI8asnX1teXlLjBgCdNacYKIAoLB73DBDyf/K5BKAUO8I6zkiNCQpiZEJCURPwQKQMQJBsumVukUBUKjucN9rySudHzq8I24n2dubOWEnKvdNcnLT3Y+9o3gqxE3KGQbyWNlv5cKaTF6wqDhjs5DymgGWvshbEqmzh3hgoZj1cvHBezwo29I3rn4cVBFY2MKOtCRFgvLFhNQmWlQxXhxxC0zmunQs9fuy4rmt2BjZbq3yFGeaL/dOnc3NlKyzovnz09G80mhW/u5KC16u1t5ezDJBdWVOTgjXnWBlzsaQQchGcLNxUrwBGwwqGZcheEMM9592o0W7FDGeLbPZiSCU5v6xb2lvL4GBPOT15qJTN1TLSWysdLS3l8JHJcuv2vdLSXit9A8Nl6tHjcvbs+TI+OVF+8atfltFDk+XB45nS2d3L0DLH5PpO6e/rKYsLC/KYX1vfiLk75EKescD5yNkuRW0MCmaWDMqJb3zrW7JyYoA2a+bWrVvlrbeulJnpaf0samv20KOHT8p3vv2N8tln12U79r3vfbd89NFHypewEPvh3/5E9g3DI6NlYQEwtU2qbDPo8aneLYcmJ1SP3L//MOxLyJMNNpObTR4+rLoIkJO6AYIRjF+aZ9RVV956S1ZUPCviuI64VOdGw4FYRk1EI5Y4CPgu9QZe2WosNUgb7CWRYAA0ktmKlUrOJKH+ijkI/CyDlY8cmSwzM0/L3BwMTuoI576aWxAqK/IgzVagplNjs1/7j7+Lsby1pRisQaSaHWMLjlRvc06lhYyUurFpZJtJTiCLJBO8NJi6s0PnMPuRa+feUU8QG7HwINe6/+B+2dne0n3oqnWXjg4Y8AwZ3dVskgvnz5WVlSXVpyz7gYEh1TAw2m2BZMtHrgFQGECT9+Cz8zs0V03yMBFup26bPdZcDgIXQC773h3Zlvg52wFASniUaEGu4nlnDcwzIt7KbQDWOp//gCa5FWNSX+hccdODwdSsPc4i4i33nGZ9rdt5Ho12cmnbR65rDRmuxebGln7kPdSp7P1sQsveVip+hpyjNHA9IvAQkHBnW3N6RC7E3jRnxoUqH2IY8SLPG53ROotay/DwiOIINbfIEkGCIH+2EqYujIHab35+rhqi6xqABr5t6BIOz+ZYRbszIV4WoCIqdtUqTEHXgwKouydyIp+xxI9UGlKXr61vlhOnTpXTp0+Xn/74R4XHBTB59e0r5c7t2zqfT548obOFXP7q1avlww9/qcbR2bNnKvIj+MTI+Ei5efOm1ubZ06fLxx9/XPZ298vXvv71cvfu/fJsda0MDo+U6enZMjM7J7s1nUcx14E1NTDQr88DLsFZxh69e/tOuXf/nmZkzS+tlPGJQ4oBrFEa0TRSNDNUpBZbLJHHcn6ybgQcB2Cqdl4A78JnQhktO03VzM4xk4zjlL2R+/LXbIJ6nbouM0BtNnvm56lSyNcS9lHlvH6qOfNNSpogO6bKnjPfDQ89ecUB1cQB2BJHspFgK1nvaT6DZrLIOg6Au8ezBEJNncQfKdoD5LYNZYNs6DhsUD2b0Q0CoBsSxlUa9zMbG/qcUZPkjEX2Teb+z63jIBW6WeOZkdr3Ct7PE4cyz0g1eubfzTn1c3VZ/kI2VKI5IBJuEIl5zyRv2c2jYXn7xbzG94j7kRag2XBUIy1+IckyVtW89Io834G5NKEyECktbNtQDxGfZDsoRYUVYOS85LOoDTjD2Ntu1rpJrub/QTaOqK+Ik8wz2haZmCY1c9/2aY7TnAA/I8fZc92EKk82id3d2oeKi8JJcJ0xjqWGInbEkbOalNMqxRZqapoL5M7cJ7BK8CvWYzYPHbFcu6bdGucM50BiI6xd1aCtWI2S47Rrbzx+8kS1m22mTNIitxAB5bWi4rdNw1//3u/rHThKYRaSfhJgd1btW0jC5wPAgCUMFgpU5I0U9ckoJ3mGBccBPjc/Z6A4hi+y7TUECYuJNgNo9qGzbQXvx8FEEAdQPHzksNgCU1MPVbxOThzS92enZ3SdI6NjpaPWKWuG9S0XLQKpdTh1VvJcvISVgJVSLl66pIKGZDE9WhmuSPLMgcLm5+dQWhB0OfQPTR4SKxXm1NLyYunt92wNghEDKrODTpIoefKe7RtocMi2Y4sBhmvyOuUzA7oRqCTBDxaOJNAxm4BkIg8nDbrVfXEDQOAWAGSwtNOPz0O1D3SdYoky1yIknWKQM7Mi5hJwSCRDyIdZShRTAVB1KCpgPZPbbFw0d9SVxMCGkJrCID/Xx8/QfSb55sCggOQ+A7QQ9El0BgbNPgVUbFVi76FWGt6ooUKoS3yY83Mw0QysFzUp8A/N4XTcA+49DRpYrTS0LLE26OeirN2ewlGgCUxqaRELCwaSi6YWgUWsTdj2TvLNuOVatGab/B0NmoYMvnHrwqswZiJEIqZEpjqjo2kRDA1nOX62zbY5SmRCmZCApC1xYpgYAHgUEgaA/SycCMbwXSW+BiQzCeU+WmnRsO5oZrv5cqK10qysiQDWDFSaDGEAV1qMSPD4/WRVKIENBitrvCEbtz2U1TfB4MkmjtjuKeV2Qyfl0JkUUhTZHKlhRaCGiQbZMgvHll6d2DPApKjVNLQTwIlmAffASh0sypg/saemBWuP9Yw9wLWr7yjhZU+zx59OT5fDk5NqhACkscf/9sc/FiMK9dDbV65ozVAIskdt3XBQuhgKvb8v1QWMze7umuIln1vM/g7PoJFiIp6pQPR2GH+bSlxYsxTNPEgSIF6XPQ47W8z7YColcMia8qwJmlUGHaXukj2bmXXgrwb2gi0UhUjTYv3Sx1ZzKuqZCFyH7YWalXe8cErNG/YvXgcGOUsF1hC3U83EtelMUvKeSbaVKIpq8gtNZrgZa0o8g+kqVpcKtWBV51yXYJjlemR2Dc8G66i0H1DBEq+dDTyvdQPBGb8B9QAyOWMqJnLsjyxCkv1prLDxDPhcMHl45smuV5MmGwvRlFeDORql3EcXl3UVtfiWipUp4MVKirRwyevOz5GfqVHHpPLADZ/c7y/++aqF0cz0yp9pbjxkMfmyn3vZzzfe50ADdfl8sn4CFCduwJZDcbm8JKZUrn831X0GsCcBldjXabEAkFbr7NLZmSCU/HC3aFpM6pnfu/tATQrZMAUrKm0waP5SpDseW1bO79BIJ29hH/OeZvr6bMn76YHxzrtokPJFzsHPcX1SSwQTkn/nXuXvJ8uUz8rvwwLPZ5hF1d7+bjBCzdLNpj0e6iJjMMPk2TPbiFEkxlmgZxM2bbIZ4/qGh3VdC4uLMazcNk1iBTpy6E/UPXnusP+k3mMvYo/ZCnjlgYhSmanApIBrLTuAcwJU9ws7mDjNmdXT16UBgQBchi8PyqGJyfJY1jebUkcoD5I/Os+AItMWd1w7uRZWOfx99dmzMjdrG0flCjCPAR6DSSolFsBrKDGlQmoCLbhfsIIBrfCMB2Rkf/f39pbevu6yvLdXHi0tf+lY+eIvnPrm98rXe5+U/+3PbvzOr3UYaySsEVbXBTZrtgfWNFW8tw2Fcg7lWR70i7KYPJf7SR6ajD6arzABOdsAAdSAo1iP5oQALAGFbWWnvleOHBkuVy+eLdtL82Xh0ZPyzpVLZR2ySnd3eTKzULq7+8vNG7f1zM9eOFs2ueedtbKxs1/mNMOi2PZzZbksLy7YmnVsokzPktdvl4FB9tVBmZ+d17Nkzzqvc8zDCoE5dxOTh3QekIuzLjh3sW2kKcAgbogH58+dK7/64JcCpycmxssvPviwXHnzsuLNJ59+Xr75rfdlSzr16Ek5fe58+fnPf1XWgtBitR05cFsZGh5R3oJtrVSO2FV0OQdnn3HvuP/sdYDSWhf2TzDQbetouwhsjAZ1XTwf9q8a2zFo2nZEdb0W5yJEG2bqadBzqDKrWK1ckMfUYBsnuMQ/SN0aoJLsKXZ3ytGjk9o3n39+o+xsuxGxp/PHyjQaFFKKyObThB9qJOIc9521A1BObmSbmIZXPLmUQMK95+emJTGGuk6zMKI2ARy3L36bFBSsZeeFXrvK4Xt61KzgTJiaeqS/q7HWVpNFTHtHa1lfXS4nTxwvz54tKS4yzB1ACgU8rHbek2dInqe5GuRsaoZs6zPzPDgnWIPccwGNzNfb3ZW6zk1A9gZzg7YijnuodHNuJQVmgIIoUWiWZ26p84zcrxV2rlUfHu4MQ3e9jAyP6mxgzZBXMGxZCrQgBhFf8VPXntxlTsamaiKrrK1g5llT76j22j/QuZgkiLRLFTt3e0efXxa0UsI4b5T1sYCxZjDaAK5nLno8XIOwFCz1mHkFQQ1AkZy1s7NLOa8aw5qXY7s95kewRmVNuLXteSM7tkBRHRSgscBskUpMtLT1oetF1oeUOKGOSaU21wfRj+cmxT3qD9k5W3G4ubNbLl9+q0wcOlQePbxX1pYXy8hgn9RWKKrYYwzQpm4HK6EZ9cmnH5d5FFtnTisWPp6aKiNjo2V4dFRNUUDONy5dKj/96c+0bv7gva+Wm7fvqOHa09tflpefidGNTDFnSNJCZ22wFohxNGr4bG+9+YZq4dnZ6XLz9t2yvmVbSs+cMPEoZy5VCgeRRMP6uJikIuC3spXOOV5uQKQDhGpJNQ1rakCyJip7m5hBqFoiwFZej3xLCvxofiQhRbVt4AXZqMimhkmNxpcSvFdMyuHOENhi/pzcOeL80nuETWv1e6muF95klbkIF9GkzSHj2fAiv0mb5bSmCu5mFXMrDCSaeCbHRd4TxY7fP+QI1byJJtVpzPrkc6ayWfV3KFOyucDrJDaUebLqdRQlYROX8eRleXTm1Hq9VzDOHO9z/9qCNN9XzaAgmOSe4HqtXHzJC0YOqBiiHNjPXq8X+UDmvEleeenLRBNIMTBmVCjH6usvvd3E3LUg2kC89RwIv64xBP6UleLmZtneBbPh32mGmtijhtkeNTK2c8wp2StHjxwpM09nyxbrSZZMdmmQzRgY1o4VFDRMOKvlwNAb7jE6L2x9SIyleWJyVF3xX6qMUINxreub6yJApUMF56VsjsmJybvAD1WvRbPkYF/EJqn9UFB3mDDF+1H7S/Hf79ihGZWa+4aKDpX27utGxe+cPb9+gd+7O3Cuf0DsYYFZAlbNrtfhFrY/9nGsK0kjYcP+ia8E2ki+AMX5fTaqkwV3hUmY0vs4AWFJXOXFiAWDB6DxOzQ6kEAheaUYIXj09/SWnS0D32KjEAA6OsryyrOysr7m64hGAXkMSSPJLQcnCQzvjY+8GDmtlp1ircHfSfgMRBvMHR0ZrYBTPidgJR6U6tCSoGEL0UkDp6Ykhd8HYxoahtG4ovtDMoYv+LOlJYGZFLYUzbwW/sYEnwSe1UTA5iR8mElKxJiOYbhpheKf9xBKApYY9VGA2HKp4YWfgyA1j0OBz7ND8sCwvDGX4fNdbg6KBgBvror/nodzMCT0fXuzkszrqz1rXQAAIABJREFUWsKDUplqi5mKJIXMAwARBRiBdcqzJpgy/FANGYb97e6IlSLZsEAPJy5iRmD/Faw/DfdSwuqkXoNyGd7Y06P7ztf8wqLASh34wfKgccKXiz7fABpMgDb49lJkJXBCMoQKATUFbBirXEL5Es/qC8mCGBUG6q2osLw171216ZvAHe0PqY0sHU/bpmZlaSb8yXT1nnNzLxOKZKF5z7oBmMlHAqyVbU02EJKQHt6cKqA00Mys/lweTtrC9iEWTTNjwwVLeJKG5ZPtTQK8zWQymBRcK0VKlcjCvo0EMEFFbpyHSIeX474ZZfJyrhg+zHCwj7DzwwR6W8VMouhETcRPvH3lTQFVJB4Xzp/X8kTZAbDLYMLuHlQ9RQzFu3fulFOnTuvfALFgTsDMovk1eehwOXnypHnqrUWADkzNX/3qVxWbG6YGKiLWItJQGJOw/nr7B8q//ou/KFNTj1UoEjc1DwOv7YF+/RwWK+xvsfgAnYk3B25Can1EQ9PMD7MZE5Tl3wEO8r5n4ujil4ahFTu5HwxONRo8X3jmLzmlnJu/nBGTz9Ppe/OXm6BqxoRHq4opxT3LVnnJbGqbHWS2SjLfeW1YeH77jGPRpMpGGftKTZfGEHZ+DzBnmRkVgCUpSY/1pIIq7MJy3WdSTvLLc+N6aLDKGiKa6llQZYOiuchgv7lxiy92n+yD1HDNJkUohZzQe926YR8s9JDYA6bhnZv2Xh7Gl8WcGxvNiiWurburR2cmZzmgHPJjgeEwHzvMiuTnHBOSDaUrq86HjGsuej2kvDo3XpC8v2SJVD/7fIxovEa+fr7my37u1f92oGc8ONjnQXJhryYAJRpw7BGSd2YHyPd1e0vkimTf8RE4u1OVkkU5r8Gsi6PHjsiWBXAcFdXszJwCuwpcWKDRPOT9Yd0CJlqOXtc1sYenp59Wt4bXZR2xB8XKxR6mYhv6DKMRwTlnr912Kw2j6cSzSnCzaugG601NqrCxosFPnHLh69lZBo5adD6LVRvDKQ3k+gyRqiEHHTY14cgplPPFPA8UqszeILdKkCo/R3Y80+M4i1QCgQCkdisWWkqbCk/iv+24PAzYUbwIlOHZEKdR0nr+mJV2gM68N1ZuPBfOCuZHOc907FdhLPtBlCMwzbfFTpblAOpJKQDMGuVLs9VqqGzIF2nKmVAjr+s4r9QAjjkMMPJZI1LGFOafMA+lpgK0b3Cg/PLxk1dtiX8j3788NqacamNjy8MbseWU3QXsUg+cJW8UsBDrOk9+K4QGVPhjz1GxIkWmoK6nyRb3XUxIxzCA9u6uzlLfr5dTJyZLb1spR4b6S0H9Rx1Q6yyTx0+WT67fLEMjY+X6pzf0/EfGRkonvvGdXeXe1NOy+Ix5AJ3l7Jmz5cH9u4UIyjOhGfFw6rHWcv9Aj/zJUVpw3dgw8pwBWKefPi39g0M6V7CHRQkB2/jxk6flnatXy+07d5STM5fi088+K28zdH1nV99/7yvvljt37iqXxxpq6vFUWdtYkQoTq8GVtY0y/XS+rG9sqVWM3RnxnhzTtnv2gWdvSs0WxBEaeX4GrnXYEyKoyNIwlI74+NcN2Kqxp9iyIwYo6zQbrrAsyV957fGxUe2FVMFbwWVyiPMDP98KIAzwnH9Pa6m0XuQ1aHJevnxJa2VmZk55O8oyA1covgC8FaUFjnTUaGi6US7CV1gVJcBNfFGNIgXXvsHXYuCcvYU1kOaZxUw57o9V8vYbN/mFNYf1Yc1kM+ylYh1DduIsP3nqhJ7D1KMpxUyaIaLvtJB7tJTx0ZEyOzujZ0KjlNl4KF07O03Oo9mpvKzPsT2V43l+i0whdaOVv+Si2GSlxRJnLw2aBOqwIOO18twmrqC88WwOq9KpuSvCQihDyRtUHxObNjZVV1ptvqrkqr2VZtam7HJNTqJeQZGzF7m1ZzY4l/EakIoc8gRKCpQbsJDleGBgOwkxslepBtBiV2rlfOaVnCtp72sbnmZ1aLL4nTdUMyJiTqBtRdvkuoCiUR7xGhqNig3VDRapdmXgHMDuk8G5mffxPVnzyTYsCDD1PTV1uD7NehNT3hZSYspLje86UEplkXVMmrRVHY2hmAGGSmS/lLPnL5TTp8+U9taiBteTh/elZrh//4Hu67lz58qtm7dU1545c7oszs+Xu3fvlmPHj5W1lVWpQSBbtnXWyo2bN8T8fufq2+X73/++mgxvX70m1RbrC2s6gbDkglKZU+PjbLGlc7APW+2WUmpigu9qRgjKzytvvlV+8OMfl6cz83od9gtnKWsm2ftJCCNW8MXvGwR3TZekOO037U+aNla/KD4R+1Hn0NSLOZ4iJEZDQbm65A227vGsCTcHWGuyMo5ZNyIuxJydbDToXG0aKp31b/4O18W6BMfQnAzZcJrYmQ2rrIPdgHczLfPznJXFZ1MuEYoiEyyNXSkPzK5FWlyrHnWtER8t1qDzNb9nWnM27OwS7NccnahTTIK1dXqjecN+SlKi3zzVGqmgqHRDYZ3keq+Rjyee05wrN5o1Dfupl1VrJovldYd9WiiOUvGcr2vczueJv55/Rcg6eS1Ciaj1RARzfORLsaOpafGyZCjXosgx8Tn5PIMoirAO39xQPKF2pmbmTOScN9luX2eBrJH2aBSs6Uxpa6+V+q7XNufV3h6kZXIZ5l62lLfferv8+G9/UljFJRphrD3WGmcBKm0UnCbzmPzGsyXWcvZqxpysm5mNYUwrz1jyca6HPSRLKuyJwz6QJw7GCQZBrE3CM/sTRSA1BHsQxYRmtUIqVTPVjiKcI4sLi4rlsncOtd7qimf16Sm9VlT8G8m5X7/p3+MdeGtsPAZ/behwJJHRULCQuJKocBCpaw+LZGenbO6YKSxbkRg6qmAaiXh6JrLp3c33YZbAKYcOG5nNxvcpjPgi6YMVsrqxLhUDSejRw0fKQF9/mXo4pYJ7eGSk9A8NaVDp4tJi6ezqVsAgWAFKKMnXYLRugeEJPrnzad9vGDir62tleXFJwULD0EqrGFwcYEp0QmL8bBVAwsx6mPkkAiQfBC8CCYkPw0+xfpIFEXLXgz1ZBgFUAa5Mos5gYFn4/hNQ0xNZB4wSBDeHdCAFqKhhlvgrbyHtfCYJo5PGkF/izxseqGJ15rA1APxgqfu50VE2KJyJX5VMxFwEHlF21N2t13FVvVce2j4QDYIYnDDLOAsZfCY5z0hu+FmeMw2bfayiZN80oHtF04bPjFc+/7d0j8/TVrY2zErifWgi2F6Ag6GuxAnwgwGfSvaCMTQ2PqYEi+HnFOMJdHNtAEQGPNdcICDZRure3aNEF3YMCSPvLZ/xlVXdbw6CVMAAbOjQCqTDUkazEcRuDpDRvoE+07k2P6vmDdxQYrhRkUlDzAWJ+5o5gfRNoVRJBkizWsFNDid9WUx5nRnsT+VLc7MqQdaUt7pBGesq2PW5ZxP0zg/xHLgoBpVB1mRq5/pyEmhUyEmcmRayiwgQNBVZLqRdAFo1YskyXx1tZvaarWNbKAGpwUwTAB0eyVozUozY4/HM6ZPl/NmzZZZZNKWoyLh7956SEFvVDamxARBOos+awBZOnxFfyJ5eJdw//NEPy7e+8W0xLpV8drSLaf+Xf/mXstTimxTbNC+5/vf/4H1dq60DusvjmenyL//VnwlAI/64sHJxCcBCkwQ1V6rA9Px2zfzKRlE2dOTnHImm2EhRrDYzbDIxtAIo1BNNjTuDiY1GhRoDsURfQcSJuPGKRkWAornK86fwys51IVltsLv4/Kmi43dyUJ+HRmeiD2PFyhGejxsljUZFXFB0KAza4p+ciT+fif1LQ1vFUbB2sJfxGnV8UUEUA/5ctNnShLOIGIo6Lhvt/F7zOk/gP++9QF9ZI1oFxvlkUMKFjfZtk72XmH/s0YhvCfLKAgGAkWZ9+PPyvrn+3aR0s0KMeAEuXQIeYQrBPMXWIVn7BqUMxvr6G7Ltxr3IJ+/XTkA6n2nGvVelInkPqjUQRWhzIyfjzIs/+6rXfC5qEk9hKPd0CwDiSzNP8FgOkgVWNZwRMKA0F4bfYd6PhsC6mPZwSANrGqYqj3nPJZBSo421ZMIDVkIARNwz2MUgZqwPrFZWV5+pWdjeZqsPmt4ALQvzC1o/9qz3PItkUZNbkT/xc9mIp1HBz8OMerFRwX0SoB5NA89kcNOS9ck1G3CC4bUnVZeHg3u5s68487IxkdYKNFk5l23nZK9oWxFG0yAaFZkzABhjxQm7zPesvXinAe47f9EQ+lBCiUgQzRAUFaws2L9iZWqQZ6q6HPe7w8arj6G//FuB+Qprvt9ECCy9gqlNrjU9MyOQSwOTAeFa28rGtgky/BzPlHt99MhhkSQoAGm07OxsKc8jx9Rg8ojBxB2AFA3vBeCLPULOyDrh+dKo2Nrc0LwDGK7sDwrn/r7eMjg0UOZ2dsqT5We/yVL+e/+Zw0NDZbgdEH8x4ggWJzSwOFsp2H1OVmqrOKfTrkt2PVK6Os/H8iBndtiRMCwuiMeKrT7re3u7Pcy+1Et7y345fWisnDo8UVbnZsr045ly7NTRsn1QyuzSszI2fqhMP50tPHMaqTsweFvby4NHT8vuQWvZ2tktZ06fKUvMZNhY154+fepMuXPvvtTJpXVfPvMiNoS1x97unuaKkcdx7tK0ffz0aVl+tqrn9/Enn5djRyeVU5IHfO+73ym3bt9WbsxgbcBIco9Tp0+VuZnZsrWxUS6/ealMzzwtCwvzZXR8oswvLJWN9Z2yr/aJmZedXR1lfZ25fV2KCaynbH6xmmkiArBUIF1rq6zbIErArG6Oy8QN9jn7AoYk+1c2hAEsO5/CvrRdrysFaA5QpuFWzXLwUGSzZxszSTKPELszmakiD21rj5K+EieOnzym3AsQ1goG57mAR6wb5ttorg+Nx86GQoqajmZiDowGFBcLFoCeuQuwTVs7qlomVQfUTcT1pcUlsYf1/VR41bDlWStjYxNal4DB5AYmqDG7i+HILZrhQQzjNViXUu+jvOpsK6PDQ8qztjex3SOvKFIIUSfSXELlynnL63Nf1GxCIYKNVXePPi/fk+Joa0NNAYAsPh/XsvKMNT0eNoAoZ1zX+pzZ8QBXzRwhLxksjx49FODFulY8LC3ls08/LW++9aYVagBzXV1lfn6hPJ1+IltRLPBQR6E2eLbMeotB4MTQ7m4P2sZ3PezYXMFZyUZzhrgohe6m/dRVwzWRwjIX4hpd21uxVlnlCvDlbFwPtaJ/n/OVc5H61KQJgLw2nT+2OGOtMP+xS78vIpDymQ7db2KLmvWra4qp2XzOZg3vz2skGztZ51wjOTIzJ7JOztqYM5PQZMa190DmW5xJUumhrCC2SYHVqWlnsLDfefdaGRroL7X2lrK1jmpppPzsZz9XLXXtnXdkA8U+Z5g2NtCJD3z80Ud6vli01Hp6yvXrnwtTePONN8qPfvQjNZyuXXuvfPDBL0tHjXO6XUrFhcVlEVNszes8TE3I0RGtS84m7p+B7P1y5tTpMs/vLa/oHvNZUXKyXohHqWRQA0PWWbZG3NzY0jNnzfE2rF2eQeYdySjXPAcaqWHpnXmy4lcMQHceYtJDKpypyXymoGqE1R52RU3kDA3fDgBeuXC4HliR6vou6xuuC1xHg41psou8ahIgfyeW5fyetDPlmlOpn4088i3Wii13TSZU4ybudTZfRPwQqaupScHPvGAxXDUwmpr8qVY02O94mbkvcYX/zjqj0QCJRkXO91CcdbPHNlIGuF3XNtTN1feayEO5blLVoFd4CbGMz6+mTdQk+VqJX/h8ceRQoyisPF0nOHXJahEAPu3iqn5P4HxqVMRzr5wi4nVfmgDFwPFUnLDmyWeJQTToiZ3sH949ZxainuP6M3cGO6vvuWZqKZBhWKMo+bmP+2Vzc1W4HNH2m9/4Rvnxj39S1qjHO4hHLYqLfG7il4hQYbWd+bexpJwxaVt1KSP2DtQkzHuvGIgiLZ4Pz59cE1ySOgHsivwVfBISAufDw3v3tUeZR4MCCNtgWaZDtsK2LaywuBZhgfy9E4XooFxLIPxiYQmO9bpR8feeYr9+g/+/78CloWEFbfkaKjDBbrFXMMGmhyn0+/vaNAII9/fKmgZdG+Dne2wwEjglDnTmI0DxM2pCADIGgKuBwTEXIm2NFAj2aQAMlzPnzqgRcuv2Lf3O8SNHdShRaOIde+XttyW7Wnq2VGbn5g1MtsAE6dQBxP8mDk0o6UESzcF48tRJse5v374t8IqgQqIBY4yDj0YHQYikgj8BDCnkawwmk3yWBG2vzM7M6oycPHRI14bH3dDgUNXd5aDmHqK0+H/Zew/mSNPsOvPCe49CFVC+unxb9gyb4lDkDDUkJUZIWm5otdIf0P4uKVbajRBjVxFaUn44tNPTM+1NdXnvq4CCKfgEsPGcc29mVnUPjTQKkYoGg1NoIJH5fe/3vteecy6FeK7lzJnTlnNAN391VQEF14qRkTRVUuZk8CgY57wI6b/SDGnsKBihuIpzIQAgwSF4k+MVsgkDa8fkAqnps3zxWRXYEbi4+dBqNDioMWLXBedENKvAma9tK2OWVADXYmqtqWkqGKjhQ+Evh2MSIGxT9BuyFjwMmp4eGWGu0YUhhsbRuHGjC4QiaCiCE11TDvxWwM88E6HM12IxBzPyuRQoGETI8zSjxug+Nds0dMuDhKtpxtqBfCeoxymRPJHALywsxtGjh/Vc2TftqBOCQGlZt9G5C9mRuH6tdzPYUpDnIpmAJ82D3fqutPFLV9vFQRd82oOMejaWTGvJKnmYdkubU4GlivkeWl2U/2p0VMBOwGEEvoM+NzsogLvxpFPUptFZ8kAVsLXfSnujwsMWHahWAFTNSSfpDHJFlgQmjdFgFfRI/ze18dkzZlh0iV3TbIIlwqMCegcC1u80yI8C/E6gawm6jsHZi/Pz+pzDBw/qmX/66Wdx+vSZGB2DwbCpxFxoCIq9QgV2yUZobRu7ceXqtfjggw/if/tH/0hoB9ZtbHIi/uCHP4y7d+7ofNG0wP6dOnUyHj18FG+8+aakUAhE2GO//+//o5oVBFb8N+9PMk3jkyBEc20WPQSUdZP0RqKEC7GtInraW53nZAs5MLfMmtCUGVhXUdjNshbDqJoSCayyzWmX+PrzkPN/RUaFZgqJ7mzbwFvXjBXpLnPQc4B2FdX9ET4jDHAksMZmek9Zt7UCaSc6zlpoGPML/VfuZySUkEhI42i/lDqy1VAUmjMT9rKDaqiyBzo6xR60tmxLnsnJhNFbVWgpJKv1u41e1IyKGqLWpLb7/ppJH0g+ZP+EPDJTROw7yQdSUACt68KNC/JOFkGb17Pjs6Ho40/wTaur62JUFKpNCLJEntd5fDkRqvvj6owM+mok8uc1K9qbD+22q66x/W/bmxd/UbzTeq89NSqGRoZ01kqGgP0hmcP+Pvl87H7Jt/EcJJeWX0LXdXXpvCJDImmMTtPasZsbm6CoRsUE5LnvNGhu0MTAToCmdYMRvyXZDNBcNEb6+9W8EEMgqfT4O5ILXs/7P0v2ZjVpK/nBprDeJC7V8G/OXOjsVJGS92BuVtHJKUbMzs5pLgUIY2ZhEZ+BrhobGdFgPdaBz6e4XmeQfSPmhSjzjumqmV2IRB68YwujqLGL5199VUNCKZSxFgOwXjNB0/MVYrWVwNLIdfN2x/su5UTLj/E3xEMUDXlWFPpYQ9iqFJ15HXMl8DsUTbiXuYNzmimA3eK+3fA2ihOZIq3dLkzNCclkDQ+PxuuvntezWl5ciitXLmdDiAGqBiRwbWjZ42vwBS6MbDZlI3xvZlNSyEb66e79+1pjnj0o++ERdIjXxM749OFDndX/kV/EV//4178XD+8/jE8/+0KsCs6Q5Wk8g6MKXlUstEynG7isa832AcBBIZo1plkBK2FyaiqWVVDMGQTJoASGih1jvXq7OuPA1Egc2jcRw10dcfzgAUku3Hv0OKKnN1a3dhT30fTgLI+Pj8bl61dj3+zBeLa8Fitrm7HX0Rn7pqZjeWkxRoeGYjVnvPTDsN7ajvXtNdl+9iMbeksxMXvecwWkRb5LoXkz7j98HOfOnpbkI3uDmXLMDyB2QsqR73mft956M7748qL87KlXTsaHH30cM/sm4+y5M3H5yqW4dft+bG1ZZox5AaApn68jI2kUMfGpGu1ZQNN+Svkgzlzp97Of2H/EztiPyn+4L4ruPKdq2jtms42j+GGfGs3BxJwbCsfcu2KEHuav5LwlmB7JfKlYib/1LCbHGnzPe8AWEthsxzrXkxPjAm1QvKEx4GavGU7YxEGkLKQH3iugkW2WZYFsW/md2fk8E64LtgAMRTW7iF9yrhS2RLlKb6+KTtgPSbYk8hskP+/PGbV074CKNVWYpTDPOR8ZHY7TJ09pxgZzrdiTI0M0GZ7HyRPHZCuxIfhK5mo4VLLlcqPG0lvYHs5A5UM1O43ngk8GFEXhnGviegEWnD59Oq5evSa/j62WRn5vr84Ja3H//j01wAroUAPC1ZTd3FSeDWOMNYQRRKwYXWZ+U3xCbpmmCufY+3gxevt7Y3BgSMUv9jXn0jml5yfpvHf3xMjYqJu/m1tqxvBF/KPXMl8mZ8Op6IxEc9uQ2ELoq/DJMG6KsLkP1ATYDdlAIbWZ7TUy3Pye96HQzt8S9xqUQVOemYApeaK97sY+TRjWHEWCkgEm3mbvqamWsW2xKrDjjmc8l6OAXLUGLSaq6xQClpAfJeYF6ac0e2JLkQxwP7sdEQyxPn74YAz2dUsVATY0zxH52MuXLuksnj9/Lq5cvhxHDh+W9NOHH3wQT588ibmDB6OjuyuuXr8qabbjR4/G+++/r8LrL/2t78S7P/6J9gdMJRoVML2CgqqCrjzvm5sxMTaufB97jV2Q3+rpkbw2jLPnYm17Zh7nVzOWZB86FK9o7gnNiKzD6N4SNc7ncLZpWlR+4MK+ZWuqRmBVBVgbBnSYGWMlAH7O2S7JXwEis5mCbXbs66G/9Xc8OwMnnDVXo6JqF46rk8kDYKDm2SQzu+RsFW20DQb3njDwgbiu7CTnqR9ZoNx/7cXzmlXBnlD8moBR5RLNfNJAQwP98vlksd+RvNfaNZZkLAP0LUlkYq0EPxjMa1tXz1rPqk2q2bF3a5afmx7et+0xesUYlbu15yR6j5/RqMAeu27nho7rP645ZKLUjP2rHtiKZ1rKGoqL9hLUkc0lrVHmaaq1ZD2rmueJNvva8Ki9QVXAI2ww0s0Vi6r5uEPDYU3nj/qLFEY6DEbFvjV2aQoBLGKWZ9a+dmA8s8+3BGY7deJ4TE1Ox5XLV2MJ1umWayFcv+Z9ZjxUCjCsAzYX3zM4RGPZjDFqhPUsDQzt0bBr8np+x4oCOLtz547AzLMHD+b5nZdKw+EjhwRog+3L/F/s1sy+fbG4sqQZadg2gE8lQU59QiyLvE5ej6/CDwK6RLJRtu8bRsX/yBD8m8/+77ECJ/odkNkugz5Dm81BtAuEHoxdB3ITyZEsbNdAMMnXQH/SLAVLcPDVLJDn7AQNVU0UJJ8lmmlqZ+KAKA6NT4zFbieazc80XJHh2hxiglQxMTTk1PMCYDsQDGKYNtehT3fpdwxRIzDidyQtBKBouoleiEPq2BOjAs1SEHcYbw47hTF1RdMBkXyC3pO0kry8EamgIIWU6rVmPIG9BlsuLQp1TUBD0eIIAxh3dhRE4hAoRkDfUnMi11eI90RwS7amwXAiB2cK2tT4MYWw0C8EtmIMSGbIlHLWvTkkSsPZUvc5dQP5e4oDpRnfTlWrol0VCatYXdV1+6EsdiY6pV16CANekj9QabkmFUg1uC+HEmUhopxWofv2QFzqvnfyWeL4TfnkM0Ci0bQwwmlXMy2eLRlJIrQPckyQyaUb68ChdMNVKMmhW2I9ZIDF9e7bN6PhnCQE7BnWjqIJCS5F5Cr8NvUym2FKuvOSyUp4hAsm1k/U4F4VBayn2woq2r7PQbiVQNZ6NiW0MigyOt7nk71QBV8xDLoIfLZMs8xBaBUAVVBVmvjNJgiJdDYMRKNN9IeCl6IGJ3TJ+9ID9ppoivxZ3YmkxqpBkywKJwVGbatYmsh1zg7zSIwwMZKpApuSCBKKIZNrL22uYw6NrkZQC5XSQngSEHZIOqBbTIqZ6Wk1EyhGULREfmVocCT2z6Jn7bPM/tjYdOIE0lJ7l4atKPV98Xu/9/tqfCIfhyQPQdPa5nr84Ad/kAwoSzARmLCXSECgaM/OzqoxcvnKlfjphx/FJjr3KXukNc0CH8kuiS+JtwcNUvBwYRT7aQRH2VMXCqoYn0Y5kRwubhiN578tm97uN3RG2ux9JX/tDYy/qp+p62vWtvP9KQJ7jd3AVUMhZYzccPOZsfSEaf0Zs9vWM4sjYFSs6pKKRtwsercV09UMwfbkoD3OxvDoiFhtavxB1SXpwZ8h45AzBYwYknczu0Koz201kzgnmjkgNohR+XypMZRyerXW9TNeB3IR1h2MCp8dJzOwfHQfkho0M03PQg0KD/zmuiYnpzRbQ7KJ2MIc1G1taaO/hTzKRNCIRheHQOpSzOD/XWixtnRde/veqPVvbzLUnvkZPanm+7y8R/68RsVfdT+1v769UYH/nZwaF0KQ5Js1p5HpAmyPGhUkzthJZIYsywJ7wRsFHwNi07IQ6U9S2kdDWPU7mEyOe0BKgezGB3mo5J4KMcRHkpfcI55xQc3NMRC8W4nA8z7hZ/gEUFRiLHZZDlMFxQgVmXgdbJCivrs5CVLUDS/emwKf7axnsYyPTwhtBfihpD+wFfjK1XXPrFLRIBvuasJ1GNEshLPWz1IZKlxnMu29aoo768p1IGUnSZ2HD1XsUzO82dBiuKB9RO0nodEk7abet4d485m9vTrLFEdsuyLWniNL1SkNYO6NGEnxYzZTkItkrQGRWBoSxBto+f1x7dq1aOzuya5zbscnRoXFLUnBAAAgAElEQVScv3TxUqI6KeQhF7Cu90RCA+YRdoQCEUUeniX7iT1TCE8VBhKQUMPoaTqvrT4X0pSCE+uH9AfPcml5MQYH+2OzqyuuPH7y37Ld/5v/9lfffDOO7p+JS5euxOVLVxR/KabE5mlOEM0IF4u4dx4C64vfcrzfAklsbW/anmzQNDUqFF31AhWBoKbIrXMFU6YzYmJ0NKbHR+Lejauxf3w0BrsiZsZHtX8fzS9G3+hQrG3uiJHDwHrO9Jlzp+Px0ycxvX827j2aj+3djliX5vJwbAPSef5cc6RoAlHkZBDtzCwM2j4NN2evHJqblf3kvtijJO7MhQKURFF5fXXdAKbnq3qPt956Ky588bnOJyw0UM74eOJWENNnz50VAvnmzRvxK3/7b2nv3b9/P27euhc9Yq/BSOhTh05jcMuWiw2ZGvjENxTOQPMSF+ZZ7MUX5twK2MFim6YNozFkn+CtYBlPf+9n45jFjX3L87L3rb/erYZhoW/Fksp8pmn/U+YW+8Dz02yrPSNDyZc2KdgDotq0jOCxI0fiyePHzfltvBiwCWeFps33fv27cfX6TTd7NmEggSz1EG81uATycnwvuQzFKAzdFb5ENlF7UPPKfH+WEKFgbhvPf5ODDQ2PqEklubxN5PJWlOfIlEh6dUezYw4fnIvNjVXJgkmKbHtbdkGyfEJUd8XQ4LCZIpn3Mo9EbFVk4bK5zRmnYU0juIqF5HU0J6b2TYtlQ6MZ23306LFsHrXsPo1XmI3YeMW3yKh1dPq6czakCsar9gfYJQpw5KwMe9dAaBrLEXHxwkXllvNI29L0Snks1oOfgTbfyUGw3itmYFLsw5YJlZzSNS15Fb+uGjIGQRAXJ2iIZ5NMROXtDMvW2jBA3jkodp6B2ABtyKPI4SUbtNMwSJF4XGCLLbESy65yT0bfWy7GKHdmNdSsI4O2iuVVcw6qSFdF0AL0uNDoBjSgND3blJsqwFbFKBRYrY6wTS/I+45B5Y2dmNk/q5gx9hoxMzURp08cU53iypVret358+c1SJvPYV7FZ59+ohgdQCKNOIqS7MHHTx+rdsDMG/KP93/6vhDhb731dvz0/Q/kh3p6+mN+8Vk8fPTYxLSMKZ1G7YrJ4bmUzufVsBiwxCdgFObksPG5PkAJBZyxXI+LyqyxlS2cC+usvABC8X9UriY/wTnN1xILlLQmryt5GeIu9q4Ko5mfquGY711xm5oJacO8h8zkqwupZmTtWdm8WgfqJClVVNdd9SKedckSFbiyGKEGGDomE6BLqgsuRPM7yVClnLPirPxd7UfsUzHRDLRhWzqeKlvsBkGCM3K+gfZgKmMoHsx5gMU6UTyUzMbKxytGb+azWU9SPsN1p5ysmkMmd2T+5qZJM5BKtrTBLvWcvwZt1Iww/Le+D4MUig1TD5F9gH35ahPD917ycvrbbI4UeKyYMyVzLv/Txtx/OdDh9/V8ahYr56UPphYA1ZyFyr/EIthUbAONZ4Cw7HGxDncAunTFyspaDA/R+KW2sxWDg/glAxpOHDsSc7Nz8eEHH8X2bsQG8nP4zmbtLxtuxA89Bi9iP8kJ8fXMJSO/oNmwuLQcJ44fs4R9RNy+fUfnRzLRyd55/PCJ5g6q2Zqy49yvYvXVVc/Z6+9PexkCAd24dVONaWIg9gKv8xnpiuWlFbOLct+6lkd82yvf+E2j4uXd9c1//41fgUNdDkoJlEsioKQSROMlsSQ4qcJSV6cOkg5NFj0xcCWLY+qcmx7thZJC6tngcqj6zCzIQjNOmJ+hL48+PIkBh5MOI8k1RQgaIRQKQOARDN25e8eOYQtU44AMhWczWMew5HpAAqJPD9IFY8ag7I2tdQ2i5N4xBhiVCigZskcQdujw4VhYfKbrAOkn1NTWVoyNjOq9l54t6R5BaN3XsO+GUNkYpM01SxFobdOhCJ2SRUqSZ2mxJtpZhl4DweTC0okYQUy2r3kTFPNwZOqCm5Kv7jGUZVATaN1mwVmSIckUqeBwYMjySkY15Hsk04EPVDGubS6Fivup1Ygh5Nm4CZWFVskfuehRqApcY3fOSWjuiY6OZoOG4N0U5A2jKdA57G4NdBJFU7MgnKRpnzGcNGVwOrq6Y3l1Tckn+5TnoIA00SZcJ2ijQoUQLHtQHEVyS0IhPwUCp1AfJLYkr5NTk0KmKClv40BUwFNNCzn4nJGg4COln+SIm1Gg1+7lGR/NSC4p/PbfLg41k4QcoGXEg2nV9aVkozlUjqTVxaZWYOhr8x4pdHlL7obEkf3SkvpwwOOA5cXApgKjdiNnvVEnnUX35L6NRrMMgdYkIzolB21vQBBVTbJqaHqzt+i89XIX810AbDZa2miyFUB5b1ozVQWr0dF44/XX1OxkKN0br72uAXSgHY4dP67gy1qnSOJQVOjWWeV8OZG17fjww48lfXDq1GlR90EoMWjv2s3rKmxI41uF6T4lhBStaFbw/bmzZ3UbP3r33ZhfXFRhxjauv9mIqIC5GUBnI6OSBBckTI/XwMEMqllTyWHl86oAXWe6HUlTQ82yMdpMDnP/uhmajY02VMwLjYwKh8WmM5rKlO/W51cQ+oIzVNHfhbAa1NhqTrV0Xjm7kiqQpq2bBprR00DCx5IOIAqrkdUaKp37PK9b+1fyNbYlXCdFhKcL81qTaj7BhKsERzYik2TeRraHobo5c4A9jl3ApraSPDdWKsEvu9le9O/t6RYrAhkSXUsm0ZY/c9OG75sFUZoPqQXLs0TekAYJzfZq3FXhoVgzFD2alPWUA+L90DBeXFxW0Cv2SVvjqtalmirVLGpvXlTy0kqCWme5/Vz/9wp8Xm6atH8mR38fevagkROdWYUOfmYZFJiKDMCzvnPNeqkh9ayH2XGricgz6xO/TrGZv2HdKSSB8ESH3bR+J74UIdgrDHOWf9uxlABJBUAH2HhOKGybYVqwj9AaV8Ks5M9+iPcr6SfADOWzjLxzE54YrEAOKvgnCECI8Z2Gh88mStKx1Y7kzjQIuRDJKf/mhr73MjbLjBBk9lqSA3r/mlGRGvt87tzcnBIzmD5Ce/cYiKA9laxHSYQQC6JTDFMoi+Mgei3vafYnDV+eEY3I1edrTRYDhVLJo4glB0CmYdmH3R0VRxVrHZwTs4U1lWTL4LD8jvzRzraaN8RK+r0Gne8JrYxcEw0GCjqzB2YVI/zk/Q8tVZTDPpsxw8ZGc5gsdpa9w7WxniUHVU1N/CgoO5odNFWe7e7GvZ/DYO3/mvN17tjR+Pbp09q3ly5djsuXr2rNC7hRtop/+ZmBO26EVpxFIq7CjRq2W/HWW2/ExUtfxvr6puJTnjkzH06dPhO3bt6MN954Xc+PgdYUDBgwPj40ED/+4x/G9spSHDt4INYWn8Urr5yI1a2tmF9ZjUVYHl09QqBvrG7G2bOvqEDe1dsfN+88jMVVy/OQ7N+9fSvWYAv19MT+AweEPkbfeWpmMsYnJ+L2rVtSnqKRNHdgVnsCVDMgI87soyeP1dSi0AAYANbj7Vu3hYI/sP9AvP/Bh/H2W2/Fwwf3xb547fz5+ODDD1QQxO9/8slHcf7VM0JkogN9+cr1WHmOhEqXZuUpZ5I0FkAmkN2egSNkb0q1mpXjpmrFTNV8Bt2v4lk2o6shXs3zstWcg5oBwWsE3JLdT+10xT5uhggslrIkYD5owBqEQ6xMUwRQEEUSWBQ9mukmiSDylYal1tQo6OqK2f0HBKR4cP9ePH78VHNBQHuqMMPgehj32MfYEzirgDGS3+uxTTY4qmaxgbq1fy//J3BYxosulBoYUHkLxWszblPCh1xtfEJ2lNwMKTp/BraDptUBzTJiCDt7mJiUhhuzygAnHTp4OPYfmJV8MA1fcjGaEdgmfDaIeArv2KeSi7UUpJHtFLL5l0I0jC/lmx1mZeHrYTrQwJYM4SCMChC9g9ojxB7EFPwNTTPOxZPHT9TIJv9kvQ4fOqwmyFaDeTIwRUbjk48+0Z59trikdWd/3rh507KFm2ahab2zYE1OVk0K3rNd6YA1bqLmm9KyLfBMs7CfsTd5pfbG1oaAgtQ1yyZWnEbeS+7EGat4ib3J89AswmZh176xCtSFJneh1owNI/NbhVTHfva/5WOq/gD4A1vPOrBfOCMCLGomg5kWZqZ6j6iI2wmBoTMamj2lkN9nZy/i/Kuvx+r6ety7eytiZzsOTE/GmVOntdbsSeSeLl28KJv5xhuv6bmQc7xy8hXl24CTyAEuXPpS+2v2wH49zz/70z+VL3/11dfFdON6hoZHNQuRz6f5yT1zLvFhPDP2pIZq95Cz0VT0OWKfYOMAUbhhaKm4ArEJRJPnX8OA0dTPvIy1qbycc1FKDmp+wWohN9J6mqVd+4a1FyCxo1PX5ByhBdDgeRDHw1I0sDKfcRt7C79cfyNf1DYr4yv+rvl5tm+VINbeVQ0iZwfUe5q96qHIZU8U/2aDvoBp9n/b2djO+XA150r5k5sCVUdqByFVc6IaGdVgqIbGi/GrC/qVh5dNd1xq9rv3ays/10zBfH6co6p91MwcAxqrvtZqxtXnY88F6Mjrr/rEC/l4NvEq5xcINfOg9gYTf+M41Cy++qq/Y50lL0jtMEFnlQc1X5u1gGKYYBHKrlctQ/YgFV1qrVmfalRQn2GvsO+ZH8T3NAW5PgAQau6mZKLqh9moGB+bVNOSRsXIMA3WRuxub8W3v/12nDl5Kv7wD/84GrudsZnzOasJpRoYs1M3PetG9R01t4di5flSTE1PqCHL2UJlRfPLVlfNqmaOSuYm3KeZk56zwSJKSjRZwwJXKbbpNftidU1Nx8bebly+5sYo+QzvN7NvRrE3QHLsfTN/6aImCJt1O+0u8ciBd9prLv81seQ3f/PNCvy1WoGJdQ9ilKFKOp3pYd1Cqr352uvSMgZNB9JDRfQu09XK8FOwq8GuTUNXVLJEdYpyTkFmh4IbDA2jR6qxoCLf0JAGUYGKpMjI7y210G85pefPFfgx2PbO3btJ8R8SUpVElmsi8AQJNjM9o0Iiww8ZLkrgLGmMA7MaZvPkKQggO/GakbFvetrBKvMPOjoUdKCXyu9haUjft8MSURQKGPRDgkQDpH9gUJISK6sgtlZjR51cIyFciE50Ss6hgClCUKehZDkEmQbQC8XiZiESei7IzBp6RWU6RGlEf1nIRwYE9yOPtKnEnfvivfgbAiTuAVSxdF1rQFJS86xZbMSymRFukKgAvOO5GewJkhN+VpJVctqaEwGLYEdyWBQDoF1Xk0Som5QtwdDL+ecJkCZ07CogLwQBr1USLTS+iyHl/Lg+aOaLoji7kMP+KIdH4wunyvNQIELhlkJoNlhYH+2RiXE/G6Fa91LGI9SogHbtQVxff0ybBMnmQC0XoJuO/KUZE1/XqGgPXl5uEthBQpNmoKmL/txfs9AmNBXBiOWRan0KYVcsKJw4fy8EfiaeNa+ikgbfYdE5Xxysrl9VsiDUWwalOeScv2silYWSd6Jj1Dcso6TPti2jBqlLv5kGjNGA2u8vBUF1Xb46S4fUOraCJX+3sb6p88weZI8jfcNbPpufVzBx/vzZmJqcjNu3b6vYdPLUacubdXY62Q+Q+zCNqllW2t0d8S/++b+IEydeieMnTjRRPhRLfvLBB/Hll1/qORCAIFHBfqRQtX/G82iOHz8uNKZQvyQNObTWQ8/97NiDdT6EfK1B6WkvapaDNHyFFiGItbydBsvnmjejYS2YF7PwNu3NtUoO1UwiWE7kjYruubDt9qeC21rzakhUo6JYBU00Tb5QRydlFVjrdqSO5ZVsA0r+yzIXRuxp3wqx7WBUzLmlxaZ8TUnmyCbk/VcBfi/1VPl83kMSWyC02ceSZLYEoZleTghqaLSuExuWxVaa4TwbkCs+Cm5+6CymBJuTg9SQbUusGbLLZ0tepI0RhSaxz4jtqIoyKpIa4V9JCMVr5O0Isklkmg2ivDajCHfMDsw1l4Thzo5mneBXuEY9byUApVXeQkvWs/PvrcntBnRRz1uMnGbS97OM4s8ponm5QVbr7rdH4hE5tUmjdtVkMiuCddQwvUyqoIbX/YmSrUGsngnDGi8ursTRI4eV4IOGlQ/Zaej8sh9Awfb3UdQLoe7xd9WsgFlALEHBy8kVMlCr0h3H9z16/EjPDBtOUkJyxfURS/l4uslYhSKeNc+AhKuaCCWZyT1Uc4L9xBexBee/GEqa29TnIbMuVnVLz51kRijjlEErgIEQ2TnPAhtC3OXEMdk9qUtde6Kk2k6+clIxGetFglaoba6FArUAHwyQf7YgGyRZF3wFxQuG7SIVI4k9M+14A84BDDt0wpHzBHgB4IR7PnX2nBoeT+efiP4/MT4WSwuLYr9RNMeXE1P29Q/GU3TthexkVgYMi2e51jTsDVwRahy/HhFHjhyJ3/rN34h//i/+TyFSy1ZKqzzRl5Wkl3SYG/+2TzV7jWepAYt9fZILQgKFvXH3+Wo8yZlkP6ej8Re+zcGpyfi1t97SfoVBcenSpbh185YaUsS0xHUugjhm4EzAsJGcDgMhd3P+zt6O4mdsy9DwoPzpo8f3FTtqBsN2QzHviVdOarbX3Oysro05I8iMYc/6uzriJ3/6x7Hw4F4cn9sfw/1mPX9y4cvY7e6Jk+dejYXFpXj6ZD6ePnkWb791Xrr7w2MTcf3Og7j78KnOyeuvvx53bt+M50vLMTmBvM6ZuHDxkmKh/qH+ODB3IJ6BMN/1LLPpyal4+OCh9ifFbWaj3X/AcPuu2D+zL65cvR7Hj3LutwQs+rVf+Y4Q0OwJipHv/eQnihlgynz55UXlH4cPzcbCAs2OfSoaXL16PW7ffahi+6bQ/j6jNHjY7yUdhm9nnZDDkr8Ps6O5du5NwAgBENpZdhQcUhqkUMV4QgExzNpwAd8DkOWTkpGITeQzq6GHn5MfBAyVMwfKFgAkwpSDKC8tbedkbAOal5YipAHEGWTN8CvIYjGUtB8ZW+wiw0SRHFQs2gIAVEBn6QzvKzNhdxUnbedcG88T62rGVpqPKGg5/tuFdq5ZCP29HYG/RsfNQKt8hxuRhG9XR0xNjqtYQzuor6dLzFbiADEgJsbj+rWr+jyGJQ+PgLZlGDh5KU0WGtWDavTDnFG+1NGhofK8jmeHjQb8IMZbY1v5V0lvkHMAptPsoK1NNbko8PO88Q/sT+wDZ5GmNHuGa1dDHWmkdUuzYV/xZTwXoYc3NwTM41qYoUJh8MsLFz3LMEEZsqWaV2EAGn+PX+G+uWaBNHLfyf8wf0KMHPt4sfQSiFgMUPliXZ9zdLn+DgYab8oulM0UMC33Io0U2B18ruTjllc0Lw6/XfG1ADZZZ7BRawX/lYcaXtEMSJuvqAG9VQyW9FN+ttQcEhTDWvP5rKXnLnq/lzwL+SCMCs226UGaDIWG0LzLM2dfjUOHDsX1a1fi+uXLMT0xEm++8UZcV1OoEefPndcwbS6KeRUfffSR4tBzZ8/Ehx98qAbWb/zmb2quDY1cagqsB40Fnt0br78Zf/pn78a+/QdiDVbE6moMjTAL0cx4S5xt6HwNDw2IzYmt5j2oR7CXeMbstbWUeHZY5uaoGLfJWpYc25bllM2iLBCZZX9q/gDrSZOxCrS8rubMcIYlp4kPQaMff6K96njR+8c1AzEOwrPAqvlYckouytMVaj1aZJkLlNkspDtIsv1JBDnXUEBDg55sS6qZKVuWP68GScXlXItzYmIjA77UVBRQNBvNeUmK1TN/d+PHMUz9vXOFVvNB954sDbfXMvdqz2dbFJOMSRwDkgd6vc0ILjksA+jMNq/mnBsyblBU7UD3DqCgtMuaZ8nsNS1j1ii8tj5TfOt8oz13KTvgZt7LuX3lOW1HMgGyADpgqLYGeEuqDcAZ9/0Sg6IUBQqY18wFE0hnaaOtZu0GGwajgnyaZ8D+X1h4JuknlEmwoYAPeS40UMVk7Esfstcl1hExyujwYGxuPo/OQF5+OF49d07n8sMPPo7H84sxPIZEs1lYshOZi3umUJdyOJr6Y6PjMTI6JEYF/kGNO+TMqXnsUCe0DyUeZh10L41GbKxtxuT0lHwZ8ZZy723kCvvke8w4pi9quwxT6sLFLz2DTVJX6/KzntdqoGfNSOV3fFXuqGb9N42KvzBe/uYFf8NW4EQOMCTRxQiqAEryiQxKIosf3H+gAI1gjSCsl4IvCPUNIxFfKK434wtbawUdUFr7BxR02QyaZsZB5QsdTpwzwTaJPT+/fv2qjA9dVYJgFf8bOzlwu1+OmiC/NNuq248Bp2O5tPhMztLahFD+ezTkikRA+rqbaJF67sbQwGCiIWZkBChgIBVFsvPo0SMjLpN1AnKSJIAkBAM9/+yZUBYY4bt37+rf23fuCsEn/cJMXpQ05NBP7rlQuQrMWaLU/6xaUGtNvWI4zZrTUNJbODAcBQUt7hNjljgHrQsIC9YWQ2jksoePqeiTCJP6nGYzIIe/lt9jfSw14vBRRebUpLXjS3p5IqCkLZvfY4z1nEGN7e5oDykAzxkllqzai8ZeI5Hsbk7oHrIh4kTGwSZrsL65EStrG3IsoiyCsunpltZ4DeTCmQmF0URs7DUlxlg7AlE+m+JVoVdo5oBwoshnmu3XdCraWAcq7raxJ5osGDlohTPNwMRHotUQcBBhuYyMy5oRSFFaq8DLs6qikdD4agoaMaLETgN1W0VFF0+cmNR7FwOjZmG00BXN0MP17bYA6ytmLJsKkuhJGRzLd3mWiopRYkRlkPQ1dtD7x8l4oTgVGGotPMOi9l1dCgjhQrE011uBqdkGlViRADO4VhrBT5+qsAUlk2qjdFQTdU5xi0BARZscloVNA6kg+QECE5qTYl10xpkzZ/SeoHsPHNgv6Y///IP/0pQPgs4O4pDX8joGTJIksdcZtk0iosBbTSNL/Bjh39WkVJfMmGxBfRE0ZYFCklY5kLIkxgp50wpCXTB3IOugubZne4Bb+6mWupp5Ldp5awhc8wRkAC97nsWR+tc5Ur6y/QOFbDI7ooLqYuU5sW09bzcBfP3FduA6Ccz4b4JRNyQtHWBEmM8QAbcDtc6gUaHLAR3aDcJ3WBJ/RugR7Hv4q5CNQuA5SWhqOjeZCfYznEH2Tj0X9j773cyLDIjbBmwX6wLUKQUOUJLes26CVSG6qOpmkEjdudmM5XWtRgW+i0DZxQS+NCgwh3YXg0sN5myATU1aQ561wj+JaZRNGDWBUnKoWZhI6ZCSwKq9Uxkl//3fo1FRxYaXzcTP+rkauns0k8eVfDQZbbn1JC+y7UJsq+Fin1vSV9gIyckgUTE2JmkQ+dR8psr5Oq3/joY5RXWYECoK7allKoQ/z5aCvLWQLcGC1AzPCv9Rdpc9W3NVjCz2AFP2SRWPsBOsbyF3uTYPcLaUJTZFiXVKjvA96H3iM+wWCDNkk5DBpFHC/cECrUJbMZ/qnPD37Af8sBswNLzaaf8ubmrd8Pt5tg8dPKh9D2DFRTJsmNF7sk3S7CUhhNVpaSgNTe12MYlmgxpMAB50jhoCWSj+Gho26KDfiEjit7X1zdhQ0rol0IcKvlsbwf6emp6UVMfFS5djdQ0Em2MOmhJc572798wAznsDyY78hGVVXLz5/ve/H59/fiGu37iR/hJmib1OPZ+yJRo8LIkeFwJLmquKH/gh/hTbTwHswOz+uHDvQSxkEvk1rvDn+qPJwYF4++SJGBxkwDqJcIc01e/fM0sA34YZwkcTLzpmppnUo0JYV1dK7CR7FpnEXhL+nUacPPVK7O5sqRE3OjoSU1MzMTo2pqKXZYgasZssWAAqDMce6u+Nd//oD+LZw4dx+MBMTI4OxcKzxVhYWom1xm70j4zGyuqaE3Tmf7xyPB7evx/D4xNx697jWFh+Hp3dvfKhYtNsbcT66moMaH37hdqFEc29rK6s6jxoqGyXhwWrINLdIwQ68dLDh4/i4OycpFk5X0ixMPMOO8JnwNKg0QIy8uLFSwIi0RC9+OXFOHnyeBw5MhePHz3UeaSxdufeo5hfWBKrYpNGWEo6qAEEozmLt5rF1fTnlm2pIh7vRTMaPX4X5KyPTW5Rch8V4ylWoCmbvqoYijXHQjKy254twv2Utja2a2XVMhGaQ4HEULclcgQ2UC7gKxSgip/toeneF7vbzs8EGOrslJQhA8ovX70qJDdzJJCzxC4WYK3loxyfak4D4CmGLGfMKvS65qRY7srzxlpBD89Sc866OnU/gMH4nmIrRSPNqWs0YnwimXU5x4ffjw4PifXN7IGNdRjXzgHYW/umpsQIgxXw7V/8Re3fJ/PIhgxrH3d39SqnFOsVtpkQri64U2DGDlP0x6ezvuTA5ICAEdjHtqcwukDh2h/w97InGYOyT7DRYvo8eqQZBMQi7EMYP9hW5LbcsPHAct5TLP7x8WSK98SNGzfFrKi8wHEfklmdMT0zozPJ+7FnShKsVWwEIGH/42aEYwvleQJ2VTzVIbYgjVeer4eK9wu4x59VPkkjVw3oPYbbD+t+aWawVpIyFPvUrHj5RZyNVJTJJ5tZUmVLjtU01vqlr2QSqjlGA6wtry7AThMElPJhGqQrQA75STZnhP72IHn2f1+v2ftcJD6F2TgnT56Mw4fm4tH9O7G08DQOHTwUt+/e1QWdPXtOTWBu56033oyfvPee9ucbaqrekawXCgvMOqRmwH8Tt1AbYB1fe/X1+MM/+pM4MDcXa+suZJKvbksqzeCVAtlNTBjEYGUIA/OIP1gD5mZwnh1XugFRzYOyFxWvuinlwfN1Lr2/QHD3tgqtW8yNZBA62v/riqNlS7JeIRlLfHueW86W9kzlBzQl009WvOHrQnbSdqReW/EnwYeL563cR88+4yR8Nw2FVj7oVLnk8kpisphkJWNd+YTeu+az5bVjX8n75b/IJXKrKQ/Js1S2VrF2DrhuxVC6wCawUz+vJCvfq5094R+1dnSdNfN+ZIEAACAASURBVPZD7V3/eav91/5zSUAlc+7l1zXZEJlHVxzv98rc2qiSvIyvJvn1ucJz6Rm15vG5eF9Njfa34X2cUwkwlNKFauzUrMQE5ij/TeCymkxZiyp/IQZiW9NUNbMtSz8OJFOC+8LO4udpxLpJ5eYT8Trvj63WbFddLzKInQLwdHWietAZja21mBwfjV/81ttifn722YV4vLAUA8NjVoNQruCGH/cg5gJNAlRScug89YiR4UHPsQRsqLjTEufYP8fUltmsRu/S8vPm0He2AX619jt+W/NlGrbVqrkODsbtu3fkP6lVuobo9SAXLoCRwE7NOW2thvM3jYqfa3j9zZv9dVgBhmmD8MAgKVhNdL2Rnq0Oc9ELRbFKhIn9SUsGqP1+ZPwScS+UfmeXBkILRZPSQAoCGWKloqsH0NgxEDCZcg+NEgcux5kFrdGR8Xi2MC/2grQSO0CUwDZw0I+BoSlB4GcEGe/fKRQN9KojRw8reOcaSawYtkhgRZeV+6S4CEMC4wM6UZrUqTvLv6PDI0IcEEAcOXpUXdKbt2+lZniX6Oam7CFjhJN5kdpcBcVqQHCNJfPx1T3hgjbOVQPLEwnB64aGGBrcoyHjJG2gIqRbzpCrrc0YGRpWV1b6y+mriupJUOcvv7cCijY5l3KsCupSIqWYMMVEMEqFrnMGIzAnNINkVwPrNGCRgjDaxoNIVbhZgU7gIFRo6OA0KnaMtCR4ZL1U3MGZ5awNnjsJOIkerJPFFZKvreawahUNswjHaxefLTWLLJIZQpM05aSGhikkDzURxziNhYV5Fa7QrVZzQzTjl8KLl9ABmiXRRL15HSseMWLIwYmdZgYqTfKAHXerYZDI6LaioJIQNbEqcXCyar1Ssy1w+jSpWC8CWV5azZp6Vi+eyRcDpvpdq77cKlK3egZJx5bkmNHXXHcFJhoYK61rF985Cx4A99WdrCRk1006N1JaBfVaixdXnd+39DaV1rgy3izC8uxhVfDv2bNnjDj78qKGn5JkMdSeQYZ8nmQJUjJEslwg5rl+EoBEhmggVzb0zp45E8eOHVdgYXRNV3z40YeyK9U0G+gDAUzxckQNMJJTmq23b92Jz774NPqhdJOpaECcC+1mKFkvlYXSKuT+cmHY9GPtLzXbHDgWat4oHBegzXRpIXv890YNuYBQ8k5OTF1ML8q2E4cqrPBG1UBqf4B+Sg5YpT+f7DC9X8pB+frag3GF8k3UXxVP1EAlScwEpwJY+5Ia5GxkP+eUL4LNYpOpKJPSgzU3gNco2S5GRaK3KK7BqNDaavC8Z3hYk98asLr+bEB6lobPGTRe/k4FZqGR3fiTnWy75/bvtYfTDtFgfzoPos9D+Op1xWoq2+EiFX/mZhS/Z/+QREqqLs9SFYMUBOcaKBXJORWo+WIzJyYn5Js4h2KkSRbPVH7Lizh5r/cr9FShxlo2Kb3DX7JR0WravnjuXzzXrd/97IbEV+1GXon01ykgytcl4pUCeella+YVM52wRdKbNavM7CNrOZPIuBGArIblSzRwstsoZeKEtfUN2VjQxAvzaG8jrZFyZIODOu9lvyQ5wYyrZGwqjlITy8hGNwZ7NHtBiLw8g8UExG7wRaOiEtjS2+V68Jc8N2I0J7bs4101s7hvGKMwxfhb/g77t7wCo6YkMWwn2n1NybM4niI+cQOszrikn9L/cGbw4chlsqdBGyNr1oe0CyzPHN5JURCEPIM9aeRw3rhWBgPKB+acI1C2FLbZnzCP3nj9De35Tz771LImQmQimTJkGShsQsp5/vI739bQWvb00MiI5jAwmJR4AFtDLjw+Nh7PFheMrlUB3QwqTDDXRgGPa33rF96OQ4ePxL/9t/+2ycaj6Eb854ammYg+0kbLi9G5bTkWsaESiVyDibX+emaej3J/bT0erzz/WRv65/Lz/aMjsa+/N8bGJtTEkf8Ccft8TWwBCqK2F4VydFNYfnyXvZpJeE+PCrQg01kzWIoUdcfHRmKw3xI+Z86cjampfU37CwiGOFzId8WOdvCjQ4Px7p/8Uczfvx9zM1PR14Xv24nVre1YWFmN7kEaUz4j58+ejds3bliuo7M71rf3Ynl9I7Yau2Zw73h+GIOSabposxJXdRhp2J8IX0m/JktNUkopL+v5cQyVXxciUzKujYYGod+8fkNzD2BbIOV45vQp7UvY2m++/lrcu3s/1teX41e+806srS6bkbPXEYtLq3H52i3FuGvJ3qi4wr7YRSKAE5wR9glxgWR6NjYEggIBv7S47GHzyWQrH1M2ulhuX4kDdGYdP6oZrXNCsd2z9tivvAdsTyTakGrB9vE5YgDRiOzsVvNCfiD3sgZId3VEb3+P577Q7IPtmKAKpK6u37yjQegM6e4r+TlYUyUHWkOLc9AxcbXmCenMWxpqM2XHHO8TyyK7yfUMKA4XQjsDUIoz3MPjJ4/VFMEesu+w6WqSZQGW/UMzk/OLPcT687OpyYl4whwT9PTZBxtr8c4vvRMTk2Nx8eLFmNrHmdmO7k6/J8+KPJQ1w5fQtLW2fijWxi/LBu/tadYZ+4mGN2sHOwJmLw0Gz39pycdQWFYTfAVVgEGdyZr3Q6OCZ4KN52fIHfMZj8TU9++wwexjaqJ379yNJ0/nE7xg1jznSdK+ypU9U0axg4YLwxgwQ6J8gfJwseGZ4dTSqG8C53K4sIttNKANJOTZb24SEzln5NrMAEATfki+lbyYvNmNn0TNZyFXsWMCcAS0SLmngnY5Gv2a5KGZLWSgmNbT4I8EpWV8z57SPJBACsrPynM3kXqFgdivvHN4cEAzKtz46IrVjS3NxuG575uaiMOHDkQn+6rRiDv37skeMUz7i8+/0Pl788034uOPPhETkMHan3/2udYUebmF+afapwzlZo4O/p0aw5nTZ+PzL74Ui42G3aMnTzWjQgxROjh7jlWliT8yqhiFtWZfqTGObDI+bBdww1pT/qjAYwVEkaysZgLSfDAgtNjDBRQS0y7nkVAU5RkbTOnFJXZy48TAHM2Iy6J9UirlVwx20CAHzaSq2LKYkzRWlD8lTIvfV+6g2kLGmHUPTceYdSHiWlhbxAuC9bSx9c3kcD5TbIP2/EeFdwByKW+IvVAukZKXL7PBDYDxfVZsXAX8ev/KVQwGqzy+siRffTPn/3O8fAtUpr9ovpftdwGTUq2AAnrNGEmppAKRVD7mmUCe+aN4rw249qLMcuZpeTZVr9DwcwNCnZu1GLbVHGlvaLjHmSwZNYPc5HFM6RkfzZJI5lc1aJ0N5vqJlVnUtMqZjVVbUB40Pq65g5xZ/CjngKI+X/g55zQG4GKbSlIam7mzvat4AX/S2F6P7k7O1lYMD/bFr37nO7JVf/LHfxarm41YWttUrklNyaDFhgDWI8OjmnNFPoUfILbs6gZ03aumBHUrmNfU2DjjxBKA1PAJ+F+alNhh8n1sCjOG+B1+uc4dCjCAjbaYuSpVhhHF9peuXBFQG5vFz0ZHx+PRo4cJoukVW6xy/JJMtkT0zjeMip9LZP3Nm/y1WoEjff2xvLTUlAeSUUodOetSUkRGd7gRI0MjSvRBs6vokVpsCsiygNlMiNMIqUCXBaL2G8d5kvjicEXdFaKhM8bHRhVwMj+CABfjgNFjqBlanvv3H4h90/sU1CHRgBOb2T8d0/v2iWpJAbxwGrdu324ihUDqYOhaHWMnshTN0Z8nSOY9GZKDAaUAS7Jj3VaGbmHM7WpJNlglNG4JIK5cv6ZAiAB1aGRY+uKy02W01aG1s4eRAT0URBcINVBPFD7QTJYe81e+CilthBHG2AMxSbzHFJSSnBYSGcPGa3htJUmFxlKTIt9f8k45j8Jr4iJ10dFJytRrSnoxBtDdW+NghCKUBM2WA4UcXEaS0D5kqdZBeq8rK9I3VoCcHWf2BrR5vrgmoVuT7YDjI5gCGSdWRUfE4vJybKThd7BDkOTnSkLF8COCfQK95hfNkJSXmdk3raYXxh/nQYGfjjx74N69e81AvgZMVQGuUB4Vxan4+RKror24/zKaPcOXJspdxZAKJvJC6+zoWWRBqob+ummIdHeXEjGCW64BhJbYIZKTMbPBwV+i94V6SYRESm78rKJiRRbNJmOTFeLARsXMthk0ahIwVC+T0vYh4kXTfnE7G2XPmlfjoArtreZd/UWhS3zfTbAJv849SFCmJG57W0g09hYB7fUbNyXhoOS1AaLycfT2guylaJVRJEF/tyVkoGqOjY4oUEE6QvqxQ0Px9ttvq2CtWTkzM/Hxx5/ElxcvaI+5gdmjggdFCJJLbCXSdZwFaOBicuzSasF+eui2dWDNQqu1VNE89UhdrDTtt/05OYCzXFE1ICRpklGx0B1CtrQQcZ4vY5ZCBaM14MtzVdK25Hso6S9kU1unqYk4yj1Ytp7tISRMc7B8pZsOvC115AYotpzPU+IEwit1ZPl9q3lSFGQzHXgGPIuSxZEmqlDcMLVc9K2GqgL0pLzb7jIXZzzmnxHQdXpuEDq/pd+dSDQjp1rJlRkbO7LNvDfPuRDUvJbvK5iuf9ufU/lOilQaoKxGemksm73hQpSTIaG3pQroxIDPdqNiXbbVw0jdyKpAXFrFuRe0j/QcLS0I2tna3S6oVNGKZ9XejHCzq7VX/DvLb+V20L9ufPl1P6vp8F8T0NSafd17li968X0BOISCeHybkgFQ+polYRSVmXC60kST2VZIDoQh9Vtbakq8/vobcfHi5dje3hAbgVdTXOnq6tDQT7TY7auH9AzX1jz3gDODXnhdM3aMQi++BjYBewdGRSHvuUcSJWKDx5KEchOeGMoSebtCZvHV3qgQEjV1xDVQPhkXxY7g98RFrAG2hgKDmJ4wKAeQtXyifeXGpJFndU5cDHC8RnFCZ4kmd0o/caI4K9xvNTZZNyRRuBf8z3e/+91476c/kR0DpQxlXewSDRO3TrWknJjHIdQ2IBgQ3Ogye/D51MRk/PZv/3Yitfvjh3/0w3jvJx9EZ7cb48PDo2rCyHZ0hAYgfu9X/7YaQsiAkhQOj47Hf/xP/zk+/fyC7AII7xrEiI2RBndjO86cPqNrvX/vnhuPkqbqin/2z/6P+Jf/8l95HVNiRwzObg9P5P4t0eOZIdgJNcWyAFisGP7lXsV6Zfjt3q7Yd7A/Nzo64t7ysppeP88vGCJzI2MxqCYT9mpcGsrEydLJ7+0R4AYpFuLcVtMLNLoHtK+srMfk5JT8IIN4uQeKsTQo5heeSot5Z3szJsdG4/bNm/Grv/ZrStDHJ6d0lt7/6Qdx4/q1+I3f+Dti1FBIYh/29nTGv/ndfx2d29uxf2I8Ona3Y27uUFy6diOera7F9P65WFxZjRs37sW5k0fiwL6pWF5ejJW1zVhv7EXv0HA8X92IASTFNtZ0L0+fPomBoWHdn9ayYy+I5R49fKRrATzEWeLc0OQiBgeUQkw3OTmtHAefcfzYMUlAHTlyWLaBnOHkqVMxz/y67Ua8ev5c/OjH72nOwdHDh+P99z+Mt988LcAEZ62vdyBW17fj3v1Hce8x6Pru2ERKp69XRQ0x9QBAaODnuBgBsK6HBpGL2JLvk9zrTkOFTORbKlZtSQKy1zwLSnMACx2bSOKSY+Xn2D/NyRL7gb8x8wc7YKq2C1bsF2LeXQaH9nQLNKazggZ3zr+S5MWuWc40rWCFU2yWbj7nu6cv9h04EDdu3Yn1rW0BRGwL3cirGAZfrxmEieTGhhFjUSAmLh0Zn8xcwwXYavghV0vMBJiMmM55zIAk+cjB7ty+K/vDfAqeZyG9YQAxi4YfSPYvOjTTBBTqbmM7Bvv7tYdu3bopQMA773wrjp04FvMLTwQQo3G0t9MdTx4vqODFepX8DWeW+IM4G9t/4/p1sRtGx0aD2Yf4Da5Z2v6dXWrict00ZMkzWAPun0e4vun/5oxgs7lPngGFLHw+to51QyaI98E/33twX80ZcpyFZ89iY9MD0D//4kITzMIZVtyysxNPF/BdDI41arzQ9o4Pa46DZ/5J4jkL4M2YJmMCP1cDxIilqxDchVyfwFGWkMLemZm+2Rw8TuyBvC6x0MNHD3XvjhmLuecY1p/xIsJbEZ1+VBz1F9HgZd9p7lA8pPEEmNGFS8dT/KX2FTOehkf0hpw75lvSHOQW8Vc0KhYXGE6+E929fbH8fC2W1FxBLG43JidG443zZ2VLrt+8HQOD/ZKB/eLzz/Wc3n77F+KD99/XWpArvPujH+nnr736ajy6f19NXOzMG2++GXdu3ZItOnbslfjkk8+057q6e+PWrduxCGO4v1fsLLGwGB6/2VBdA7ANKGr8dg3WFRhjz02vKvqTrxO7N8EpKb9o2RiYnYBuVp1Hy1chp2Sgk2SOurp0Ftj/7TEZtYYCcbCfyB+atZ6MX8VwZlHJLzscbzmGdL2kBmBnENnMYSSBmQxfx5mOTSrmlF2jiVnM/Zwd0MzJc/6Dah+5lbgO/V+C9lRnSDR/u1pB3Yvi/wQh+KJZkszNBQRyjtHOcGh+WFtM3MJofZWx0PL77Q0452XVEOGeSna18jwDnFxzoSFfcXGdZcXqCYwhHyB3qDpAST77fQ0s5MvNiBevscAYlRtqTdS8yBmh1VBIFQhLZJXclhmAza+sI8l65PXV7xQvJcismBWVOxZgTCob+YVNHMr5SpxB/CV2me+J7cgDYDxgR6n7CdyZeUxjG6Ar/hog4/Po7WFWWWcc2D8dszP749DsXPz4x+/HzXsPY70Bq/OVeJTz5WRjqQswo3eNWXSWMqN5ATP48MGD+iwkialPYXPINakfEkNRf6IWwRoCgkXumgbj3ME5SVEq39CAe1QaDsSdW7cVAzCThjhmbGIi5heeCYDM5zAXk/oksY5kV/eQX2cGT+aPku7NZiLKBN9IP/08Q+1v3uuvwwoc6XdA62QMWQkbJ4pvRaUkGHNx3FS/Mno6KKWVl4GHi6ytGRbSIQdBsZfaiUlB5+D3ZWebzxJyprNLSGiqmRehV3ZEnDx1UsESA8xwujQqMFgklwyiOn3yZMwcmImf/PQ9HXSSSILwkrxwst0wxTGlBzCWFBsLQQgDYX11TUGGUXyWH8CgoEMq9BxFHBWqemJ5aVk6xwTe6AA/W15S95M1wpiBnmw6x9RuhA1AUEcQx/2cPn1KAfCzxWfNoLFdwkfwm2ZbwcO0ST74W9acpJDigp8HCLrnSlRVuOrskJHlnqogxjNt18MtdIC1ih248ncEubwnyCS+SiexinkFW+A58wwxmA4MjO7idQRGFTBp/VOShSCToL1QogTmln/y35DsVjGc12ofrq2J2o8z0mDRvd14PL+gznfRrLlm3pMAia4yARxNrDLkvvYONbOksSntdxcjaFKw97gGOtu+bgdvDprTqbfJPmmPJ5rZv3dwZF1Gn+pCl1e9t4mweHEkQ7NYrNC8zckrCct9R2DJvSDTYCp2l2QKWI9PP/ssGTceYs95U8EoHb4YRYkOFfpEBeJ2y/NV9NILjQrOa3OGgM+247mW7qz2juaJWE6pEBNfsW+i+Bq1X0X1Ckrbg8/2v8s4sRVD1sWn9r6QCpOTceKVVyTpgPb1e++/r8KUEGCxp0SLQAIUMGtEcDz/jCDDxQQCAoIRrS0DJA/MxeQUzUsXH7ELnL0f/JcfaP4Jfw+qiUBKRfBuox6wSwydvXL5Uly5cqVZCFYjrsPNBwKWkkYzbbQ0qv2MtXckf+bzb5RlDSArtoUl+tobFQ4c/V7Y8jr3Jc/RPJ+JnKEoW6+XbWg0VGip5kV74OnFr+du9kLp/WvftumdNjtxe0YjOzkwKqhkcOrfsi/VqPBnwnAwAtizQ7qajArsOAmWm1wp5ZTnRowKodtbDUAKCxQTKuCWbXcnXsdUTdnm+ns9SPz4bGQZ+EI6So2/XBsX+K1VX8+rCrpeY6OVQcpY+snIId9rMmckS2M9X9sS1t2NIw1LnJzUWW+x7Ix4qoK8gctGulY7j/3Ce1FQQZcAf+BGUp7JfKCFmKoEphqypfHb8jmt5sT/iEZF7b9WE8iNCsu7McjOrIcm0h15EZh8WRDhTIJ+L7QV94mtILkpJoLmbHV1x/Q0hVL0x8did7cR92ANjE/G0OBw3L//wGCKlDTC52NXWF9+ZgbqXowjjTM2JikQfGedQYr77CvrZbuYjV0v6TB8j4vG6Hmb+VD7iddIPilRbkq607cUElBSi2kTSZq4lo1NmlyOY2Aqar+npIH9ttkjunZk0PbMYFXhIvcv54gYiL8r+QfWjz34T/7pP43/8B//gz6DRgCxDftsVXKctiH4aRUgk8lEgkfx0b58PV47fy5+/dd/PZ4vL8coNnhhIX7v3/2+ivvYYorLxHi7xCG7jXjnF78df/tXflkFZRVOtxoxMjYu+aY/fffd6OjsiXUNKWzNxBFzCpmY0THFhg8eMn9qWww6iie/8zv/q571hx9aW5y4AfvMPuJ8Eq9VvMseEGt30+w9XlMxTu1VIV6lA74X+2b2OaYiJunrjXkGL/6c2BUzIyOxD9DKBtIilrbD3rjYibyTWbQ8a2IdCqMkxpYl2NKcj6WlFaEIKYgtLq3o3h3PNyTxsr7xPMbGRmJudn8ASWGg9ZtvvSU/iw+kaY9m/vr6Tvz6d78Tr7/2qucoNZCpGY3f/Vf/Vwx0dcbs1ESsLi9poPUzCoFrG7G2ZZDTxto6TitOnTgejx7ej4l9++PR/GLce/w0Vtc3Y2J6ShryNCm2tnfj9NmTMb+wqIIta33s2OG4efNOjAwN6hHg55FoVFN2Z0d2AkYJ9n9yYlyDsE+eOCq7ymwB5kjduXM7ZmfnxKy+fOlSHDt+XA0ygFKz+2dic2M1+vo6Y+7AjNiZNISWllY1hPPKtZuxsrYW25IfBcOP/c4ZV5kD7ZueMohGTbyt1IIPXQOxAkURBjdjE6q52Bqu6nhaPrYpvelZddgx2wLHCexPirUAquTPeZbI/3Xbd9BM5PxR2OEVxCqwYHQmkYZVkZfCc288X1+Jwf5BDSE1e8GsrOXVdaHA+4eGY3RyKhYWl2NsfCT6EjyjxnHKPakohbxbnnkhPTs64v6Dh7F/bk73Wn5cszVSd5u/UXOwZDmRw+hmTtUzx7kdXWpI1d9j58kb1jfIdbxW+IntTUsEaV4eQ6lB2VMI3t6KX/7OO7FvhmbbRly6clGSaY0GAK9d5Xazc3MqfrNHifPwEdtbnsvDDDsK5HhvMy+HlZe6+ORzxz5EfhF7DIAFGTKYevgs7LkHmQMw2xBQjaI770WeDbtf7IyhwXj8+Ek0dvfEIkTGSPLCgKk6uuL69etqyBmQ1iv7iZyxBgdLwhkwUEk8ZdydcyrEsEwplULqYyvK1onZKeYmNtuDwHMXaj4J68Y+Io7lmvmq4jXxFnuGTQYiGgYKsxs9N8G22WAbx4WVMDWzig7iv7KoWbTOVzUH9+7sqlGERFs1V4mxa+Yae+fwEZgMj7XHyDlZH8mKaai7mXHIznFGeDbU2QeHRmJjq6FrxudsrK3GL7xxXs/s5t27sqPYjAtfXpBUHDN03v/gfd07zMBPP/tEe+6V4yfi6qVLYlaNjY0qPwHBjT1aWVmNH73749i/fzb2OrqU/zMzi248zAwYK/heYgsxnATec3PK6gWew7kwv5CSNwacVGPJoKdusVbIIwCV8jyIQXmOvAfP1IPda4iyY9RiFDXnQKRMqiRxkpGOf5OdoumU+QqsKyTBnBQ7V3Adwk3WKliriZDsRMUIBYpqe20Zu9qPjqcd40j2tAkOdJ3DDIuKVZFBzpmMbblU7SYB1QBQaD4hTbxiHNeMlpItLmBH5ca1IVv5l+/LcXjNY2jFrC2bzYuqcVJnyOyJllpUxXU1dF4MpybrIPPAnBPjuXS292IkpDKGmhxkjYq3dhV/qR7TTKBbTUHVmV56PspNc6ZQi0HSAlO1nqWfIV/cQ7FZdL2SnTaTuflVjaeco1BsFe295vu8OCdM6htZV+xW88v7yZ9hthG5uuJdzq3OiZnuNOyp/yGLNj01IwnAjo6d6OvBL+zE4YMHoqtjLw7Ozakx/fEXl6Ojt0+NYc49fnrlOTYf+UtqRVuqG2IfsC8wTPdNTcaNGzesBJMxOmxNGpFu+K3H5MSkloC4n7wagA0NZWbbEY9ojs/AgGbmwhIRqBiQMTGUAExjAnATlxVojdcCaObnAvim+kd/vxm++EI9l28aFa399813/3OswGkl0i16nwrPGLqUt2iow+8EWyh7ZIo4KDmnAANSQ5lKUqRkPmzwQCnS/bNsjfRcVVBFooihrh7aZopjh+SXNsWwQEYGxNekDi7oGB1CSTj0WosXHeTe3lhYXBBiuZCWXBvBN8FaDdwqXV4VM1KDFJSRHFtSdLdVeDDTgOu0A3RnmetHf5hAdHpqWtdHwkbCJ4cH+wI6Z1dXPJmfb9LuuBYSeQwfBQz+/tixY82hfwSyFEMwvDLecrA2yNXpZr34e3WQZUy7TMXs9NA5tHe5Hu6HhIekFJoqRk9JCwO0xYCxIbPj33XBRIN1c0aA/nUBzgiClr4jroTnaKptq/hVLAsPfPI+KQpgId655yp4VDFN6KrUUKXYQVGEYIgvPh+tXp4f98GeKF1DdKsXl5eMWkMPVjNH+hWMibkD8hhUZxryanwI2ZRDP/mXNaFQzWdBbabA5IFdm2beuLrTwvtUZFHNi3KcQrGh7VsBi4v4lTS5oOvXtKOH3Njwfi5WQXUQeL1ZEkYq8YxpxBw6fEjPjmCERgxOUHqFa2uiE6LRXM6cs1ZsDAWWqQ3bjsRmXxU6ol2KygethY5vL8jyq2ouqKCee8dDf2G3eKiaCmNZxLM+sW0BDl+MAemlZqDzwsp47epvVcBNJoj2B8EQAZgaDtZMPXr0mGSX2EO379yR3qsL0JbOmjt4UOdFc3JUzOsQKkPa6T098cUXn6sRBjWTcBJ+MgAAIABJREFUAIZEleRESLjoEKMH7er3swFCQss5R6OYggOFThoVLh7sxccffexElHk+kiUzyqu+hKLPomOrEJvrKqmekocqyZacoqYg3PZJcibNhKAQ+16rknVzQd060HypeZbPpYrYtqk568HVkKbcWPv+r4ZcRah8fnvwquD6JXQc61TIcX80iQta3J6D5Ka2Zd7UCBCqyrZFjQrmJ6lRQQORAm8OEdM12iZCl1eDoBhIxQ7TkN9hNdwpKnjCjkr8/t9E4Ffxn98Vw4ygHUYFZ60KyNr32SCQv2ub11HD7xKOJV8G6hObomKxPotyn5s6Fdw3r5tzo4GEbuo250Eh5SfmG3LoTlSVkHaYBl6Ub96XZ86+wl+CDGb/2a5XouREolBlrUZWi3LevhfLl78c5VRR/Ouinyqy/6y/+UoT7GewNOozXr4einCjSNFQGM9mcenjurjlJLoYC5wxknwPdDTaGBtBks8XDEYKLXwOZ50GBDEHyChkInm/23fuSY/cSEdYfX4t9kJ7J20lDSKhrEDPZyGAOAUUJ5/LsGBskfZpG0NFzfednaYMSDXE5AMTNVb+QAw2ZlH1eYbE1gYauqCPHZcNUpBmiOnz5SY4QJ+ZTA72LCzR0pmWJINmyGTzuqPVPJOd7bTcnQrYDI8d6BUD9X//J/9YqNDHTykESbBCyG7kYhpbgEC6VdAfG58QI4kGIcUgbLZR8A/j7/3G9yWL4WLgeux2dMTv/j//Jp6vrUYXQwrDUnnYhM693fjld74V3/vur8Wd27eE1sW29PUNxNVr1+M//eAPYgOJSUAWWaBQXAoim6J9zmiwhIsBBcRip06ejFdfezV+/9/9++jutWyY2BbZ1KG4yfsJ3Z2D2BVHSUrNAy79+N2c1IyjjIEoOiG9ucHAYgZ/9/boXpd3tmP++ZpQ+H+Vr77u7pgeGYoRngdyB0gprW2oaIg5HBkZk7QRa8mMJgpjB+cOxieffmpbhZSq5EuJVdG935Fs6dLyqmYl0NDy8NUNFXQHB2DbbMaJo0ejpwME34bmEvBMKZYikcJ8FmQ2J8Ym4h/+/d+OhfknkkU4cvhQ/N//8l9FX2fEoZlpMWJANy6tratRsf/QISHO93YaMTk6ps+C2TAwNBqbjb24fvt+dPb2ClgCUYxGhRkC+CrH4MSy2GhiH84wLGcKg/zfk/lnYkgyTFuyLXfvxpEjR2Ph2ZKe5cGDc3Hnzl0VETnLYm93dct2whDat29a/81A3ddePReD/d2xu0VRhOItRfHN6OkbiqXna3Hx6nWJU7KrFBelvFIHjKR0GqMagsleNqRFNkmMShcniJc4w9gmnhN+S3KzNAEHh2QfaKQZ5O4GWc2rw2aVlJvi0ASSFVp6q0GB3bJHbiw2lDOR57DPd2B6MjekFwAA7KrNGBjoE0CM/QpY4+nTpwJ2YQt6+wZwvLG4uhqdPT1uGiiP6Inl5ZRZFKgLFqllFYmDakgshfnegX4XtZpDju3XfE9u8pK7CMlNHpbz/7CxPOtC8FKwgRUmn56AIYOiyAE8c0z5z862pDUUXzQ245fe+cWYnpqIkbEhNSoWFhZjaGRKNgUGJkUmmhGcZTf3dgQcYH+w38h/sbPkJsS8agoq1HQsQuOLPA0fgf0HdEY/CdkQ3ovcFRDF0rNFS+CSnzWsVc4aE/fw9zTBLDvY6fUQe2/dc4ieLapQTT4kSTGtl8EKkodNBiu2zw1UAzyqAMjrPLuwNQOv/IBmzmUsz/rJLki2tFP3XMA4rhXbBviOOI7mDvEw7205POSWh+WPAQKo0F6yelnorXzFcZJjM0A0lrN1s509zvkwIGjULJTMDTlRvX2eRYnp94BbZmyOCNR4+TLMScs9YvPN/neIi3KDmnZ5DzThYOqJkfp8RT4PW7Z/dkZ5BTb8yOHDce3aVeU5586ei88++1Tr+8Ybb8SFCxd072dPn4mb16/Gxtqa5lVQxKcBRjOD5ixyUVPTM2pSbjZ2rCdAal5glN1dNYLIaSl68v7EEsTG5Kx6/gvPBBLkS7JGJV8qKVPPu+Gca87KgAFXOm8Jfqp8rGJ2MwbNzi0/plAzJcPMrHAjUjlUm59VvMa6ApZKBq78aCpYuCnh+ScFJuF6lReK6ct+daxhYB35gHNJ+S7yxbbCu94v419LrDkf0tyTrNko78H+cA3UedLZKubOe2wHTjmez3mhav4mADH/sBoBNa/CuUzLg1etpoBJBjuarV1pVb26rrH+uwrMYp+S16YkbQGIm9ei5oQBnKrRcF/ZYKyGYwGvqkHRfo2t/My5EOe5Gi7NuF72I6WDM3fxgHKDXVwct13HoTXzt7bZhbUs9XqTnFOKquoHzRVu/U4M2Hyu2EOBVwE0JCsIGyYGcIJExKDIOgL7kf/2bHEkyKjfEcuFZlP0dG7HQHdHHJ6bjc6uXdnYjc1G3HuyFB29yCW6ySPJJmpsYu43YuHZgvJAN0o8KHtm35QaxQVW4XwRS9BYRgaKa/GMw07ZZ+fsZueSl5EfqnHb1RljgK4442GmNfNymY9J0wP7TMOCz9GcXIFP/AyK8Vv70GycXOZvGhV/ldD6m9f+TViBM+Oj6tppMN3zNXUIK0FT8VcOzAGwBlrnUGUKcEal090D3dtCnRaF2fRSa6fSSGjsGr1AoMuhHRgYiZ4u0PfWD+/sQmrJn0/SiyMeIeEYHNJAPAryswdmFYTw+RxepI/wKWZsuCNOUEKzhQ4pRXsbNBexcX3qNkPfl4zTmgqfoHIYrqWAWjRJo180Jwktvh4PJoXKSYJ2+/YdFaLQ+MSQeAhVj96TQoeMdHaRKYRjWFiPk6+8ImQfQSaGF5QDQTBGquU4beqrIFz0XYyhnkEWv6G18RpQdbrnLAaD/CgEgtYkkwKCejUNYE6ocGYvXN1ZSX8QUDRlmBiC10JDl8alnEkiG6rwVWgPNXR6HCwqOFLxiAAZJIONNT+jMcO90OwxKtaO387Is0m4VpITocPyM0mWkdcQyyUdte47Z2Mg5YHDd3HFzBAKTSDnPXDcbA+ehXTO1TDr0jMjOamArVksazvE5XCrQK9AhBhTA2+NaKgCfxXZHGA58G7CnzUXxJIwRoQ4cuZvpHG7uqr7Jqn7zne+o2SQ/cOQUGQ9CJg3treE+iUBAEm5tLgUa8/dpWc/WV87h2ynhn+7xmXz+rKhw22CXPu6L53fpFQqDEjat+4hk3EXIe0oa1hx7YGSBnOA6SRIiHLNPEhJmYSGO1j2Whk5gpSCNYtZGyVeoHwpQm5tCeG0/8CBOHfubHz00UeyXwyqu3nzZiLhqyFFIozWNgOrjPaZnp7W3oRqz54AuQbyk72iRFoyID2xsrwUP/zDPxTzAsTkFoO1989qTSimsMdAY/O3V65cjqvXrup8kDwKfZsJs5D5Qvm6aVhFSaOAvP8rAFfBrS0QrpZZNY0q8K75CnoO7fDLIs83A+0XmTNf5dHko8yko4rK7KNqGr1AxdG1tQp1lg3yZjDSiGTD7JWyV81rL9TTSw1PbT8NvfYcFPY9kkZQbCugppnNea0ktpFNoGYDNRmBrAtBJcUCrXMG+Fm21zXxPLAB9dVeSKfphE1doRGdTSUXgSyv5b3uVbTdNsLJ9q87xifG4tGjJx7Cu0NRALYeFPVcszxDFL9Zs2bTpwGThKFsG02Go/wVjYoaXKiZ4B4crb0D/VuNQuZbTAq1Q7CbndBm46kaI9VQeLkh0N6EKIRSnfdao9qzX2cn6n3LttT7tX9Oe/Oh/fP+olgp86KYnppsngt8GPEC6w86tZpnblAYPQuiXYmffKZZXzxzCgD4fdaL80vhifciKapCFD9DYq8BunKdQlCPCmXYHhDZoB6FoM8ZTCQW0hHPwYLVBDNN3EO26znXWZCGbqMhO15fTaRfp+VaNHBvbVWJi+UZ8GfMInEsoESXBrAkEbeVKMn2pz+RLW0yeNqvwZIJVTAlPoP5Jd38PbNN2LsqcqkQxlbajt/4/veFwv/gw49iFKkT5mZt76oIA8eH15K8HT9xPC5fuSybJ5mO9TUh9B/cfRC/8w/+Xhyam/MsjL29eLa0HP/m//s9SeFQMCL+4rn2MDCxM+L0iWPxd3/rN4Xy9jkMzRF77yfvx3s/fT+2NKWXYaipo53sQYwRxRXFf56Vri/WCoTt7/wv/zD+7L134+r1Wyp4UZAdoPhBXs0SZhN3E7nC1EJvL3pUnFZJNPcjVu/6uhsqqd/Nz4g9Bgc9Q6AB4KexE+vb25KydHPd7BfiJGZ9DXT3xGBfdwwjoxMdirVpQtKkELMW9P6uGa2chX3TM4rh2QP4MpDd77//QZ4R3zeNfwbILq0wv6BH9rmru0+gFc7GJAOoN3mOoO57NG8CBGJ3d0c8X1+TbdntYGD4ITVF7t99IH926pXjcf/u7Tj5yvH4O9/7bvy/v/uvo3u3EUcPzgV2XQCT1bVY225EH+zpjq5YXVmKwwdmxZp49PhhjE/ti93o0bDqrYb0V4Qs5zNLk7qLH2JvO92U1/5XXNkjO7i6+txMtE4aGeOyAxoovo3klefxsT7Ms7p65aqeEbHWF59f0M9gYHBWiSeI8Xu6Il47dzo2ni9J31ozwYTI3Y7u/sGYX1qLi9duZgEpm8Gpu67iHrkOOtODQ2YxdXXE2sZabBET7xgZS1GDWEZnN5HDgCDwQcTKVdzjHNEErDlamhFT/jVlFcuuWK8aRgM20LHI1CSyp2vx6NFjnQOaWbBEkEY6cfxoLNCQ6Ix4+xfeiL1OZnEsK7ba2tyOzbUNxZiKafr6YxN2IgPVaRxt0gBzI16F7AIMZYEYe4a9/fzzL+TTxVAVmIoB2faHNfeFNQAYwhdNiyqM7XEvW9ueJ0QRfs85mrT9U3ee8wmjRn6uG3ktnv2G58owv4Pi+U4jvvXmm7FvajymZibjytXLce3mzZg5cDier23E0/mnAqIpH15dEzOK4dX7Z/Y3S2tr5MlIg4wiXbyrOJ19dfbsWeWB2BtARHwJFMaA6Y1VST9ht8nXkMHlzlk7Na91/vZkQ1kTzSLY2jBTHybbFkV+z4Bj7RYWFyVTRDMI20pMTbOYZlOLTV2yYc6rOCsVN/G9i/oGl3nodiHLHZvX2rOXWEM+12yIlI7KQjR5lRsZBtNx/ZoFtGf5zv5BcvAeyyiurtrmy28ZWMXniKWrHMP2W+oH5GlbBqew7yQZuuPh48TynBveZ30T38jcKHJ8rs+5wYnjJ/T5sJt53zWhq80m2dqg8T6gZgTvLbm8Pu9HS31uKUc/sH9/nD53Kp4tzltxoLsnbt24IdATqgoXLnwp//vq+VfjiwtIEHbH+fPn48Knn4gZMr1/RrE+s50OTM/E1MS0Zlns27dfNukZ8xaRbYIRsutGolhhsRvf/va3487t22oANpkrnQap4Si2svEk1nVKEeNLyZXIuZBSo7ZDk9PNbZ9T2ZScd0gIK5nA5+jqA4A0a5M1Ehsw6ywVO/IMFNeURFgi4ys/IXaowryeRZ7vYvpoZmVTptbNfksW8WzdmCoQl9hhkunK4nRK4ZWv5TqpNTjeMSDDzTbvKd1DsjpLMqy9IK/X8QEtskHeV9VfXoxKec6ed5bALs15MUi1lQ8kq6DWpa1T4NSq5mkkS0BzHmjSeN87B0nWtvIWA0abIEY1F2rgtVklfD4xLn8rVgy5TjJZMkV54Uba43HH7Gbmac5EMsYrVq34v/Ib/q2B3cpBkpVCTGOf05ptoQ8tUI7AVK25nvJTKWWolxVDtW0GIvbGeT61mg3FlM0aCg0IYqGMf/lsnk9ja11QtPXNnejq7Y/+3u7oie3Y21iJYwf3xevnz8SHH34cYxOj0TswEo+ercXmrqXeYahhC4hViK2pNzSVAzgn3TArduLA/hn5IWI8fBn3jN2Tbc0GkKStyPUTvOC+nucFqalE03V4WPb+4aNHAm7w2PZN7Yu+gQGBQahxegbHThw6dFDf44M5Swb/Opp1g9w1MtUDvmlUvHhwv/mvv/kr8IrQ5cwusH64NQGNXhVCUWj8XSXzok2GkS8K1tc3lLy9jBY3ejaN/S5onq3o6+8RDbkQRR0d3TE2SpFg2wyKrg5Rzg/OHVCQgB4bn8EQR/6dfzovpBgIBRoXfCYzK2RoO0FF4Ix3mugdGdYqICnw67W8iejQ3bGHHrV0RV305MgLzdPZqUCT68fgqXBIgIuuY0+3CpM3rt+Ip0+eCs2joIqBuRQKoC33mdaL9a9BVqBn6JAyCJJ7o8FBMQr9OlBwOAcQF3IKhR5v03B3wMugPCPHtOYEhRSlNxgy7sKgA75OBXAEtMXM4J5F/x8wy0SD1jQc2PNDaq5F/T3vhdElyWvSsBNBwTNXJz+LMW5EuElkR8mwSeaBuPngYbB7CrZ5rfZOFvlAjZQMUzlPOTsQZEmHRhOZoLeCWb0XyMUOZnYMaJ0JwijoiH3Q0yu2CvvXaOJdIQFhZfBcoAzvNLi/7VhZea6iNDRBklPLhrxAXPwKo6ICNjVGCl0gWZusKsvpFwfWTQyjvHLmQAZfZNXNgm6iRdjTBKQ06bh/3vOtt95SsYHnBoUYJ0WixpBSEl0Ka/wN55ZAFJStkAmi2rsJRWDnBDi1FsWwcNCgAWkK6ho/s1HBhTqIMpWU9xfzJCncrCUJt/R9hWBzw9Coj5Y8jdHkLcqx1i+DtxeB/CWXs2fpkETby85UUX8PuYtx2YODh8yY+OCjD+N73/uegg3YD26Got3eowBCDRIVBtDo3lWjApujIbusHUEK56vR0P3xMxLs+/fuS+aCRiGDdvv7B2N6ekaUdvYhUhdnzpzR3/zhD3+ohMP7oYUOgu1UxfRCs6gpVkj+pPAW7bo5MK65rdq6Fm1NzFbzzEFLq6nQos2/7KWyJ/T1zqttuPcLTZCUN6vP8If5HvW/yQCrIF5SDtlwEENNyaltlJtApigrEE8aMxaXBE0yg9L3R3N8T6hsDcvNpomQ4dnkUBNMwX4WoxOFxf7mDNGokD8Skt1BdJ1w9i/BZhWG2wvsBJ7sH/SBW7wq+5TW8D+jN4t95vdpyOYhe0CRm8G0nPO6f6F9Mhh3YNnZZIWwpJwW9ie+CJ+rxFqNii6daVPn3RCRf8MuC4XlBFOyEshVaBgy55x35DOzUZ+o2/Z7bf++nk/Z6NZ/v6h1WwnM122iv0yjopkw/iVDqGpUzMxMZ7GhoWJOzTHinHPvFIH4fAqQFI82tmynhM6VnIgbFfZDHTr7FCxA0d68dSP6QSGSgJAk9fZoaCmoc6E6JQ83oMIe+xE7rOJ1hyUKjdo0gtUgjjXLsXR1NQtX1Qyr+y9pKBoVtdYlLcTSuFmH1u1CU3KI68LewNxqTySLwUgcwlchxNgg9s+lC+6jWw03moG22eYeUdjs7CD2IwEzI4Si9clXjsXi4lPFERSB333vJ7GLJIWakgzM7ogeZCRB+e7uiOGxRtGbggfswI31GB8diWfzi/Hbv/m9ePutN+Pu3btx9Nix+Pizz+OHf/wnsbIG441r79W/Glmxt6OE83f+4T+Io8eOxpbWdTAePn4SP/iDH8bjJ/OB6OZGykjSgOKhSAc4te5ZAw3+3vOcCTUUOjvjW9/+ViyvPo9PPvsshkeHpbvfo8Lhbuzl3AZgeqyP6hkvNYPl5zjPpbmekgpCrvf3mTGCZONgv2IADQ7WzBQXNOr7KlA0pfKQbxHrwm0RgXJWPYxYiPFtN/t3ufO9nejr7Y+jR46qiU5TioIrzTQ3TntieNioWp7xbmNLMeK2pAgHZCOIEzSMG4ZOYyu2KAgzk2NjPQb6zMAdnRiNQ0cPx63b97Doiptu3bobwwODKqB3BWyAgXjnW9+K9959NyaGBqIPffqujhifnoq7Dx6qUbG9R5NpIJ49fRqvnT0j1CPsnOhkjhDxXUfsYvc4V+urAivhT4Q0f+5GAc8EdgiJO0CCmekp+SHWjLVnnZF7/OLCpZg7OBvPFlckz6Ti4pcX4+iRI/Hk8WOtDz/78uJloewPzOyPzy58GWfPnBJo5+qVa/Fr3/l2bK2vRG+X14OcZWhkNHaiK7Z2OuPy9Vuxjr3ehCmhiowlW7a2VTzu2NmL0eFhxavMEGCO3bKk+QBf9KpQqIHfmn1n30aBlbkwNKTEQk+WADIP2AkNox8ciBWkgwaRSOwUIp9COPdPPOv4j5Oxq4K3z3Jn3Lp9RwPqD87OSjMbrf5jRw5JCurooblYfb4sO8qg30dPluLg7HT8wptvqVCDdFOD/S4tjS75GcBaQtKnBE0xqMWMkAQRw077bBPX15S/qfm503BBO4tUyoPaGrY0wvDVyk9ViPSg2wJAKe7cS2R2cxhrCNC2us7cGcco/DvY1xsTo8OSMXvj3NnYPzMV0zOT8eDRg/ji4sXo7R/VnALeE9QqZ5piFCx5rvHg7JxsOw0LCmQgbXuQBln3AGLJEh+Y1WvJ0ebnn+VsADs4Zh8hyYctJPdj+Cr2kaK0hporXwTh7ziPOGJ7l2bWroBWnXuJuB0cljwQrPLHj+c1XJ7YgEIbuF2fcdspsbw0DLnVSKpGVjXTiXH4khTJ4GAzj6x8stwz7+tY2k1YmKb8bTWdWBv2nNlA3s8CNdL07rQsFpKWsKNWlz1QnFiX9TPyHsUB7NJQbG1vNqUxad5gW8QqyJknxHUu+Ibs6l44tnFxcE/D0ZkdxevICzk/yPrybDSnUTPgKHSakcC+wkZzDnlPrksD1dc3XG8YptHSGQdm98tf3b5xU0jn06+cjI8++ljnEAbShS8uaK/R5Lx26ZKaXeOTBhSw70cHh+PYkePx8Ycfxdj4pMB7d+7f14wKGUGcExZfDczd+KW/9Y781JXLVzSn5dnCgj6Lc42SgxocAo4CpETyCxaKGfz4BrMuN3M4/HqCh9w8cnMJedw+z3cCtJe+S7KZW9tpd2iybWS9IEGnfEYWwh3TZ26YzLkqfhfLoFg7NEFq9l6xg8V11pwFNwGwczyHYhmQ7xn05Ni97qtmMlROoIHjKXtWr2+CmWRfUj1DftdsN35f7NZmTqR91QKK1lmq/LTFNPL+s6RtSfOmDG42F1oyVy15Pt+H5XN9zrPJkZLIjh3NYKjP1p6ohkKyeuu6FdtRX0hGTeUW7UCqfCfv9QJs5TMrMKP9jpUC9HkZd3gtC0Tp3zUBU8wjSTURLrjyqJcBc34/g0OqdlgMrfpc/T21kpTv5TrVBEiZVGp1nH8appxLgIE8P/Ymr5NkeWNLoAVs4sbWbgyNjsXTxw9jbLA3ene3YmZsIH77735fjcsepDB3O+O9j76I1a1dMdxo1j1bWlEtkhh7374Z+SPsOXZ5P3MnOhyTwxLED2jeC8DbwQFJOPLcPK+MOpZl5PD1MBNpwAsosQkoYVM2cW52VvNqPatoO0ZHRmNkbDQ+/uRTz4TLWZabG1sJWGW2VA5az5mkzmgNlFM+/k2jotzWN//+z7ICJ6Ce4ux29xQ8SLYgh1LJSO1YJ92Fp+zUts2qkGFLB1KD3zRgtch20K8olnRi4Jj7AHagQ4kmKDyo1CTz6EF29zCgekYHHAkAHDySLry/h9bYqVFcBDmGgYZaKtZHZ4cSMxckKKRiwIxec7c2JQ54D6FTCX5Nj5Q0RA6c473QAC2GQG9q+/YPDcT0zHQ8fPBIDRKKoRTkuaaxURdFCMAJjEBPGOHgbjidU4w7Qc8XX3yhgI/i2+FDh7TuGgpO0TaHVbuIYUdYjqSkrFz08vVx7UZ/GD2Ko6/iLIa06JcM8ymDV40AUSOlY+m5ESREvAdJIHugaMzscwcANcy1JQ0lo9gcTpvMkyyAVyApBIf0qZ102xFn84JC8Pqa0fNZDOf1OB3WjC4zBSPMr+mQyBc0VCgxg8QFGJ6zqbKeZQEtVntq07IIBPqgC/kiGCeopxBIMkbASbJLU8bXnOjm9gPejorIho0RIilf0+Q6umzrl6eEUbIIKjgpxIICgZRNqs+UQ096pwY3qpjWmRRt79XHT54oGaDrrqJc0tNBmMEmkeQQgaWky2qAFs80ZUqyEF3IKO21QnkQLH/Nl9EzRfM066kYFm42lGal0fd1/woE2yjCrJfmMiQNWO41GxWFTKlh7e3UUunxU1ReA1VhPWU0x7ENBA0Mur5+84bWA41pzlYxdQjc1WzNgZEVSJC0iKGBBnpevxBnGm5stgP/z8+8J33PINVn9s+ZWg3jqtGIQ0eOxMjIUFz88mLcvH1LA7wIrIBUVcuq9FUJ5irArSHnFdDycxJl9lazkPtSo4Ln1l7krT1bUjgvFJ0d4VbE+5d2WW48ZPOtbe9LSqvZmmg1KuqNVbxVYZ5kEcmJ1hyMssVCQyclW4FzG9W8owM7TVHOhVZsew36FPOgbS4E2a+G7Kmw4ABcezLPJOdvdGSk2chVYTYTi3Y2STUqqkhca4udwO7hU2qPNhOSPEMa4pdrpX1FEyAZFQSZSGYUqozn4yKjv/B7JcNGslaFAXJVCnIUyYSMzEYiiZgabe2D7HJNOPuSMaR8TqGYRnbRqCXZ6EHAdeYrgWunvnurtBpJ7Y2K1j225nLUz17eVM1CbiZX9fv2hoc/62dxer5+m+r6oyOmpibUdC+/6OTV51u6yck6EUIZlGcPKHnk1xLNlGxO+ZLNrZie3iffbYTmkN5rLXX9ec0KKPD1NZkInh/sSDUzNOy8ISZnFXHc2LLERSXWNEP5XvIpOUC7fU2wX6xFNVgq0az9UBRyIbzS53DPDOj86U9/2pSTal+1WlvHFC5kVLPGMV1KPCXKjXPrweD4DDdeujqxYY0YH5t0gri5LtT1wwe3pasLe+zP3v1xLK2uyhdRIKaQSVFWrCgfbsUXa9n85f0pfqMf/9q5U/H3fuu35N/x3b//7/5DXLtxU5I/JJqbWzv6F8kjCt3MSNg/PRGvvXpeBdzlpZX4/MK7+mPeAAAgAElEQVTFuPfggYqJxDti1cJISnYMMYeS3+0dFXy8hzp1NsZGRqRRfpAYrDPij/7sR5L2NEMJ5Id9uZmPnbFn3Z6v/2oDN9RMGCGEVXAelhRXDa0lhG7J1Rgs4LOZTKtOo4zZzNZ1d1OJIqaANjuWLuEL+SZi6pGRwZyhFhpoiz0oOTpiIr6mpyclfUnTpzN2tGb4xsYubGTeC9mhvWhsbWp23PrqsmpnyBp2wABpbKkYxlo9ePg4evqGhQYHGUxhDamUvcZ2rG2sxsnjR+Lx/QdxcGY6NlZWYrCvJyb2TcXjhaWYX16O/uFRnYl7t+/HYE9nnDt/Oja31qKjqzfWN3fj+dpWPF/fiEHmt3TsiVHBuSKpZxgukimc7ZMnX4lr126IsUGDhPjHwzRhPGwqtrt+46Yav8wJeTo/r+GVZjc34tjRoypanDp1qjkY/uDBg7IHxMIz+/fFytKz2Dc5FgM9nbHX2Iq+npz/RT4R3bG9S+O6Iz6/eEV/k4KTamIqC2rsRRd+B3+m+UEcrpDUGMVeGkzcG79jXzxnHfGfW8yH6FMDVdJQAozh3/zsidmJmWCAlOQOdv7EiROKAR/cvx8TkxNqPSJzOTu3n3Eg2mcP7j9U3DI5ORFPHz+NsZGhOHL4YEyNj8fa8+W49OUlNe3mDh8Uq+D2zTua13P+zFkBfeYXF8WoWKGQL+klI/clydXV5SaYUNDZHM1YiufCWa940U0MI6wVG2aRivsXO4L3oGGY8wd4HX6ZOQgUYGmQargvsod7ewJ9kd/cf3BP+aZaegl0Gezri6nxseja3Ymzr5yI/TPTMblvPJZXluKTzz+Prm500f03nDUaO9gJCtystQpnAqbtiQ1BfqqCbzLojOS3NKCaQ9QOAYKBoE0JQmTMiGFpmMEokq0nZtg24IECFzZUTbmhweiACbO9qXscGTarmqYyxS/iKxq1Ypcgk7uzLYag88Ziepo5zFfF4eV7q5FRTAveG19kO9CaweV41UATo/HNRsdfFcPCOZjzsYqnmv8tqVWK5sx561NxjhyNoh5fhZ7HZ7a+t8wU14GvL9kmgdMGBlLCyM1b/HY3dnuPNfS8Bs+Dse3neczOzqoxymfevnNbTIPadxWGGDBn8B5rAPCL2BK5psWlBdm148ePSe2BBidNNICHP/r/2XvPJzmzLL3vlPfewnu0RZvZJXeXlLg0iqWC0j+qCO1XiVJQohF3dtbMTJvp6W4ADaBQMIXyvioryyh+z3NOZjame7kMUhEaRldHB1xVZr7ve++5xzzm5z9XzX/37l3V9jyPTz75KL76kjXFcGNRe5R1sji3ENPjU/Hb3/zWZunRFS9hcKUpNmeYJJCSCck6efDhA635N29W9Pn5nJzHO7t7ioOqB4TicG0lcKE8JRheI+VHn8JrijVGfERujOfEn+ueVw3CPafJqhotTzuDMe1dWTm43jclwjtzOw/02wfl27kz38tZ3JJp6vLZo5y4TJk7fE6Nwk/T7zPkqlkbJVeZ4L9kRKi3UJ4NBc7okMMT80Brou0z166zLAfg/MuDeefrfg/9n2A3KVyo7i0mhXsyAqYlSE/PQ78366LFjOjIIPzY2qwn57Rt2ehWD6Hlw0EeZ+ZE67UF0Gp7RqiXILlY19bVR6rkxYM4s04q53Au7wFJSTc7TmTc6PDLUH2VMUZChyUb3jkEqR9+K1uqdZJNo9bzLlaL2PcCTTvXUg2WPqjkp8QB4oSGt/ISI6f3HlB+iwJC14V8zo6bFzE9Ny9/rIGu0+g5bcaDd6/FH//hzyTD+puvvolm9MTTF2uxc9SMa9evSSISoPGhYnSvABJIWxLnkYVnP7E/Z2Zn5BVBjOaslaz00JByfK4B1hg5MnsO0Cn9J4Yr5BYvlp+rvwWoYG52Tq/F8FMD4/MLyVVS6y0tP2/1L92naMqbhn1bwPFaOzX8Mhvqp0HFj2TpP/317/MduDU83NIbZLOQ4BfVk2YbsdMoE58Gonpl81/IpgxiMptWM8YMjBaC/MIHGg0DDSku3Gzp7x+KkZExGYHpYG02YngEZElEo2mdS9gUFBa8mhEP/RoCINUiWhaFaNJDlVClPmOhOTC8Eqo7kzU1UfiMhEIZjhlRcJ7a50oaNfW1hAMIJJrdJEuLVy8LfQS6WtS8NKXkuo046NP38bmQ5xErAFTGMfSwwbh580Y8fPhITWQCH1/zC/MtKiYBjwO7kNwceDYd5hqdQIkqm/QxswiMTMJoXNJbot8ZcV/NGx30eW8K2SsEBAVyornVBE40l9kVThy4b4Vc5nUlO9Hfr19LnodfS4KJJEkJMCj6lIaSRJR06J288Dykq5vNTO4dNLh6L03Wu3s0fcack+fT+sqpPQWEaO+ZgEEJpNjT+j06FpWORJP7QbLKYINkkvfm8GGCrecLa+P8Ira38PhwA7iFeE3DKR3i+QG+p8fYMvVKYHl+YzXq3bBrIzPUjCi0AoyVlO+qBELXf+rkkPWBySgIJDVHRcd0EkVxO7+woN8zWOTgkoFro6milu9nyLP8Yjmli8xoaICqSoSbEUwuYFqSGGqOu/H6Q1/lQSIUQRaWnQbalndLn47U+3TDvz3I4Nl6UGFDLjfZ3bTU/U/9/vYdN0NIDV1JP7HHLUVy9coVHfyglrhnmFutrKy0inoVi7yPKLhuInMjynysCkMl7GIHeTggbw8QpqmRyWsgoVCyaTMzszE1Myf0BcknKFRi1ObWRnz5xRctnWmuR0g2KKlCbFFg9Im+SrJNodRqKJbME4OKknKpAUH+2hohdSSGFX9LakvD0Y6HV2wL/VXHv3U2k3/wYZc/yVuvVy/e+VmKUeGkOJkS0tQ80f2uolf6oZl0ckntpiv3yR42StR76Ah7VyBNwfNHrqvMOC2vZiZB+TJYo9tat2YPSLMlpiYnFG/rPJJtdcpO1ZorBLziXO4JrqTMSssbqY0c83CyvUY91DGqzAwaPjMNbTHruCcy6M7uYibxltUxvV4sP6FFDarTvulAcIuSnYMKxaiSPMmCiZ8xnb/M2I1y93lN4U1x56fWllgo2rD9kH4XgfX9oUStkx8aMPzYevqx7/2hv/9P5VAq6i4ipqcnhTpimEARDuOufCiqSGXv0pzT5+pyvKhzhIE87+/m+4mH3oODaQw6aJDEwYGeH2sOtOP+vk32Si5jZGhIjYpmFkzIMtHk4dnzzFvIsmREcG0ULCVf4yXgeF4/R+Onhti1jvi1GBWtIi+RgMhLfPP112ra8cVr8/0V9+Q9xTrJwk7FnO6H14rjbfrXnNs8tbffXlxGmrIee9T0np+dk3fB7VvX4+BgR8M7QBnLr1fiuNmIE8mPDMQohWV3X2xjIt+DpMOpfrVecrfPHyRGukLDno8/+kAswa+/+TaWll+pEW5WBI238+gFUUchSr52fqpCDiNs8gf2D+ua90Wej4gxPjGS7KIeecS4SUPj3wwkSdKkVjBrCW149u3u4WE8fPJYeZPuSaH6uizroHwXxVKakR38qlqzHkIajVjyCdxrUPY0y2nOFkMZ6SWxnzpYx60hhRCtbhLB9JWkKtpDDBKUk4G6xn/LMgts8bNzDOLJm9nPbsAIsJPvQWxhqI/vAo3vi3NYfAZ8SIeZwUcaRYL6lgmreum8B3r5sDWR29yUmThSJuyJo0Yz3qxsSSKMM2tybFTDCuLtxPhILM5Mxcnhfly/tKjcHpPafVghp6cxPjUrOZOLZjPGh0dSY/4gBodHY3vvKJ4j/YR59nvvxNburhoAhGYGFbu7+7o+ZBpAGeMvMTiAMNaFro8v2MnjE5M6Q2DNMiirhiH7nuHhixcvlUOwxxlMLMzNK/9GngY5ya3tTclI3bpxNboZ3p01oq8Lls6ArrGvfzBOmmdxGtQ1PWo2Pn66JCYIz5Y9wTCCyQVMheEBck03dKk/YMcJBJH619p3SEnOzGrYJHZn41gIfs4TGNzkxEjoHh0cSQqC3JncVbFNg9hTDZaolbi/kpVtHAsaxvAAFigAnaWl51pfUxMTYqrjT3H//t2YGB2NlZcv4s3rleju64nZ+XkhTVdX3sTu9p4G4X/w8ScxNDYaL1ZeBepcsP0YdJplmIA3msKYKg+Z5c61FIJaHlo9PcqfqI2cmrjxxrpGsozfAzYS6jnPU635/n6tgTerb9Twt/QFzUczYgVqi4gXL5Yz9ntYQOOLQQVrtPfiPO7evCFGxfQs0mAn8e3jR7Gzg4xUv+qFLeQ18A9JeU7VmjTSkWVl7Q0OSZYJWTLqjkKot2IcsrTpGUWtIqafgHj4BNBYtCmyvARgTV1gBD+hHLG05sV2v7A3CZ+RuMp9I6+iScb6ge1npmjJNDmn7JS3rSFDyRDWGcOZ2FkDEDdYIyVdWPmr8xlLNdeggudZg3XOHf7MM4PhXBJSDD74GRp/7C9MuIm9IJVnp6b18+w1vjTIKZnU9Eess1aDeg2BnLsRY2nW877ke5IC60dyasisjEZTg0n2vaRWzy9yTxzGnbt3pC3PGVSgQMkm6Uw1A70GZtQDyCZ99PFHGh6urLyMa9evxo1rN+KI4TyyoHt7YjvAiLkHw/Hzz3SPHjz4MB49fKg4AJvr9ZsVre1xfDNm5+PJ4ydiJB4cHcfa1pbAEDA2yBN5X/ISPju5Cb+nd3D5yuXY3dmWHB3nE+uO88V5oR3YlG8zFE3gqGoWmBLKD3vU8zBQyzV+NX6VJ6qmM9inhkR6yZQCqvWg1y4TdPl9pC9EAmGcY9vzqkqYes/yPmFdVBM81Ws63tceEiXxw2c3+78tQas8J3259LxUN7tBLynnlIgS6I/6ET/OlKvSYA+GU7JpfmdQIVCkAQtmLdTQxZwLDVNbktPtgYz2bf59q4eQg4LWoKMutiPmCUCVrJFiFRSDwXmic3r3d/LeULd/DyTVORjimaQfhB5ADiySea6YmTkN66CVu2et167HPZwp4GB9zorXvhdtny2+l7XoXkVHrdOR2BdTuJQddH0JVjNoC0CrwVk8b+Ks5Uw9bGPPMzjnnshvUtKADDMNZtWgC+Y4QJdT6naISucx1HMeZ4d78d//8Sdx69plqSJ8/uVvY2hsMh49ex2Hp6GhPnm/2euWW2TNk0tYvhcfp0ENsKemJ+Uryzpnf07PzOjzMZDki3P5zp07kizmTGYAyRnBIJ3eZd1DhhuADDhTvNfsf7e+vhF7hwdt6TKtgy7J4Yk9g8Tl4WH61Lq+Iz9yf/AnM+3/VC3507//Ht6BGwM2SaP5LD24nMgLbQWyHpRVGlcJ2YAGZivx9MEuVIOSRUunEAzZ3CQpfT0D0Tg6Nhr+DMRNiDI7Ojwm+iN+D9Y/BjG9J+TW1MyEmvhMG58tLcXrlTcqHq7fuB7rqxvxxeefq+G3tbUZw0MuTjVgSDNFI4/se8GJh96vg6KbMioULs40+QRFSSORnz862Ffjw5qPSBgwbBiOd997L5Zevojnyy9yggtKs19FAIaOJF2TE5NKNN20Ct3PMjUD0cH3k7CRuHLQEYwpsviZkiwqNIzRjySmnrZzqKrJPmajLwITwx0kZ5Q07u21Vh4JNgeCP4cPsDISrUaG/i6TP4pMHdpCG0C5dFKugyh9Hvh+Je3pV1Hou2p4l0m3EFJJh9PApEyIcvJea6QMsCjgQY5V0S4zbnQy1YwYkOwKEiqeolv/j/vGvxf6goTYRUyfAr4S50Sa2Fw7YnZutpW8cN0cSKwNmpEk/RRNusaUj7HpmL86G78tnftOzfv8vevT77MpOtER3wcQO5EotJKQLWmWy/Oj2UUxjawT1841cZ0UAtzj8YkJJeZ7u/t6RgwmaOaC/GVN8bo01Hd3t4V0rUKgqPjtppWTESFRaCI323r9naGMQotiqaSxPMG3TqYSfBk4p0lsIsdL2qJQ5G6mez+WaZmQGdCcO2j7eYq39iufufSJZf6HXuOVK2rgPfjoIxULIC4fPX4cT589s3cK8lSwIHrNhDCSxsM7ngPrji8SDaFmc4AhKQESkqFBN4eyeBJyDLQJhoEjo7FzeBhT0zMxMzUteibP5LvvHklX0uy0NDrOQRANn0I2Cd3EAFj+G06ESzbNiB1Ttr8nQPY9VgPmclCWk3Zc8lJ5D99uGisG5M+XXqy20fdW9lsHVw0o3nrfzj8m/rfVEHAz0Im00euw5zyAYn/ys+zptz0hqgDSfuhzEe8mqk0OOUdEvU1DMq9d08TVXE92Dn/fYlTkvpW3izwqUopM+qrnHuTmfa4rL7mKipvVVC55Lp0fSZeun9H60SDRxWI1+41OYgDh99WgIin5KgTy72wK1619x37hGvqEvkJ6xsWX1gTydVWQJjDAjdFewaELRVUofiMs8z56pVvWRwNBAAXtoYpiXAdt3H+mAdTB8sgH3zlg+LHhROe583cNKjob73+ftElA5K4uJfvQvjlzKcJZU5LIyWEka8DMJ8eyMsK2oSuGn0bHcj/Zuzo/TpEgOYqx8RHlKvgFlGH1weFRbDEMgBnaY9kOnpFQvSp2vb+IzQINbG25aZ1nlKQTe3v1eQ3k8LOs39cAnThW97Qad/yc4svpiRiP5GHVlPrwww9ia2NL5q81DFQzMHMcAQUEJGkXu9VgEGozh2EqyMDYp/QT/ya2Kf4yPQBILmJuejp2trfivXfuxocfvhO/+fLLGBoZ0/D7i6++itHJSaF6N9c31LgAdSokHANITLRZ4w3LbPAMYVWwvvv7e4Xe3zmgQdcjXfxG80zPjAHE8MioPBX6e3tigUY7clwpqyNZi5PTOJERJyCRgdjb3VIhd3R40GrCIe+kfahmoCWEiH5oA5M7cs+OaFZ+91DDRM46DeU95rMsInsnB2VqnLwVF9WsSdZnoQVbwws83/oHxJrtNK9sDyeSQFEDaWDXejU3fs1ysdSP2B5KgQwAUK52hiRCj5DYbkJ6yAqgpLT7GTbQrdK/nzHoIKfAMwcftyMhCHl+avSf+7ns7SA/ORwjQwMBWPTgYE/n6tjEmD7P4fFpvHjxRhJh5PCsX6STZqYn4vXLFzKtPNrdkgfF6clx7AI6GR2NtZ3dGGAP9fbF0f5B3Lx6NU4aB3HcPNKAav/oNFbXt2L/qBFTs9Py0QAogLwTqP7xsQlJrZJn7h3sa0gBEIozluY792V5eVlMKeqPa9duxC/++q90BiARSXOUBgEszC8+/1IoaZDKxIGPP/44Hj56pOeE4TbmuAtzk/Hu3dtxwNqSXAMDzoY+w/b2XoxPzshzj4HP0stX8XptU2uewQwsDpDzzeOTGBkaEXvz5PREUmegPsnhd3d2WjKtxOZLi4sCRPHcGTgo5xgd0WckxpCjEHeQrtra3pIvmc4qmPAwZ2ZmtM+IF+6LIQvDMAVZQPvCbWxuqlmLlAWMCqS9Pnj/XUnaHeztxfLScw2COYHeuf+OmjDLz5YVBxHJ/ZP/7h/HytpqdA/0xSbx7szmnpU/lwwrABrOO8nWbO/oLPe9vSIwEWtPrbRMtlnbDGAYSLx4vqxYhsRZtQu5TljpgNW4jmIr4mnDc+d1eTYM1ciRQNobaY5IV0Q/5qXDw3H7+tWYnZ6KmbmpuOg6j9WN9Tg+Oo/NrV3VI3ugZEG44p2zvaNhEcwK1hxNaXnexEWMTY6JKcDnJL6bfVlM6QvlmRoIZAOYHLKAatSDzr3Jb50Xc33EJHIn2AdI8BVzgaY5a4Hz7unTJcVoUPUexBiAYxS4WcC8dg3o+Uw1WKhmIc9U9aBqK/t1OaYaNFLAsZJJLNQwa8/fE2oUch38vId3loKiNsEHhZoMkB4m5EgXYkQOeI89wdBNIKs3b7Ru6rNQGyJ7xeuQv/E5QR9XjqJa5MTSxZaodp7pzzmYzTvWWZ/OdCOvLWU8OTEeH3z4QXz7zTeSoCq/kAKyGLTV5cFQ1sEwJbi2w8M9XQdnMGC4P/mjP9J9+Mu//LnOl48//Tg+//xzgR7eeed+fPHll4FM26UrV2L55Qudb9OTUzE5OhHf/PabmJqaiaPGSTRpjNI7KeCc/JfO1dsAqMN9Z+h4+dJlyQCz5797/Fjob2WH2dRXviGfmAQKZv9DbIWU7lHfA+N1/Lwk1QuQ0+dnsWzrXhSbt2S8qvlcMrkFwCkWQuWqnPWdtW6bmeAsTwOo9LMxW5jhLYyPGhjZtFv1pe5F9jBKsikLcjP6Dbap39eaVR4t0IFBPWZeGTwr2SfOiVINKfZRJqHOS9teja06KZvn3iv0V/wDaq6fOqdwXtBmPXj47IF01cOV9xVIjzhP/WCZTnuy2PC+WBgGT5a8svPzkpgqgJHjfOUlNhb3ffPyKFq++xM84wJUFUCQe6Lft1QlDGas2olXcVxxfeD7pHfImjulh8ntOkFZrbzGjXh+pIbaAkhltlO1m++VpTFp4nNP2Me8jMBDgF9SrcTDbQ//+ZW9id/Vzt5e9A0MxST+c0f7cX68Hz3NRvzpP/4kbly5Io/Tz3/zdYzPzMfK5kE0kNU7OZXkktiLmNkfHKZUdKgPo+FXV7cG9wBcX7x8JYnByfEJ9ZeIM8+eLuncBkB6+fLl9LnoidGxEamD0C9Ub05Se4dmTE5P672IadwD1azHR5KL4s/EIvYiZzfxjTyQM7Sk2hiOG3hcg5qLn6Sf/j4F5U/f8/t1By5396ioF9WRJij0z8aJEAlKdoTcciO4DnH+rEIJg0AZeKGVaNo9gQ1mQbsB1xunJzTuGBCcypSazIpm00D/kJruDDdGR/BfOIz3338npuemlJRjPqbmZJolE/RpUvzql7+K9dU1JQoUU+gJiw6W2vkc2mX6pFCaqG0lrBxUHAok7wRlJVlOaCSPlGZGFHs0f2/duaMJ5+OnT3OKbYSO0ZtpdJSPnKBKkk6CzmcGRSc2xqK1LdU4AckJAkVGTx5EkJyVV4Om2KXJ6I5i60DmZ0HUCKkiVILvuQqTEyNFJWWVyXIZLBkl4Yk/36/mb14DQ4ZicZTXiBolhUDsYENwj3hepg4ycfY9VLOO5CITEbEFslln3U/LBqkpifYl8jCJapCJIyTYNN5SEnHqZjEHj/w2RBc3ZZRioJqShRbSoEcSXm15laIoM/0G9Q7FGyTuypsVFRo0K8moeLY1AKmGvhKgjuqphhWFUKfJ03moV4JSybR/LXmTzp/2sdyJUpFOfw4tuK/FOKEoIpFmrWgd6ZCC3QPq90wa7Bvrm6IDknhSmCrxy6Sc9cHzLt3jQg5pWOAPl0lusj5oWKGh0Fk1Kv/x91GgyMuFZ54N1LoHlbRxXawvCi0349rNXaESUt5MyVp2bJW02KjC7eWi2SZzAL8H06Gtfc4wkqElwz+YDBubG2IUffvwWw22yuBbSMU0KCMJ0X5JdElbJxXd62GzUwYGpfsrTWhpZaafB3TMYRuUc89Hx8bioqc3RkbH1OyZnpoR4uqzz36tQswNgT4hro02QzvYqKC87do75SlQUlgacqXGpJhd2Ux2Ctrxlc1ONRhTs5nPr0Z5ZqatgUQmhWq6lWZEvpiS0Lca79WI/z5jor0GnKQWyqYeWRupz9CpKM5OsmzQWDqsjqlHv0M5LllBEKhIa4H+57VgjPFxjw8PtTaEHNO6SHQdTVCtxTYq00NGFws0Xkhya+0b/YlBuuULFAdTPq6Kcy95o/C1H4WgyrMiqdl+IrmXi1FW5oLJRLM/TrKFaFTIy8l7gKXuIsAeHVwvzUM1uFNCguYcBT1fFJiSzys9YDUcibH+XNqjWmVIGFqKkXuleC8Gkoc4QmqnrFm9v5dM5zi21poHIG8PG35sQPFDWc+PDSrqHv/nZEr6iPKXGRHqiIKFGM55d3hohCP3XH5GnLP4zuCzJe1mwBRGW0v2KGWgXGSHvFBs3twu9gBkkFOAXEUPuvxWJLmCYXQWrPJ0SCPQGsSpSE65DN6Tew+jogrrtwcV/Lsbb+3BsRC8vb3KJ9A2J54IGJAIQlCbpyfNePj4kZF22ewRMi2N1csDpu0h5nXbZo2ZAdnX4xzu4sIIfuLA2elF9Pf0x/lpnu8wXBem4/692/H69WudOzdv34n/5c//1+hL6acrl6/EG2Rl0nRezfuBvujp74u+9KsZR6qzcSJZNprLPAA+L8withBSm2oSijV0qlyKYcbE+Kjiq+XeTpV30oySJ4GMQsmpQIn2q1BE1ksSKtJCx2/iTPcSBLoapngIHDVjiCbw/m589fChEOictx5U2MiTeNPF58z115XMxu+dUynhUkMkDetoNgj4g4nzpAYV1Qjr3G4+bqupYFaE47D/3qAWIzl5nkZL04RzTMTkWmzbbg/R2PdoKyPtQwQSA/YI2TCjjjXA03WFCmSjBx3OSgqRPLp50tC+WH/zJhbnpuPstBHN86ZYFXx7o3Eeb1bWI7oHBfxAomt8jL05FKfNRgz2dMX89FR0wegYH5VZ+nlPX7xYXYu5hUUV3Bura/HBO+/ExcVJnJw14vyiO/CRPTg+FVr/XCxUYqdzzvHRcdUlYnlnc1W5IbIQ/QNGIMNKPm6oYUhTAWQ+TTAGA1wP+SjrlwYkPng0pt+5fy9+/evP49Ligs13H38X7713T+f6+tpqvHP7egzT9D63sW+38lma4AC8TnQP8dfo7h+IL7/+Jg4bXI/3JPdauRveVgODikmYMPNvvH5fyqCyXmhKqBkjCVjTCsntxsbGHTs4lwaQI9oTkEUN8j30rw2soKG6eMk+CZsbmzE6PiIQBzn7wuK8/Fd4bQ0Izs8EAnqzuhYLM9Nx796dePPypZhIrLOXK6/E7MDnA5YGw0xqru2dvfj0009j6eXz2DnYj+0d6kSjuNUoPD8Xs4Hr4T6zF2BHMaBkLTO8IX9jmCT/pwRUWTbxPBYW5pU3gVgt4BanG7GeMx2TcYbB1ILV4JbcD4blDCJPML1vSq6MGCIQDHJrALhY43GuZtXk+EhMz05pmMFg4hn2xfMAACAASURBVNHj52LJ8Nr8gKR9B6izBnXWcHYCriNuCUmcZt3I/uIHMzbqus/eIPZEIv5I0iMbhVUrmb0wpmempmx067ySvFsCEHTen5/o3GftwLhA0pQ8GFlTPh8NOTUNK6+FQZ4seO5NnUNEksqxVNtlblvnELG/zscaVBQIrQZQvAbXBEuGHM7AMPcIqlFIrcF7AgYQAK1ktGCyiA3iZhxxhu8T8K7R0BCjPahgsGuAkepZneuuD8X6gymYoAT2kPLrHktDsw6QlLZ0kesKzn+uibXnc/4w7ty+pbW3vc068qCG7+UssYIB4JiGcrYPPvhAgMbV1TfaB+T8DOTHR8dkns4AVQbss7PxxW++1JD43ffejV/+6pdas7fu3IrV9TWd1VMTUzE55kHF4sKlODhuxBH1tHoUFwJKsjYMjgnFWq4VryPO/+mpqXjw4IGu+euvv5H/ltZan9me/J77LrWHLvtuUDMRY/h78l/3EwqsUqbMoMAbekb2wwGkBbL9++AiMWokq2cvnZafQZ6JOsWykV25Tg3PJFmUUmgGGXod8ux4pm5Qt9H4+nMC/yqPrAa2Bn8p0eta0gcYv/fAxaxR9Sg69oE9n/zl3NYMsMq7tI/4M7l01vDtfNc1fYH0HJsqd/Zwoz5nxbQCIxSAyMOvYn/YRLxev934N7un6pgCefneFFDB+Tr3wwATX0+9VtWZ6mVV3afvavvptb+/fR2qgbL3Uyxry0+2pa9KKUODq+wz+Vmngbm+v2PQk8MM5d7y7zPqvyQaWyoVHQCeKpSJE5YSNtiLM72UR6gDuJ7Km+1r0hsX+MuMj8X+Pozn07hoHsdw70WM90f8i3/yxzEy0C9G6JNnLyP6huLl+m6cd/fH4NCw6n+uiwFs+c8xhOezGiRpLwv2OPeVuMJ7EteI/+plpQ+m17RjCzGO2oyzFF9avdaZGWzEUvJasYP7+vTaAGOQqWQvFeOS9yIPYJ/yTMyQc1ysHLFku37yqPjPqSx/+t7fizswn40rNiMbgY0jU7j8exnDyHyoK/A6OCMJzOlrBTMf9nUIouVpap/pdsQwe1QEGuS9RnFQbEEb50BV4076owPxB3/4qRrX6AVDb0L+hgSe7ydgkuD9xX/8Cw9T0nhtcIDiiGbugAJAHXxGE9Lgto6fi0cKXcRabZolSivFoA45S7W48T0Q16/d0Ht/8/BhNDTBN5VUkkKZELqp5eEAVGYGJyBpCCxF+6coIrnggK8kW8dGK4i3zYo7p9g1tKhOJUmiZbj8syq4U7bJaP4ydkq91JSL4jr5fKXtWPRIH3CmESqhkeG4ByiSnsrpdX0PgZQfqGluITYLLcB6oEnd1v+k2TieU2+bkWpCn80WPhfoVQ2O8nDj+j28Ac15qrXG2uTwGBlyo1NDj/we1hiBv/R/OUxA9/E6UGNBwIGso6Al6ZXUVHe3kmTWFwUdes32McFs1RP7atLpnrYMqArd0SmbkthyQzD1JYSEGi1t7Uj9fcpz1YFSclidyYQS+ZbOpuVv+Lx8boZ3pWfshooHAaz36WnMwg815ecaKLIY9nBfGZKJHlmJ4A/4VFhqpm2Y/b1mdUoz+eoKlWGkmwzoe/taA4KSgLKniL1falDWRtcUVb0t/aRmKwl0h44/zVqGFFwPTR9QRzBFbt28KS1m1u3z5WVpTq6urcfe3m6LEQH6wMlcl9C83GNrtbrYaTWf0/CPgSLSUW2KvB9oJZncS5B1NJ7Gp6ZkpknRSuEC8vLZkyet/cfeZNBUeqiOK3gStGnDQuaoodiWgKq1XwhCJZ45mKjhUDW3Wwl2Nq1bTeFkQ+hnO2ZklnpzPORzqDDORKsGG1XA1mAxM2An7SnnxXlgBBPMJ7NVasjkgYDXR6G7K4mW/nKi4Rz72trJuhfEFgoQ7hvPvNkUEpPPhgQHAVsJvBC2fGuPktLu7pRq6fHwwvvPRQPNKz6HinQGLEmhVQ8yhxGFQPRnarPQOpvJek6JUizUaLvAKF3Z9s/6dfwe1SSuvdCidZc/TZqgJSNbyM+K+/UeKjzTc6JlCM4bcB9Sd9/P1kZu0IQ1lJHkFAWgyoRWMaMhV4ccYhUtnYOJGrS+XXz92KDih4YSlQB9v4hqD0X+rp/53eTpQoXrwsKcdcq3d3Te01xmCKCCJ4sk3XeaKkKNn7bOK9Y7RTtff/RHfyQ5lYcPvxXCWoPyHiP9ud/cN5BVFLoMszn7+aKROShvqjPFApmU571kbdikkmGbfW6Iu8SbGlTUunNM7BGiCrRrsTH5e8ta+N8x6eN1aJZoTYN6bZzEgw8/VK7xV3/z14r1Jzm4kfRm6nSXxEitbf6Ns5CGptFZNjLtVV5D4w/2Jpq/nF0I2jjvY4JAfnZpYTYmJjAZPVJD9eNPP42//fyzZKBgDNtUQ4bCi+9BxmV8asKgiNxDsFFYjmoegSzDhHzQlHrOa5ovfD/5EtJtz58vaeDIa/G6BsbY+0Ea8tmsI6/jvtBAU8yh4YPpMQax2QSRdMDefkteo+u8O/qHB2N9azMePnmiRrdYmKXzLBU6Vcl58tnsvtCKtYeETsxGK+vCGtxqe2iMyvnIOcZnFbsv14aZWI7/xZCwsTlxLYevYv3pirzGJQ3nRpz2sZgSjqfkWhS8+HHx2WAYjI3jJQHaGc8Re5ARO8mnOAvFrEk5RcnmIWdwYjNb9lfjaD/Gh0F6Y2R5HBfdHppMT8/F5uYu0TaePbPUzscffxgba6uxv7cTVy8taEjRByMGSQjAOGfn8WJ1PRavXI31tc14/eJVXF1Ep3kiEFHq6uqNo8ZZrK5vR/M8Ymp2RuthZ3dbn+ny4uVYXV1vmYdeWrwUr1+/knQjzxbENM8BMMtA6luDiNcAbKAvVt6sxv17d8TQhsF9/eo1Nfzu3L2rYTjs2jt3bitfAum7uDgr2aMrizMx2NcTp40jGbADluC+wUShLumSzBbOH12xd9iIx8+W4oSGhfma+q/qCjXQVMeMCnHNXmSv+9wD4ICBs2UuaDQCYCq0O/mLvfUulBcCHqFZTDyUpJ0a/QsaVNDomJ2Z1qCCNTe/AEP3RKxb9gnDqNFhTHWPVP988vFH8cu/+WWMj4+J1dFonojZsb27H5cXFmJ+bja2N7flEfLBgw/jzfqqWOYHRw3dk4rlxJ733n03GifH9g8BTFEyqcSvwUEBTAAMSZIw9edrg9kbCv+OXa0pgwmYCdF4N0CL+1UDAIGWYGHBrAFwMjQsPx1J3zJwBdUMG1s6aacx3NsT1y4vxvgo5qZj0TfYH/tHh7G8vBpd3X2SlWIARe4Gc7mYDsRKWDHUJNRhB8cHyqNgBrAPuaesn5J7NOofRgEMWuevQpNrTx2pMQZ7n73O55ckDUMdgFyJ+oZlRCOXvyOX4Ys6d30TxshZ7MHgSMa8m7Ae2Bj17QF9/b4GFXX2c6/qXgqImIOB+j7nzgaX1ff6GVnah1+rmV+sEQ/XDBJR80wm4pb+QipQQ0ea8Ko5nYNKBlha8/ZF9DPvAMClbDH5uyR5Mt9UfNNA4dgyg8nW1truH4jBgWFdH3vBZ8K5hno8L3KGhfk5DT1hKxjFfqaBkNHsXrMAID795FP5QzBUZIhHXkTfYWxkRAM53h/1B3yIfvPb3+q+f/DB+/G3v/xlDI+OxI2bN+LJ0yd6LmJgj47Ht18/jLn5BXkDvXy9EjsMfABPJFOE56hBzuio64/AbBqQIMPjScmfPX321B5ZmTuzr4nrMjpWTeP0n2uampg0o4Y+iPwm2F/J0EkzdXIj7ilnF/tF+Udvrz0dpZLh/LZyYeV0An7k+VWNfzXDy3upXYBUvq/BErVDXk9JwXU2t1k3kkRLFmPlpZXfyoMUD59B+6Iou9V5mJ445bVG/KW3kL4UxMsa+BbosMBaVRs5v/3hHLWk5tp5bet3beBRh0yZBxv+fNr7Anpyn2GMmNnQucd87nMee4BRIAbVIgI+mWFddA7ytHbunlLdem7OPasWU/aQPSPdS0li+TNUPVJ1jdk11Es5bOhgkihHbtUNPKO2Z55ziPJWNIir8s56PuTK9fM1YKna0qywlOZNQC/fq3PupKkaEHaxBglHmc/ImxXvCnJsg164Jpi+gFcEENlYjaHu05gc6o5/+o/+YYyg1LG3H4+ePI/RqYV49HwlXq1vi41H7GffS0opQULks+RKGpT0DcijaWhkpCXxynuWCbj2DL2axnFKU7kWIKfm883PzcWjR4+V8wtsOjGhffDs2ZJ83cjf6EsBGOX8pe6wGkSP9p3OnfRM9P1re6SqDkyW9E+Dit+tHn/6m9/zOzDFIX16pmJdNENoU719Spz5s7T+SSSQe5LkiOnoCmyJ/K+BgBgWSTk3vQxEqvLDGBwiyW5oQODmeiMG+4djsA+WANP8rnjn/p24fedW7B1STFpGYXZ+TocviT2bdG5+Pv71//6v1Xg2mshmWxSvIIuqoaREq5p1GIJLF5RD1Ihagr4Q9A0a111x3jy1Rid6csOj8gEAaUMQwagNbeBCcTmo+yAvcC3BvxAloKa40NaBoUIJCivJramWNY3/fkOoTR90cG+b+VaThF+RKpKGH4U1jbgT6LiNNF32AcG/1ZeblknRy4O4KMA23faAQbJU2RSncetpdYHs/bo2NnNiV/qUouGmPh6DnUqGWUNuljvxZG0Ucti0UxsflXSQP6Ob/FX882eKNp4XCEAaN/ysElAVjEiGHalIIDmWkVoimTjUj45BHjqhItBL03BgUMksxZI1YZ3wQkvu1HItX4bOLd5KlAtlncjlOmTZHzQiyo+iELxmsLjRoNdIWGUNl6wdadN3SQukZBENH2QKOCBBa/GFPImMky58UIHmoWhhr4IElibs4EBLAokktdgMnYlaZxPSAzIzb/hoJMFKdoSWM5qJNcMwq6idRogYlatYgASDEBMeRFQjvBIWNfDSAFjNmUQ000lwEiYhcA1qRPtvyYJ5L3D/7t29Fzdv3lTSApIJzdatnS0hpNivpEig8lRg0bBT0uZCyNqlRmioGSx0ofXWAZ5gzEojU1qjma4KDXnSiPm5+ZTaOI2FS5clS2JpoYP4xV/+pWIdCRSF11kOE400yyGhmsZORMU2o+neYZpdbAUnohbrsYZ8GjZ0gN7tw9DmWbRi3ts+FEn7LbZFaYhK+zyTfZ6hWWRJ7U26rzSak53Qlhyx/I32SA7eiDs8c5pnlijDZBgJLYbBfl0hl4QeNMqEfcv31Odu7wGfKTTYuPaRQWQJuyU58c69ezozQIAeN6xNL28L2kPdDEFIsM3mYVCuIiCL6mJ30UTRvch4JLkZ3Uc337wvjVSq2y0UkOTHvGercC/GYDuOZzuxxYTxddvLxwk4a1hN9DTEa9GzWXym/UX3RRr4IrmYz6nYNaCgW4MqrQsPkIoxCJuCZ2GUuZsJrB8VNLmXW8PqjqFMraW6Nv5cRVBnjOgcOLyd9vx9hw6dg46/78/4vVwYz83M2OQOhkJXV0qvnaqRAJKTPUec1NAMrXjOYs6e1HHnjrFv/+xf/ln85V/8XPGD6wa1yK5TU6C/X0hs1i86/gxFZKCYKDYkHHh/oW4Zfp4yVBtrSTy1ytdEhPJMaFL7vlqWQJIMERo+E58rd+DvhbjKtUIctyxAt+Iia4eYMzs9I2Tyz3/xl47tfPaURyuwBsUaS6uGiZJWVG7n/St5FJmt+yzXwJzGMvJPp0hCWVKIs5EhxuX5uRge6dfAmHU/NjkZI+PjsQuNnSEA+U0Tk/KGBuqXLi8qdjLSZo1SdKL5uzg/L2Rrf5/NCYnNSGzu7u9pf5p9xCM/E0pZnl7J7hkbGdX6BrBCTkUzl/yRtU9Tgkao5HEaINDGdK8oNlkX8rA6sLav7tnpRQwOD8XG9lZ88/i7GBxmiANrzzKBrBViNLEYdJ6K0jS/bKMP3ZwzAg+Gq8/Jimka5jebyq/Jp5S7ALbItWTJBksseEBp1KP/3kCEGnArRuN+7V2fRf95DHHm0KzvH3SMiq6YmpoUO4ac+OBwrzXw55nt7R8ZyScmMZJZDBxKssFxiHsMSnCYZtBpQwj0sYnRePVqWajCyYkp+Wn85jcP4/7de5a26kXTGSmgZowODcTU6EjMjI/F+uqbuHz5amwfHcXS6zdx9cbNeP7seRyRz/X1xc2bV+K8i4ZXd7x6sxEra1vROD2T7vvm9lbs7m0rti/MLSjPIxYzJLx953Y8f/ZM65UGG2uQvInm/NjYhPJ5GvYbm9tx+dJiPF1aiqmpcXl5IR+0uLCovYVPw/179yQLxb4m3+I1YIbMzU7EQF9PdCNRQsMrdcLVyDxAkqJH0i0axLEO+gfiyfJyLK9sahhyzvM4ByRh+U7ikJoyvT1qRCK1xDMTIEPs7obyVJgUnJOcl9bivlBjA0lZ1jfNfvaGDIZHQLkfa90yvOG5rr5Z1TkKS1EeOhNjGioRJ2EWw7jB74NrGx0eio8efBif/epXyu1hgM/Mz0si6umzF9Hb1RXXrlyKibFxfT4ktFbW1+KLr7/ROi07NwZbxF3MybmXMF0rt6hGJ41Pajr0vCsGsv7LY0DD1JTLk78XuUUfMsKDem/qFeJVyXM6z7QcTwF6GHIIwQ/LKmUfx0dGYgy/la7IQcVITEzZrB094r/92y+jf2BI7BgGpiB2Wed6r8FB5SvsL+I0e3z/6ECG46wBYhwxCqYL8ZTv4XmQl7O/eF4MVqt2EEuh2xI0G+vrkg+mblJOjIdf/6Ak1mg+iyHXZfAfNS/XyL0jjjDk5f+qZzVcpFYqzxx5NLj5b8ZcG2hVA4k6j9j/JXWqXDvzvGKd8kw0EEsgGuvSctHZ2NTgwMMRYhZfGoKn/wTxiS9Ag0SoqhvIG6lVO/M3ARO7e2JAgzxLOtWZRUO/2CrcF+pB9ir7ivrHHj6uPyyzkrmV5KHsWTQwYFkg1Bmmp2fi1auXqiHpX/BsODsKPPbHf/zH8pY8PNxXM5PIu/T0Wdy4cV1SgvhE3bp9K0bHRrXmN7c2tf4//+ILrdFrN67H4+++08B8bmY2hvoHJREz2D8kD6bHT58lgOZCEtjsJ8B7DBEB6pDPcm52KlYQ13a2dwymC/sW2g/TUpi6P3nmUQsiS815DDtULCQxQl0DcM2u/dpAFmVbWQC54d1WgmAdulaAxYgktZvPxUhxH/37wwqfa9WwZx0mmChH+c6rqC3sxSk2TPpfJAxQ96UAkBr6nthfrNZ0K3/PuskSmP5p4rL2RV5jNcnrjFaezNmd675NYe8out5OeDt47tXvqH3TCTSqAYoADOqleYjoa2wPKvjZYon5WdS/tVnTVgto7y/XsH4+UpzQGdJmQAjLlKAkAaayxlMNkhKarf5O1uPtIZMHEQYyOMephrxiVA4Ya9DB5zWLpbwrSlXCi4n/BIZBtSEHS1V/6VknG6bikXo7rIkuN/6pw3l/8kcGj+xt4ixxjTzP8eqkJT0MyAjARuNwJ/rOmzExcBH/4p/8ic7wtbWt+ObhkxiemI8nr1bj9eZu3Lp5K168fqn8mPvGva46VRKoZwZdI/NELgc4kn20tr4e169fV/+NPIIYSQ+VISaMLYAHxMyZ6SkBl5eXn+usIK6hCiHQnO6v62OeI+ofoE8AISh/REkiwVHsW3IJxVg932QEZV9VNVrv4j9sdwd+Z+H+9Bc/3YHfvzswp8BmjUglPalrLMqcEg+jzKvwB+HBJijJIfkTZOPViAdoSW5yEgwpZs6aGMshMYXWGwZpZ0KnqDnLfjvjz4Px6c8+0uGjqb8kn85lijmASXVvryR8fvv1b+Prr35rjcVE2JCM8xmruahmYBp7c6gVLZLJJM1P6Px8RkspHUtbF61XgsDw4JBkXWhcPHm2JOMdgn8vSJ4TI7P5kpG3NFeNoiTAliQTVFYlvDL9Aq3JTyQiQeapRUFsSwTV9LyaGZXYFyVStMc0LAIFRVIGIqsO6DJ1I3pVstIKYinNRECspFs+Fzk4oJDmwHOThAagp9QUs5XQGA3jwQONdF7b8lBovlsCzO0kN2GVcKXxMs+ORNKUNyNs1LTMQQzNAFOg26hmDRtS/5T3LQR4vYcMLjOjqgOSg0XoHoI8PhQK4j4g66tkATSU29n1wApZikSbO2kyq+OHviqh4/O0fkYNRJswu+FsKiSNC5maZiM4IRJ5/ZYiakn+5ACjkLTSW8yhgA+66Rbd2kgbtLv7VMRSECFTxoHOtH58ckIaia9fvZR3A/dSSA7WfTJGnFxaq1KJpYZvRgKbmuuvug98n2Wa6mfadE8PuDo1cv2aWsti55jJpESxpDNaWpWWdGndo7r/JNOSXwH16UQaRNJHH31k/47jY2m/UqSQjMuAkhhwjkQEOtpGIYlimuaxNsUy2prPh0knjUKZreH1gplWUsFpeHWifNDG53poDo6OT6o5ybP9/NefiYmhxi7SHBRLxLkuo8o0nEmkiZN6Dypqn+cS9t4pEzoZH7fZHG1Gj5OTSuz0+RK8IomDt56Zk6BKZCw9xdpkbRk5Y0RtPeei4+rPyVqqJmcN2qpwETuJwo9iMFGsouWrqPEg0U1/D+cqiedXM1tc5HC+1JDGN4H4AYKwT3IRxJg//Nmn8d57H8TX33wTL1+txMbWjuKyUEFCX0N3bxuTFiunrQNvxhxxTms72U5ao631n14auf7qOjnPpBNfhncZJ3xdxZhqa62WbAv7Ws8kjao9dE7GRxaLNRihzaxYwpkpQ3JLhjTRnwdBLrZTMo60APh+m11oGJ8uiUZbm6UjUzjQWekTYh3sGhYVYsufp7OBYUo+A7U2q6zWx3/poOLtmPqfO6gY6OtVgxomE+cwBToJPGc1TSKZNSZ63uvawx6fGbB8mpYVHBzSOedi3wUhRQTFF99J02wjY4oMOpvNaDTc1Bc9e3DQsiV5TtBYYXAqWRUZqBtBxx4R0y9CwxPep+I7v2cPlEeFmu2YAEr/3qhh1gFNSKG8GseOkzJ67lEMfOedd+IXf/ULNb5pfFragWa2UVgyfiyz1TI4zBhQMmA6f8RxcDGJ+y/PiYYPDbQLTAk18DiPK5cXY2piRJ5YNCxglR0CdFBx50HzaaMZh3v7QsHfvHVLz2lgaFDNcEl2AXY5NXW9mIM8IxpOQgV32Y8BpgB6wwxxFK8DiZGUhZK8nr1J1HQgvlDonsOeAnRjuRYKTKHZut0w45kf7tuzRs/i5CwGhkFHH8Vvvv5a95oGD/dX7APtRZuSUzgqXuWQu+J3xWI3H+zD5M/rNcdn5M9mUfoe8x4thEsH28RNXw8qKmeh2e08i2FIyuhJHiqD/cV5DA+BLHXRikcBr68ziPxbeQxR4Dz2dg+V+9qHxA0TfrBQlKWbXw1HDXxPm4Fc197OViwszsbK6xdqNIP+6+nqj4ffPo6FhUWBSMjx8YzY2d6UGffc5ERMjgzHqxcvYnZhIS56++Llm/VYuHw1Xr9eib3tbXkezM6MR/RcxMjYRGzvHsXTpVeYosXC5UtCu+8fwJDtkvTT5uZ2S797emY63qysRtfFmRoIE+nhtra6FuOTk2r40tiGVQGas2SDaCaw754/fxHXr11RHNnY2Ip337kfS8+X5d3A0fryxYu4dnU+Zqcn44D1O9gffb1dakLbYJlnXewWmrDd0XTiEY+XlmJzG98NmkkXihkalAOYGRzSdckzZ2RYa5HXVAOJYWIfPmX2JGOw4LOS5tCgvAtAQ9PE1HAQptX5eQv5jIQlawypIJ45e0tNJdVDRoPrjAZYlJ4GM5MTcf36tfjqiy8EgiKPunTlckxMTWowtL66Gn1dIMKn9LrkM5u727H8+pWaJix0D9ucIyJRI7Q7SNSeHmt1Z+zkGvGgIaawTw1yMDhEvhodciXEwJKZoQnLnpyY5DNttQy6y/uGDXf1Cn4nGKKvq9krOVoNX7tieKA/hmm29/XG1cUFMa1nZiejqxeT0uH4xd98Fs3Tc8lyHR+fCKVPHKCmsA/eWfT19On+ab9cnClm0azni31HTSWU9zkehZYQ5b5QrxUog4GKAT7W6kdKlAZ6na3Kw1MS5sJ9SX0fDTtQxcQR1iv3htpYzLSU6+k8p/mM8m9K1HEngK+GENVQZR3xd2WAXY1cf06fezIM1/OkcegBvV/T+QMAFTH8E7znuoJcEHBTr/YA9QnxiAE1Z7Ebi5bJkrRXemMpT8uzElAJ7B/uJ4M3M4nMmlDNr1zIEjc+N3pSyx4JlxMx8eyLhmzksD7n8dFhTE9bVhfQE58VGTgGepz3nG8MwckpPvn0E0mY8bww3GXAt7W5qTXOMPjZs6diITE05XoPjg4Fnvzl3/4yJqYmdE4/fvJEOcXs1IxQ2etv1mNickrgsqfPnytmEJNr+F0DI6RP9axUL7tvIJAjDB6knNSMnTBjHtP1lI8hnsi3sa9PDELumZi1nAew+vV7N3YLoFR5us811x/c09rDtZZ4LvydAHfJpjD4q3KtHC0kwK3FpkoJTIMJfY7pc/Q6J6rmuYYVNWCgXkxp69rHnMncK4Nbaew6H7L8mRn6nJ3OR6yGAIhDeyPY62ZhsHaLwVDsfw3DdP0G69V+KoZF5ftZpuQBbDBBDWtqmGDWuWsuft7PDhkyapD2+e0emVlLfCa/v2uyqsMrNzRLqvJ1945qCKS4Sh8sJcDqszrHtqRTfZU8r4BR+Vk6n4EBGqlCkiAz13W8PgMV6kcDFkt2SwOYDsUIvl++lJl3ekDGgN59BzN77KMlqbPsR2gwneuJ6yXuFeBR9TRrPGXoK5dSfpUqLwJ4pEffKeDdvoje00a8c3MhPn7vXpw3T2J7+yCWX63H0PhMLK9tx95RM/oGrbahWjtrVuILZy3ApRKzAuTAHwBAGHgH83JRvYTqszCwx0z79cqK1unQMB6XPZZ9z1hEPGSQIilk+hunZ8pVkPtmwE9vg5grzhyQdAAAIABJREFUsCXXnXvfYE/3znRWAktpMeYTwvLToKK11n/6zX8jd2AmzcoIWtLAHxpyQVzyHKC2MwFVyZPGLdV4bzeD2pNwNQgz6GoaieBsFwkFB6Slkghyc3MLokXLYLEnRMum+Q6VmiY3WsMEKQISwwOQJH/1C4zxzpU0FoKHIr0tR+UGXyFB7LFhFgOJEMke0hjsbjY6aCyua2trQ4UMRjlQfh8+eqxEB+RW0eLqmoWIUuBv0/qqQc6hsyvasg2SlLyntqCKGzVOEjGXND4fJm4oOrB/n1lRxU2hUHg97rs9A3zIQWGlAOLPFD+FYCCoW8rL98RoB9MLi3YntHlPjxJgiiSjLKFJdhhFSV/SshRG+fjwJYDynj5crIWvA6wDja/PygHE5y0aY1baBNlWklTBtzwesrDr1JG05iwyLi7qfC+M6CiEft1HN0TRrrZupZKu1HxVA1FI47bsgr6vY0hRjbVqqFVj0w14D/eq2cjza9PYnRSURFglC9w3T8ZpELu5U2uoGtBqYIn+nWakOTjkPpHsGsHkgRq/p7ig0KGxzrq5dPlSzMzOCo0Fusf6qqutgYMaKpmoVpJaTReGOjXsczLWNnymMOCrtPa9jjy09OFZxmY2DlNDPJOzQp3LdCwbLNXgqYaLD12QPpZo873PQUcmQXdu35a2NIgGJK6++OKL2NnbFb2c75dsCMO4AYynbGLL/6Bkq3NE0mFt0FDRgmYyaFn2klCJoPkYLCTdWkXo7KzYW2jUUij39g4IqUqBwKDCiCQKWSfsyBZVEqMEHFmSUxdlNegsTdOiu+tZpH6pUO+a4DoR1XpW0mefFrOZvA8qTgsB/EPDtWQIeHBrpFwNpiiARCsWwsa0cb1G6p1WL8zoX6/1ioUlF0JRybWC2pLmMJ4qzVOhy0A6GvPvRiIyELymvRpMXa09xQMBbAPSmqE1exGTz/ffeyc+fvAgvnvyJJro5ff2xdNnz6Nxchr7B4dGJ6dOZ8n71b3iXGkl58rqM8nPQUU1ccsAvPZ5oUC9/tPTp9gtiQbqHGa6FnHs1vMUMej7sdyFSCEaSxoq76sftNYuI4+KI2qOsN953iX90irIjP5nTeksyvhHEqthcYfpttdaFUHpjfHWvalGSWlB/38xqPgvS5lAs3fJbNVDaAx0C5lmFJfWVRZGXA/DRHKDQmASF0oGqFhWZhWYiTI5NSEwgsZAFyHDbNYtTa+ThgcesDHo+BFzS8ecNUxM4nl1ouuUX2RDx9rlbXnGGlTILLvZVByvz6m9mIUJSE3QWhQ0xCb8HZBPojhCI/vXn30Wa5sbMTA0oIGK44j3qZkV6RWUsGdih1mEZgsYVGC93T6Z7nqtnZ4SayxbIpnE/b24dvVSzM1NxfKzZ0J8joxP4I4tfX5eg/jXODyOg509NecuX7mse2lvsGxIZIHKIJdnRNOJ5b+wuBBr62tqFhW4gyOFRqlRdgAzhvQ8KNJmpmZ0rZiLugGRbE1pZ8OAsvQTwAoZ019cxNTEROzs7Lak4DTU6u2Nw8ZRfPv4iQYBYgRyr2CUpEcM+0+m4BWvsqlgDWgX3jVMZo1UPHH+5yOPdUFDyxJgzr/eHuA69NK4aKMmuQfVZNTwiXxHw103o2CdMFzC1Lc8vchhkS3RQEKAGprfXXpmNFZpOglAkShMsYzVGLRpo5o+yqt6BATgvcSc6wf53h/bWxsxNTkd/X1DcXSIKbSHfiCVkWs8OTmK8eGhGOztVmOYfYsvwnlPf7xe34xrt27H3s5eNI8bcev69TjY34mzLhCtXbG+tRfLr1bFbbp7/37sHuzJHJ11Mjc7J0CGdb4tu8O92dnasucJ7Bw8KtRQRe95JFbXkPTpFgiBvBi5HZoKd+/dlawT95Cm/8uXrySbxFpbXn4RDz54N1bwsDg8iPfeuxPN46NgUMoJJvmazLsxcpZ3EveSnIcmIoac0R0Pnz43WEdgLwMkDNLps/dJMsJATtKkYPjDcyGusN9pVPAciQUlrQuzlrhPw8uSEDRmh9ToHcrGNK/Lz4DmJAayN6hljHq2DCLPG+YTP3/96lUNIXd3tuPVy9exvr0T4+OjMTk9pUHr6spK7GxtK+7wvXMLC/F67U3sHh5Y+ooaDgZmfhZiGWvMDVM3oiqmEQuspW+/ggJt8cyIyaDcqUOLgWZJIJ+bDAEWFxZkZOqfc47o4fx5XL1yRQMzpJHMLisGZVdMjIwErAq8U5AlG+zrjamZyehGivjiIn7+i89icmZOr0feghQd+SQxhDOdNU4EEMtXKG0jsN1AdhOY+8t57X2f3j4amAMOMVqePUYco64sMBIBgrVhhp7vm+K35GEA37DneX0Glh6Gsy6ovYo9WU1N7nflvc5fXIvVwEHxKZ9L1en8Hb+vprTzWa9p156Dzu0wds37ToyqPJprlSRZq2/gfIjrNYM2z2nuV7KfWC8MYIhVVReSUxOvWTul8MBQkYEB+fxnn30m1HIh6YX4JlZKW596PlHQ/L1yHn8GA+/w9vG64zm2QUyW+eIsffbsmYZlklHKmAcYgKEqZ+vipUV5UvB5Li3Ma9CHXAyxh0Hp+saaDK8Zrn/79bc6q67fvB6//vwzxa7piakYGRyOh18/jCtXr8b+0bE8Kg4ZsHCOal9+32uh8kzyFNYJZxFSa6x9mI4aah4yfGco2Za91iAeg2oNQfrFTuF7WHeux82UlI9ZGhgrjUwjZte4bqI7/rg24JkRm8i15DvaIdWrPpF2R3mbuZle7L9SPGAPqJHPcFNyw/V9yeTIOkPXLtBH5tXKkc2OBWCqugLAavoxVpyonovTcvcKrK7huFfXolyiZc5sMJOQ/4lrLGDXD5VVbaBAJ9O6AHpl8O062PfQ4LCKhR4G2reHf696u2rldk1uUGxJZPn7SuLVf3DfoxgVjq9+pgY9aajU4WFRPgqu4dsSvI4DdUZZcq8lCc7gt75X7AnnIFKMSGBODXwqxpjJXR4iDgn8b5k2D2ANICrWugc+1b+RF0R6vVZ805pO7xTl+DoHzU7zgMdrnOdIPtvf1Yzm/kH80Ue348blOXkAbmzuxtKL1RgYmY7XW/vRMzgSh+p9DsrI+uQkATBdofxGzyIlPPE8ZV/Q46P2JGaRw3NGyA+RWJNS5PQa9cwl+2VgqvKxvEaun3yAn+NecS0MPxlAr2+uRW8PuYVzV3vS+ufLm6QTEEMroEBaPzEq/ssqzZ9++v+Hd2DmFAqfUcucMjIKTukXHzFpKpgdTEtJ+F8cHI3cUILXwJ/AOoA+wJhqu7jCZA9TP4odUDs/+/Rnsbd7EKMEI6Fij+Py4lzMz8/FyQlN9B5NTmFWgFyBfvk3f/O3OqyFBDu/kBmcEtyui+gRaiP1pU9PRW8WhR29OhXwbZ1hPpqpd2jsG+3C57u8eElBBjkIjHUo/ggyaj7kYIPA7GTbDXnQInWo8CufzYMKU+0IwjIEk5GwpXRqQl+HeB3sxapwY8mJou5lshbqMONXmy1PtNBYNPhIzi2VhOyPfR8oYKT3mAfczs62UDwkiGVIJVQOkkPNE1GopXlNQ0R68GZNFAKQqXoV521TH39ONevTaJqkuwp71gwNek29tb4K3W3UhmWPjNbnc0hvUP4HND392ZSEkMBAbwTBI0RaDqjSyKrkvzpRSU5onLCTZDPcAq1mxIEbSSBxKmnXdSRDqNVETYR5NZqcICUTIZHVpcla5ld1kNd94fPTJJD5ezY2qoiohEqJqD4j0h8gPs5S4soHGqgZ6bTPzcX62poQhgwlKOxgFFCM00in+c5rc+0klewLhn4MLWo4ZTS6tWLbTcpsTbcSfz+f0jxVwpqNW+69Bg9ZLJI8yuSstf/PVXgV/ZpDWs2wepaF5DYwPPeG730NHVXoyNfkVEPEBx8+UKOQz/vNt9/E6tqa0A78Dw0fJAKmrVD/hW5oNGJ6ZialW6zdOzRkjXWvUzdQBoYttcK6BsXIZ4Cl1Ww09Wfi0OqbN0Iws5cHB0fU/PrFL36hv2ddgKZUUpYJHc+pZVbdjW6maee1dgr5Xo1N308nWMU2KlhP0Ty1TjLRLlk7FcT6+3ZTPmsFv1eiNPWcae5C3faCU1ysQYV8IWha1qAiB2Q1WSpEepmP14CS5sr/9K/+lQxcKaCJ0d999zj2QS6XUXq+ZpmL1uClYqr2NjE8WPMnkgGkKfTu/bvx6ccfx5uV19IXB71KM+u4SZMgYnf/UGamaI7XcKG1n1NWC9SXmvbFlMhSSsPs0lTNfVfIMDXwSAxV4JffgJNryaAlWrAdx4t9YISRCgSGIdmlVBMzh36dhYheT5JCbmpoEKRmaAdbg+GdDJIZ7phJ4dtpJLkwNarHzeAow26zOfIzpCRY6zwpdH0WciUHVWvR3/dfn1HReX794FDt78yPYL71xNzcjM58BodiNxATU6ZCKHiGVimvxI0Cjc0ZWEUWjYga1lnPmyE2jIpxse8sHbOvZ0dTQ6cEjTUGE42mihIa8jTxNdiDIZp+TtXYqT3lBsmA3g/GYzGOOnXAGYISF0EJF8upBhb8Ojo2onOL2E2jkLgDwhSdaporsIyeLS8rhllykt51uyD3WZpSih0NtNqDrCH2MHt3ZHQojk+Odd3K2848qObsBoU6OzMZd+/eiMePHsXo4FAsXL4s9DXGwhWHLprnsbWxIc1/0Kog6Fi3SDB6CGCdeuQL6zmAtKWRc3h8qBiuIlaD99Bz5iaTn8pUuKdXTEjiMg00mkJ4lDXPyD2TqanBhKUIhQRtmE0Ia4Z4XewHnjVn5fb+Xjx++tQzdFXd5/JVMNPywk3lRGZXEW0NbRf6NRzrXNMaChODUiKPohW2I2eiDKAzf+jck35tbwI3dTwAl5xk6hSzDgWCyfOCZhlgGzX7QOYfHklmhAvhvLl69bIRd2o8dcXx4YGajqyhtbVVNdnUVK7BvXI+a+6zbsiNjk7O9Jzj4iRu3bqqtWAwhc3WkVzjXtMnWH2zon10cnQQ927dCFoRsJUPjo7jvLsv9hvNmF5YiOXnr+Jobz8evPduHDcOYmiE590TmzuHcXLWJU+4XnwHBDAhv9mJqYnp2NvdV/M/+jAghnmwH2cnTeUHsPCMlHW8ZL0sPX9Om8pMj52duHT5cmxu0OwckvQSbEhYkuhBkz/euH4tfvPVV3Hl0oJeb3N9Pa5eWYy+HtrxnO+AelxLGIxF09qo3jMkg2jownKZmIpnyy/i6dLrHALBgKWh0h3HDCtgq8t3wVKl9k+DVeU1ZZY2z7mdU6kEy/qBgQVrsNDNYt6ceXht0ALgIRqzx1qDbjq6RuKbxEU8j3jvnXuSpXj29InWDXvyyTPkaC7UuAEZyv5ZefkqNjd3Yn5mMj548CCWXjyPs+6I0dGJODk+VU6l8yybMMWGqKEya5s4h0QNAyaGQPblUTKS8nQR165d1f3AdNSedq4jyQlo4l+6tKDGsaVn2ix6YgvSPAcHR7GCJJaMgV2rGETSHf3d3ZIjuzQP+2ZEZuM9fd2q8f76V19F/+CwGZACQtG08/CzABAnxycaHqkhd3Ya+4f7rleSUS75Pvxocjhd4CmDO8wKJ9aJIS4JnW77yUmWxoxP0O81gMCPq2oQ9mP58tEs53X4In8VW5r1meul0O+szzqLCqRSbAkx2pIBW/VHfU8NlXiWxAq+Ci1ccZAhmOIiDbyUgeb7eE3eX8PQvl4NAYeGBxTDGBJyzlJ70oTkmWmwUyCPrCaoQ6lnGVKzZ9dWV+P+/fvap//Xv/k3Lekrs6XNeOR1CHQMziSfNjikZ2NWtu8Dg2gWvQbFp2cpfdev8w22BGtVLP7zc5lns6fv3L0TL169EoMSSScGRHs7O4oT+Btub2/GlauXtce/e/I4rl27Lv889sx3T76LS1euxGeff6bnujA7H10XXbGxuhGTk1Oxsb0T/UOY54aNsfHaSN8Z7oElipHybGp4bjNwN1RXXr3WXhfzMYcQbBXWopqhAjvY30g5SHoTuZ7u0ZrR2aP1XsN21xCWZU2J795esxpzCMn3Y+rOd3LPXTsm+CjrNcv8dIDwMs9kP/ElZmuCLctzjbVWA7R6rjL3TnaBZcZzWEI+cnzUAtJVs7/6AU6C1FVpDXfYk3yV96YkHRmiJpujanuduQkoMpDK53FL+aDFlcyhiv/ZLEjib7JRqmlc/8aZxXrnPW1+XmzsAq/4PcwMcZyvWGrwCbmm5Xn5TgPh3Ncp9rafefn+uFbUrciBpYB/YnZ6eFmgMymGIGuY0qCKJ8r/q8/hHLg+j0AgYuXD1PN1iL2roYhlfn2OucZ2XpwStAmYqtyvwHAanDedv/I+ZgVOSg6txSRKid66hzXoNiPMbH4PKprJYOiJ06O96Gk24n/+H/4kRvq6JDW//PJNPFt+E1NzV+Pp6/U46+nXvQKYJLnznh7vmV57RnFWS46wuzdGRodpTeoB1aDPwDJYdB7gcdbC/BbACHmqM/sa8RnX1tbMmG6eSDIKnzxiXPnS4QXFvVpdX9UAgzOZM97+tPjGtln2LQnhlkS0+28/DSpyKfz0y387d2Dy2CZKnkMYzdlC7OYwooKqkoFuo0z5fhV6mgo206ivEGZtGRJLktCg7oqTpumw/+O//LP4D//+/7GmYl9/HB0ciL7+zv178cGH7wuxTDFreY/u+OUvfxXPlpZah6vQeHnQkfQ0MbTkkE+TVwVrmqbZNGTi7iaAmQB8IjRP9XsQsBGaZHIQQAHd3d/XISz6rhALR2ko7oCtYsAQeAVUkonSfiZxgq7tqbeRPhwQvk8uUEqvs3NSX0MKIRXSDMka+6ZCVtNX8jA67M9ibHRE708ioQAvGq0RpBwiRrnYELR8E7a3tpQ0Sa4HmZ9eyyvAfEFCA1prJbzZX2wl67yHaHqdE20VsDZ6rINWuv4k0jn5Z/2AaNE6ywaaDZgz0U2zq0JCaH2BnJA0F6aPLuSUsDGRz2rejBoPkkSJ1WCqjPb8fRSbh/sUt6Z1UhzJ/DyHFz7ckQMp3wukozyZV2ma71WNQq3lPFRFTVQRQvFn1EY925qaly4q95sGBQm0Dl5ojyWjlK/pRkUWvzS/0MVFrziLVqGiz631TZEtBFR3b8zOzShBx++DL/xVQJoylALdxnpFb7gQ78WsqSSmnknzFG3Ytg4mn8fMJCeXRV/UsI4kSQ363kRZedhQUmFORIxosWlnu1lrnFOibiRbk8gxfSCjy4QKVCPdQ61bt27HB++/r7XK/y9fvZJO7MLiorTN2Tf8yjP47LPPdd0k7DSHVt680T3zM/dnYu3IaJI4NmS/AxpzGHVXPOR6MdCDycXAg8Eoe2x8dFToq2+/+VbxQ4M+NTMbQo+KtZEGztx8GTp26noKxe0hoJkRRtHyeW2eZUZFq2GtxM+JIkkYX9z3ViNayWh2uOpoygzQTAYncSookKprNPTznU0yUX2VDLvR226um6arwiTN4EgUQeeCKPln//Sf6d4+f/Ei1jc29R4kfCCHe/psOpwKBoly8/VKO5rPQ9ZHw09DDUzIkKToiX/4sw/i2tUr0kj/q7/+a2kJP366FOOTUzG7cCm+/uZhzM4vxsHBsX5+d2cvXr56GSNDw2+h+1xp1EBOhYgSdbPsykvJMdqSO+xL+4u46VVMOJ+P9hrpHFp6H5lyrmKApkEWBEradebkl37jHSAUujwljIR34WiNeRcPphZrAJEa5tqrYArOie1+zaIl6/Wkc+rrVcMlZdUk/STmomn3vE7t+zobqxB0sfBfb1ChQdQPfP39hxXm5eCTQJwWGGAHIEGfZBaE9AM1TL7A+dzTFY0js+dOz2jIENO7FEv3d/dyL+S6oPE/YN1lcgnnKH0a2p80z3SO2ffICF7WuobejaaaqMo58EaQsfeIBhIlV8J+9QAEmbkNS0slQqzknfh3nj/gDfIpXs+FjFF0NFQ5W0Bdi7VpeL6kK/7g05/Fo+++i28fP44+zkI9425UdMxOq6I12Tr2RHGxWsZ77OnRsfHY2NhUI+SwcaD7KNN6JDvxk2kYhX9x3oy79+7E1vqqDMWnpqbFfhVgBeNSNPvPL2Jnc0vIU+Qw1PAYpEA34paBNrFRA/nBIW0cBiMMbJ48faoBDPIZyLBoKIEMh3TqGbC6gcivaPGTZ21ubQVyN+ub62IOEIs94Aat7f1LwXhp4VJcv3E9Ntc39Jw4Q3jWeN2sbazFyhrNa67xQpIWDLwvGNQwJOC+56CwGodCBWbeU3G0c4lrEMrZWGi6LNbJz/iMJQFRqMZqIPbCYkm9eiFcU6aK/VxDETVD+0CVYnp9KhQ6wxvONHlVsEd6AATtx/37d9ScGwK80sWwj3OKghrm7YgKcQ2wiUPIiajJD3PABrU01bv7kELbjNMzgAfdMTs9pZ8b6B2Ivi77QyBLhGcUDAh8gwb7umNhZiYGpTNN7n8ae8cnsXtwHAtXrsZLkPsb23FpdjImxjFSP46JyZnYPz6Jbx8vxeDwsCQs+fvNja3o7euOa1evi+2AWSaDjYWFOXkxEF1BNmpoGV3ylwHAoTV5eChfI6QbX754HQuL84qxfNYP3/9QRrdEgtt37gigxDObnpyU3AtSMZgud+Gb0NcjiSk08rnnyjeFrHfTh9x5pM++AV2YvJPrjY7Hs6UXsbGFFwSIeed9IPYtGXUqlofk4gQOMctJ8hAtvykPwoodDENMOTAGzfLcMvq+ZEsYpDLc++STj2VEj5a2ZXF9BrGXdKbJh+ki5mdn4/LlxXi5vKyY8/7778V3T5/G1s62rgUWKWzJrrPzeP3qVZydnMbHf/BpvHj1Mta3txwXL5CRcY5Ovnv79i1d06tXr1vnSOX+gM5o5D5+/J2aOAybjNL3kUjzhvWP9jfIVufRDFpCHhEwyZ4tLWtNEx/FDGLFnZsZQyN4//BQTCmuGeammrV4EyBhNNAX0xMTMTU55rqtvyd6+vvj64fPYmcPFlJ/jIyS2yDRVDVFU2dDMQYww1aDrgPFyvqvM5vz1QwyGuS9OnMxW1aj8hyGyanPHENGDOfLnIj3ZB8y0NEAvBhwqaNPjr29tR3HjSPllEY8pxF3MupYw8QYD0Ms36NhVeYhyjWV1/RoPVSdpTyV4U/WjK71nJ9rADHowQ/vx3ByYX7BXkMDGNlPKv5w7/if36txyfACI/rMW9mPDFMLXU5tIzDc+blqM4aSPHf/6n4BuST+LMi+kp//+Z//uRr1Ps98LeMTk9pfMF96ARiWIgADmX4apiEGEblZb3ddM3EYL6PR9IwDgNCnNbb8YlmDQyR0qaVYD8QQ+UkdHYlRwTW8eLEcE5PjisErr19L1uzmjRtxtH8grxvydQYVfC8eFUgj4uU0NDwah0eNeLGyEk3O7WzsVkyvQQ7PjBhBbs45OTExJlagnmlJJ7cGRd4HHiB4ZcmrifUsKVaDYBggwVji/C3GJfeauldnVqpY8P00SssjR/kir5o1i9kObc+JFmQ+m+1t+SFvbw/0LU3N2uAaWEslbVd1aSH+BUykpyEfDdaSh5NiHwE4yb4Br1lSSwKgCSSaKXau9VYfRCxSxxt+Rnl8Dmp8xnLotg2rf5dNUS+cIUttIJ/NbWZK2+TaNTTx0QNuDwgtT11N/beZG8WYkGJF7hviC/e/wIGuu216rbwgawet+5Rjd57f9rpwnUK96h4OfRpqGT53+WeU7JTBne7BeLjNoBkAi2sWay8UoMp9NPUKyoskAa7EaA3lAaSqbvEQXX2TrLX4/PzZElCp+HF2JlAQDGcpiWTviLdl3ZC7EIPrfrKmDdboanlVchuGerui9/Qw/uWf/oNoHuzG5PhEvFrZiKWXazE2fSmWVtbjzdZuzMzOybdqeHTUMbArxKpj//A5eR+GmJevXFJ9Qawydva8lU8WqJjPxzAelqmGPjwrehEzU2JgERs5+2CHM4yAragYNjYuL0zOisOjfT0j9nrVCgKHS/K7X6+LxJVqe5Ga7Ykr76OfpJ9+sN786S9/j+/A5FFTG55NaMkWGoueeLeR1m580FRKYkKLnqomUAYcJQ1QWwcGVehbR9jBx5rJJMIfKIldXlrSBocWvb+/q8KTAosNODA4bP3VwwM1vdCctZaeCxIaZEI9p8+BkyGb+BKwoSvvbu9I703NPOm02mivij2OGwpVEi5+dn5uLpaWnkuypAYzRvrY5Chzypa5EH/HAMSNKcup1Cic4FOJdy2NakRV08aN/TbtjYYEwZqv0p9ED7MOIX6OAFf/RuLMgVT6puhqUgRwzpLkaDqu4jq1ICUFcZpm4UYOEWTdWK/DxPqnSiBkOIkxtHUVbQTclg3hOYjym002H/rCnLWMf6zj72RfQxHuEw0jJBwS5VLUYCVY0p488c+kVAWJvho/GJPy7EFSgLDie1PvlcPEVFR0AE2dVtOm2yguJAaE5kcq6cjITlM8rendajpmDqI1k4gBITPPc60lUs2NPFONhZQOm5a2ERiJxCgkRBqalpmzkrYWauP7wcPSU276W99wWIMKEgQhTZLiDKpGjYm8j9KxBPUyOBgfPngQz5YovFykWg+Wfeg1UNdbLKO6RhcWbmRpX6cRNNf6g1/JKpL3Q4vqnsiINEbXwEEImqR15hoSojSRNkKKnFrT1uwdN1TVEKY5ODYW7737rhppxA6agTQS7t2/n3r1RiCSPNDkevj4Ow9ckwbP33PYYw5qqSAzqmgInF4gMTeoJtvw6IiKEdDSTp6gw1uG4fbtO2aOXVxoqPrzv/iPQltWwSe/ldSV58I84KpC1KgjrZBkEynpKDPxDpSOk0m+74ebuz/W9K09Vgm7E2EjiKSNmUiqSqjbRUV+yo6MXOigTDhLxkQeI8SLUxe4NLxmpmYly8G9o2FzdHISN27dFCIdRhpyV0rKzy5iIA2sFY9IWEs67AwD6UijUqMO//DTDzUMQuZBPis4s5XUAAAgAElEQVSPHsfcwmJs7OzFRU9vTMPeODqWxi8MJZtoNyVxBluKBoul+YyENvKy9rD14YUUz3hq+cIadHto1DaGa0tqdd77arLXGdmK63kOVPNS9OhkLXX+PO9hFFIObXKDfW+vJWXbyG1L5VSx17kfc2l50JFnSCG2W8jtZG3Us/Xn8zNV0ywl13KRGttVEmA51PjROJAf5u3780P3y+u71nbHGk+ZBr+Uz3o/FytRmkFkXXA+h4a3XbAHzYZqyQC2BkRVpCWbIAEA1uJtD/ZKjq38pRT/GAgiv1LnBmAKGSAjfQCDC8k9o+JVjFPUwAyFwbF/kEN7xxjkZ8hTaHaU7J+0/4WUv5AJp35G/kGg1NPfQAh1Awy072i4JVOHIcyNa1fi/Xff15r/9edfxgXXTczi7EwEpovJNlKvHVvacagYPgYBJHBDv1oOpBikMmoEcX7jRmxtrMXo0GDMzsxmI8rmnSo2T06ENKXRBKOC5opMcWkuNI51PmsQkoAKob/TI4TBOg08ntH+wVEMDo+oScW9AY3LOmC/wC5hgMw5QKwh1tJMQZ6pEMTFoJG0xemZBkbkm8vPn2vfkft5bdnXRDkklW3Jl+R9q7yvgDxmTHqAb2BBIQrtR+VBopsWQixj6J5MHz4nyF2khyp+COCSTBhiRaeHVCciupiaPj9ScjKbBWKqaN1a6uHk+FhsW3xNiKP8nsySRj5IVNaUTG3FDrNWdyHwfe5bRoK8D/nIycmZ2DnYjb3DfcV58usemiaHjZgcGRfDaHBkRBJkR0j6nBzHMIOK2ZkYQkY05Y62dvZja/cgrt26Gc9fvlTzcHpmUnJhNIcGR8dia+8gll68DNKjmzdviZ2MTBRfU7PTes5q3vZ2SwIGDWlp+Hd7WEg8eL70XIbP5ESspa3NLfmt+Kx2Q4N7hlwqTEB+5Vpv3rwRz54txcLCvPIHcqi7d27FYF+XhhXKjmjanPv+n5w1dU/PL06VA9JAwH8FWc990JCjY3Fw1FBj/Rg5CeJOF+4difYVGOb7yOPao4qCeYY5XragvdlAP48b168LoSn2cp71MpNvNoU+Rx6T5+d9nUPw7l5LUQr936M8997d27Hy+pXyaUxAqZterryON2trqg9uXLsWYyMjsbmG2fhu/OwPfiamyvLKSttPIeWB2QPvv/++9ubS0pJjggYjZtnTFAZIA5OFXMzsBMdC4i51GHsKhpkalIn4BkRD7ACgQ+xV7pQDKg0IaFRlHUYKKcm59FAwTYl8j/0wFlOT4zE6MqwGrkEhF/H1t4+FbOfsoR60jA6gCQNbyreGNcdQ0P6EMFaaGibTwB4CHV/Agm7vSRsEw6JBpsfNOcXkbI7axy5NnysHKE+7Dmlanw2+VzSvxAbGF4ZnideD5NsKvWx5FMcJn3XuW7NKfSYUm1VsLHlRIq3ls3V6ajLv7VAMjwzr2cHgoeYcGrIEyZBYVAxrLVmi2CU/DEv50ZCEzYisEf6O0npPBisDA5+dBkTA0OKsk+xZ4yQOkJMTKOYoxsZHJeHiOr0nbt+8FXMz8/Ef/t2/jy+/+K0ZE4wne/ticHBYTFuG7LCouAk9vdQW1H4e0Pb3w6roiYH+oTSvNiOS50Ls4J6xRoknnD2Y7C69WJbBOmcfsRsW17WrV3X9yBXiH8g9wTyXcwZfjG+++ioefPhh4KPz9MkTsRBokjL8IG8dGRmL45NmPFt6LgR31eGFmGdozjW7Tj2zAgIghgHW5IX2NYN59SZEHDDqXusA6Vg1hJFSPVLTFJY5cQugAN8tmW8Zr3udcC7wc/wdv9e9g4WUUrkaBmT8LCS/2GQ5qPAQrECp1JlmAnpo4Ny65B9ZKzxf7pnlDD30V5wq8B65X342qTCUyXYOScrnoBr+ZvQhI+7GvdlC2b9JUIH2dacMXZ772g+p7KC6TdLglVW3f1vgA7MDYF5kxOjw+VOa6s2XINg2UMp1t/PfFiMyWUhcf8niceECy9ALY/h7YhZwi7mpvexgISZCDlx0Sug+pXxyfg5fij9HXVa7t9d5nVmv5pCrM1+UWoJ6DW1/jdYz1z0vBoaHs/4qdkhCE/H7S5+LytnNOnfsV16f/qX8NLH25MixgnXJV0kF8ucCsbJG1TsD+AajKKW+e3i/85MY6mrGP/9HP4vGwXbMz87Ho2fLsbZ9FANjM7G6vR/LK29ifn4htrZ2POSJAgcMiOWrIXzW0Awu2WfEBhgUxKyr167Jz0rDHPLQru64dfuWBvunTYAffco9kbVf30AZoDsuus5jfn7RvTWGWF0MsSMGh4bj5OQwDo8BXZq1yfsALJBc7QmKG/T5+HOXpDrpYfQNmkF4eHj806AiV99Pv/w3dAemjq3fX4h0o6dLKsjyEZ2NKydfyDJZQqT0C4tuXM1HT2ltZkjxSZH64MEDUS7RdtffYZ4WEWPjY6L+MySgUQ460I3rPqGDKAYojkA2E0NpxCshJCBnUOeFCllPUOW1oIOX9A1oSpIRppbHx4eZLHaJogWaD8QjybMSBSFIrNmpBjeHqlCu7YEF38M1OJj71CgjKFCAbQitE4H66mxoVeOfXwm8RaFVQwo0m4Kek0+SYdEWi9ruMbya9wTHVpOjC53XKWve0ZxOJENRBWksklAzFFKzNhGcljIwWphE3FrWZsxwMUyELQNFkdinRF0or9QEtpSQkxsnJR5KOHly44nv50vXmkW9sxHLAlXxr0QrDZitpdnQs5Chdxpw8V77aQyIzwnJw+joiAoADm4GUycksaCEjjEe83MFFSApCWcUrWeje07SUAiuTHhInLkmIZ1Sm7iVQGkwk4gK9zpzWNGmjGZmYqqrzC1NRW9zjr4fTDxYy3smNHQ2Oi5SEiYpmyST7EEa6xSWll3yEIJkGamNN6urov5XY4h34vl5CGWpLeWHJGnZRHej242Y+iq059thzygIawjLaEtmoolKSfko/q3koMwicHOvLQ3nV5WMSpp+VaOwCkQaCKCTKKR4PWIEhvXQsFnr7A0Zyg0OqLhmIEO8ALWgoRVDJ1hVaQ7I9ZOo8zyHR4eFsuJ+4E1DAsB1iWLN+52TMA3pe0H1Q83cWF+Lf/fv/m/JWLFHSai4D5J5UxPSpqrWTTf7pNgl7VjgxM6BojNB9P34sUHFjx093i8uUKpZ1441Xu9qUMjI1VIQ+veMTZ3N7nYjrK1nLMZF4A3UqxhOQXBl8XI2CY1Ma5w2Y2JqSsOinf29OD49NnW7eRYDXRTD6WPS5c/K2hwZHIozZEbOzuLqwoy0wYUIxkSxfyAeP3ysInF+8VK8XHkTFxRiAwNx8849odmIC+x1UG6Fen79asWoMzxLaLj2kwR6bRJrPFhzg7HOumJG1bXXMK+zSfRDjfdK+FtFRCIQKcqF9EyvJp+j3qM1tNOvPTmwyohQjUifK7UWaq34z/4cPzzIqmFCfR6/V/68DA7bA7I6f8p/pvZkvX5dW71nff+PrcH6vs4hzt/1vb9zDR3XW4NPD389qAHRPTjEPk5EVw76jCrCI8FIUuK/my9pRAebruJvSQkUijfPAElVgB5LGRf2O0VTsSD5tWSQrDXfPpP4fAIOdHer+cZ7CcggZLvXPYhGNWpS/lEsqjTJ8yDKQ/WSSAR5yTmpZwet/AhEpAds8Aru3bkVd2/eFXr8l7/+LC4w2KMhQN7kQ78WTx1BrTXPWvdZC0Py1D4RoK0Vr4yea/kYlRzB+YU+D7GzcXQY46MjMpAlzjI8ZmjOOc2QEPYHUhZXLl1u6bWzmCnWQJhy7nBvWF/kB7BWCl3spsmxmro0OMkvSspRuQQ5QBOD53HFXdYHe11nOV4MiVZUAzLFpokR5TO09JzmKc3DtmdVDWNVTguUYMCIGLMd26zWYcuPqWNvc99omPtZtnMgaaIrlnm4hU+Fik90iVOCw75DycCoRmbqTJecAh+n2M78vthf7YGSG0Mzs9NixY4ODylGIGE1NTkRQwP91oRWs8D+JXgzMehtHB8JFV1NHEAQoH65hzAHJ9BWnxiNV2+M/sWIeWp8IpoHRzE5POpBIY3/g/14jWRKV8hEe35mSl4VZ/IjOI/D4xP5H9y4fTe+e/ZUBfiDB+/H9uaW5IP6aJKdnsbOwaFi/ugo8q1uhDKY7BnoU1PPjDbhUBLtiLTCoIaF7H2dTwmMYQjBPdo/OBYymf0IWAVg1MuXL9QIgmmKnBCeKgzBdvcO4u6d2/Hy5cvo7+uO61cW4/TkSNJBQmUH8g6WBaN52jyzyTDgE96LRoLlZcmtemNjazter2LwfC4/hFNJ7HL+AsT43Thea846+xkl86juEsPU+5OmPjkOg075MXUZ+a4Yn8AR0J98P/mMfAGSyYv0hNl753HtyhX5iyw9faY88t69u3He3SXJG0zG8auYn5nVQGp3ezc+/uST+O0332iY0Wg6b7Okjj8bgwpqNZq61YDydjL6FPQqDV7iRXn4MGioNa7mKKzT/Lyqv1KLnTqFZ1YgNUmDZkO0gDW7ewzUPKgQSOaURi/xvddMMPbD0GBMT07o/bmHsDXFHtPrGS3spq7PTpkI09xFFpeYRO01NCi5VTOMz8SC4JkLEX5mNrxqBfkB9cSpWJCwjmHS+n6VZr7O7cwHibEClwg165rBjD43MxVnDw6U+/DvkrfN9WEGslHi3COpHvT3i83Hr8R44jg5LblqeUQQgwDywECREoAkL5FXa+fKYvT1mPnAmXZ6wjUPB5JY7G/iPueUfN56eyTNSrxHUovzEiYIr0/9zvcBMGNP6uyQyax945pNjNAt/8LwhZiG4gEydcRRvB4wpv7220fxb//tf4juvl7FFpuhT6gx6P1JPcrzA+Bl4AI5QfPkTLGFs7iAfM1mw8BK1cwXcefuXcnrIif28NEjxb1rNCRfvlK8u3cXs9zXqr0xxeUZK+6OjUlC+qvffKl1hkk9/76xtqaBDf2MVbH6RsUye/JsyWtMw+/sl/TDfjPiXbnqhRlQbuxbzgpGTflPulHdExjL87oyKc+9SI3EWjfoy/K01US3tBl9FNebBbTjfQqoYx83y/pwLhtM6cazAUKWkKovn601SK9hWfscNbDRaxOFgAJE1s9rnzNk0YHezh6LOaDcRL6S7TpS79cJrEqpbta6aoLMhVQDSPKV3o7VB9q+Ku33Q/ayvjoZFZ35r1kB2bRXbCoJZdda5S1Q+bhZElYZKNBBZy+oBooFfqjBn3osUjNovxexXjl23nbXETnskv1qSnm1ryLLvI4bmnVnux51r69dd/jFa5hYvlrtvoDBx8Va5XsL6MzrkDtTI3owkaYfCRar+FeMK4E9UwrTjE7ff/Y7so7lq1VrUICQHPCo/pN0nhl2Aqiqz3EaAz1d0Xd+GpOD3fFnf/oPYmvlZSwsXorfPnoar9Z2YnLhWmwfHMf69q7yin6a/kh09QOGPlSttqfclnVkpt71a9fjrHmqvU884ayH3Yw0nOrN8wv1X8gp2HuAHePCoOFT5Qld0Tw71vNgHeKBwVkzNDgc29t48QzG/uFeDA4BirS3kO5TAgEw8yY3I0aKVaPPSz5i2X4GoT8xKv7uqvOnf/09vAMzTVA9bjAXzazdQHOgEnolEY4cLCRdRAoCqORCUstPhxhIo0TXEbBAAEAT/5N/9CdqLn736Inoi7wOfw+9isT4u0dQgVN3MIllFFFj4+Pxzjv3hVgBoQPVm2Dp4GXksyaJQsr3q1ghiWdQIWkIGQseCYmjw1u+BBjcNGNyYkpNXgz3KFRIoGjqujntxKCFdksjbN8HH+oE6mpw1USfgE6AosH5dmOr88/t1/GiKTYFvy9khzwFJLlimaCiV5Mo8hlI2Em0hJJL2h0BkOSRZJECj3ukZpzQ6jTrzyWBwesVO6MGCCTqGA/bcNzslGIqcIAIfXfq5KIGWJbFsLEfiQz3W0MFyceg42f91NLxq/fiXkuaQsg+e25wGPPvmhbrBhqV2tk4BdHHSKFYFCSKfCbrGHo9uGBAC7JPjZOTYyfBKjASccCbdjbj/RRS7z0PQRJl7mElfWUCRfHcbmTqOM9GtF+jmtIVDnTIp8SYqZUUHD/caNQhqyLGhzXXIXkroRk8wNE96jb9kASUw81JfL/+p4jhWVEM0PSlSFUhmAlomaHXfW2ZcXXIOBmhbPxVZ3rTGeL4uUKl89qWsfGwxMM2DxvVXKKBUB4teemuyxL1KxkVo/Wr0a8B3eBgvPfeexrIXL50Wd4UDCrUeNrf16HN/uVaWTcgOkmOGF7xWSiEjESybi4xh8KeRGBsdDz6B9HB9nVoLx0dx8jwqO4f8hoz0zPSPeazIDXFevw//4//Teg8JVVCcOfzz+SaNSNflvSmKRRd52Ds+3e1oxFd9+NHSCw/dsQ4npQxdtsjyAlgyjlJgsONPz3fH3i2lupz7NIeVwPmXEgT6a8y0FGRx1BmMBbnF2xunJrde4cHsbWzE0eNI/IzS4mdXkR/d58SV7pLNFsYpPFPJJM0qe7fuBx/8PGD6OlCCuYkpqZm4/nzF0Kc9Q8MxdXr1+MhZ0SjETNzc3Hn7r04bBzHq1cvtU4XL11WAUBxyYCSPcFZwdoAHen7IChhspCINTDUPMywHrybB2USWffz7bjtpLxtQtcZnxQXcmhdw3QSSvYB69oSY9aELd3WlvdENuX9em/HgTIdLHTS78YPfq4GwFUc1DVVVeMCx9i3QoXJnC39NHjeZoF4oNIuZDJCdlZuP7AYa93UPanc4e3XUaTM2rCuxNKBbcSZ8wmjivgsSE/Q7Edagj2GhjVFOJ+fOOFzwOZzxHqKAs76AlP4nrooL0RpaSSzV4mdvH/R0Pk5TGgdphIt2A2L0RJTYl9o+GxQAN9jb5O2VBuDTBoxmgm2htoUKzRjehSXKKgLZW/jVBfeI8NDajwcHsEi27OHxDFyP2fx7v3b/y977/lkW3qd963OOaebc5yAMANQpGSAoqgiS5JLdtn+H+0vdklVdpVs0bIJEgIpYAIm3pxDh9u5T+fg+j3PWuecOzMApW+Gaho1uPd2nz5n73e/YYUnxIVzF+Jg7zB+89HHsYW+fW+fJZug6Nee1Ew+vZ5tlumVX3NY+1LKzxUzz8ATn3Mu+ruoozOkIySDB/KU/RH0M+MnLevOTvlMsCeMjY6lzGSX9lXFEMmgKAkAniPPlHHjNTRjeK5cz+Gx938+l+Kcz2EX7EGT48eEBBgUe9hw7CtqfqRsmueiUaXEeXz2w4eP1Dh2Q8rv5xOc93WcUnPWRQyfgN77Wv1BFbgSTMOZxVnjoo5jZRXoWPdZ2GReArjhPkDZMmb1OVWsZayRG6vP9Fx17CA2ZgJJiuFZEhnIRSUpTOOHTAoSnwP9vZIcohg5Pjoi1D1MBLZh5jixmiUMzFBl/VCsg4lJ0ZIvmIswBSgG7hzsxcGxTetHBoeir6Mr1pdXY2xkREjGjUYj5pdoVHTE9Nh4jI8M6j8iGc7n7d2DmH+zFtdv3owHjx7H2sZGvPferTjYpSF4GJOzszG/uBCLq6sq5oM6hg0LcIZ1MjE9FeubgGgwiT1WUZAYmSYgoCTmB+NLUZPmFTE/18/z2cX3LmBbjwjtj6wE486cRaoIJgUAhwvnz8WXX34RZ8+e0x797MnTuHH9gs6pbhp7+9hku9BGkRoz5t4++xTQnZDXGybu+KbwLPET6e6Nh4+fxgpIfIpkyVTV3GvvhLXvp8mcEVq6tUE2m5UC/+jzbAbsBhtNmJ0YkinxgIqsYOiXlt6YldvRJWS14hJis+4uxUOXLpyL6amJeHj/gZhMI8ODMT49KZ+u1/PzsbXeiPGxkTg9NydpJWS1Hj15HPOLSyrWi1TWBrA5ffq0cgD2gDKZJjfg+lQgH+hXo44vGp21DvgZa1SyiyVDpLMqJPNm0JQlSIjheJ68L3OHPIc5QE6x9GbZq1br8Qh9LrEn8Erg1EZ6ikJ8X0+PikycfR99+lv5bdAgNagIWVzWhI2i2cO5UdYhY8g65/OYS7Ce2VflMYFciMBbKal8bDUCrg8UbeViAnywhySSv+SixNw4OEiJWs8l8jt0zA3mSfDI8bFN1LuNgudaZEbd3ycWH8xDxbw0DcjZ01fFG55zu+MDy+KxX1pqyR6TOlM7OgX+UK6QICb2ju3dLY0PACGuFdDA6spaPH3yrImM53p6e7sly0csx5ySR0dKVGm/S7Y99zozOxNnz5zR+uVnPFP+AziEHMvjx4/j1u1bkomm+D/D3OzoVA5w9969+Df/9t9Jbg3G9e7eQXR0AcQKFTAp5LF39yHxlZ4/nDODgzXvwkVEWG3JOto/2BPTijkMmwiZs5W1NcmSLSzOaw/AS2V1dUXrirFnDQJ2ZI+HaXj366/UoOB1nFHXr13XPPr4408Ue42OjouxKSClAkrne7wP+Zr87JC52TfToTtlhcU6EdjOMoqME2eLDIAPyQ3xGzLogWcnv67ebAJ2uRFSDfdas3xP7KGUQzabIiWNm6oPKc2TDOGK5yrOrGa/AYA+VOu8rnyWPwu01gQGKSVo5dMlV0perzgtwX3NXLFpFG2Z6yqUFwuauId7Z89kDNUszGCzZJxZRJY1S2nnYkHkniFGRRv7oHK1ivMqJ7IkldmThfkqX4b6XuXzVRNg7fhnJcnUnuhZfYAve805f66Yot6rWCM1X5WzpXScxonxbDPPrppEK+esnLvlh6eGRD47P74W2LLpJ5Lg0fqZm3ptPqNteaO9/Zz3FGBEewnXmb4g9gR0/bHAmRVzMlc4q2H8FWukAINqbKSM4ebGhuo9PFvOK9WTBCjYDbiLxzsbcfPCmfjJe1fj1bNHceHCpXj49GUsrDWid2gyVhq7AvnAbuLakBCWdBwqFHjD7Wxb+YV6y+5OnD1zNsG59t8UWCHldJlvAkeSbwMKRDZKwE2z3WBJ7e0SFw+J5XX/weO4cvlCrKysxSCgjOgKmuywostzkrnMnqgYZndXrC6auEuLeK3hpdGrJijvKUAvze3vpZ9+V5nk++//oY7AzKGDFjYLU9SdwBp90CrGsFDVpEitXumpF2ovmxlaqNvo8KNB6OQWyu7tm7d04Ny/d08JLok5ck4ggghqSdooKplGfRK9A0bcs1mAasZgm8D01cuXKqJzGLMhuAhJYNsrmSiSLL7PpqVC+IERzgR7JMNClGURms2NQIiiJ00NCgDVvXRhuM3MGu+DNLoVCiYpxrVJ16HMBs6mLGO5kxaqwGdHS7fwu+aKiyd+BvKPSGYAn1VeBWzmllAw06LQjDwX7l+apDLBG3DRJYN+BWupd4xEFDRe3pdNnmIARW6C4KbhUzYxJMNE0ZcCR2ZL0s6ujn6QTA4lxR55KCeD1ZSo+xZiH6Tkzq5MMLlHDp0yhm0v7Ls41Qp0ZIgXdOj3spBBkGEt5QrqB/sHlSjy/irG0GACQaJD0YiRSnAsv+GuO9cl7JS02+034R/wf0av8j8FQ4nm1HPMxKyCNRUyO7yGWoe8/y4Eh+SvQF0Z3Wy9xe8u/5fWo4KZRAHzHjY29e9XI4h7YcyFfpV2vucHrzFy2gVR5jYIVq63icpM9JZqL2V8n3JkhZrxHlCmwN8ujApF2gszx8wm5qwCnmx6FvumkChl4vVNtIxGOwM4Sbuhf40nycFB3L55QzqxsIA4rKVjC0q1o1P0ZzOR0M/tiwUZLmNS6bXkhMneI/LIiNCcp3mFFiTIh+OwDnfpAiP7JK3tjY04e+a89gRQdki+sHfdvXc3Pv30E0kHkFDA4uFPF7P9jNj7SqNYgXmtl7cYPO1Mq/8SRsV3z5uad+2MCq0FNfqykJASdtWg++YTrSKxANnZkHUD1BJpZKwkEJcvXoqJsfGYfz2v+SSWUnQIUcu+2jcwoIQOVLXmEkWUDideKh6KDX4cXaD3oiNuXDodNy5fjv6+HiV1585fitX1jfjk0y9iaGRMiDxoso+fPGnqO3MO/OSnP4mnL16oGEVzlj2F/0jgKHYyfzg3OF8o4HBPIC35n70pnAgY5WTEnRMoMwqFLMyiUnuzon0/r7/Xnu5muEJ5J+6ZdBQtvpBWlnxJ5iKCDJlYtPbWMkAmmK+mRTURqpj57ZOkWVTOJoP2jCxOqJlV2o3eAI1ESgkY71+eX13oSjfR3S2Jm+9qOLRfxe9qVNRr2n+/ZJP8PX16ov3aOpmp3c7kEUK0Dxq1z3Y3KigMTMWpuVMqalDQ4RqKXaY+GQhrySKlYX3GO7W3sV+KPs7eiXwAcxpDScxqaTqqSW9JADU009RR49ll1qDmUaJu2dvrrAZswd7EdXG+4h3AF+/P+UMMwnxFeoXCK6hUmeTlucQ+RdNvfWMj0aFIcEZcOHcuLp47H50d3XHn7r14vfQmTpi77L+UQpqNijJU9F6uXgPnSTbutL7xnkq6fPlJFROIJMvrw3IC4xPjKtCMj42qEDAyMtZEhRNn0cCl+CtZs9IVJqnstSwP5//mxqYkaxQ/AmaR6fO5eP7suaVCaaJQ0BVy2YhO5rAL+uhU76sIi/8Q42p0pZP1Wiulvc1Yk+BRxOJ9QccSnxoEbk8lrwH7ypTcmB5Ss2nsJgFfkgXNz+LfitvSs6pivCrCSLaLtZTFJz6XmIr5y75M7KlGWja8XUCsOLG15qvZ3NqDHJsUgKKAI55X+zGIZML+bgwghcT7UwycnNT4DQ2lZCjo2FwPipFptKQeOOclhdn1jU3LWTHm7GVdnfFmedkyikODMTo4HLuNhoqGQyPDsbqxFs9fvFIxe25qMsaGBmJ0uD8GByxjsbS8Ghs7e3Hr9vvx648+jZ3tvTh3dk5nKJ85OjEeiysrYs4xjy+cvxjrq+uxRoG/qzMuXLwYrxZea0yRrAGURGOabyBvAgKZL5oXxP8aD2nQj6pwiY8S3xfDYnNTDQoASjTcmJvEDxSueX7ybBkdDTBZQzRIu7KRBfs6/dYAACAASURBVAdBsp0UqA5trNnJswgh9z1PtHrVGACQAguQz3z8/EXs7O6rWb4PwKsFis3tsf1sd8PbcWLCRfR6740yh00ZlANp+Rs8xCssC2FgEUhsNXDEDO/1M1Zjg/WMJ8F+3L5BjDUXy0tvVBRubG/F6Ph4nDpzWlKrL5+/1GeNDY/G9avXJP8FW7exuyMZGz67ikiML+NHbCV/tJRHY5/hP9aifLASCMa/Hd+62CcQ2cGB9ruSgVGD//AgJicmxHpYXFzSfZLTVfxBkwl/m+WVZclfWL2FZ3GsvRBvIRrdMCrmZmfUsBsdGhYTB/+Buw8eSc5IjJz0F8zWtEErkjCzt5eANJLiwzMMWSFibue7jgdKutBMeRWNJYXTMuZ20fZQa5O9kThRDcNEpBOr0EjimYHOZT3SEKGJwHqnQcC/GYeKjS1r6L2BuSlTbmScBWbb075Nc438qfJdXXtHp8YBxgzvTX5IU4Dh49phAfB3rrW714h+tNB5DkiggOSnoaNOaAJ0WFN8qYHb3a1zzbkrzxvPkL6YmppQbq/PHIGZxRnfqUbj2hrGtjuxs7MXr16/Vg4/MzWl5j1+Mch3nT41F1Nzs/HFF1/Er//Tb2JtY0tNwc7OnuhEzpJz+BjwgKWEyRvYa+SXIaCl/RXlAyXVAGv+F0iDvPjUqdOae4tLC03vCuY0ChBIFTKOp0/N6l7ZM/CqYK5R6+Dsv3rlSvyn//T3cfPGDUkhwgIRe67Hnk4wP2BZOW81+xqZLHnXbG3puQgAoUKl/RXVxDuECekYhfVH3aOnG+CNC64Vw7pYb2CS+FN5ptWZWWoZxaTnd7knry8ze8hvtOeQW3V2CPjJ2SaWdcbR3sCyqZ8q2Gb3GADkJpHZEo4p7B8jAF53q1gvoECbObVza+eyyOgUaJPPajKBm/EZHkyWu3bzM+OCzOvtZ2OAbQHM3DBoMSjt1dfKjNpxOXW+83pyHud5buhU/qUdusnEdJ6hOFGqBQkyyj2i1chB3cD5Y5lxt0u0FlKw9lI9yWRNtBo+Bs5orDJ2US7hHakJyMiDptlgaIY5imVL1ikZMJkrNZsvqoEYaMmXzcNbMVM1nF3z8FgTG9eZpf2tjc3ueMoM3vLJqvyHOQ4gjvVpKfpjrSspIQiAOKSfoV7C3zV/ia0zR2W+4Ue0u74aH9y+Gj+4cT6WF17EzPRsfH7nYWzsnUTP0ES82WjEHo3a/YNYR1pYwKhjMUzFWBI7yYA9vubm5uSbUbJTvL7iucqX2B+J5amF8vvknOxZAz3dsbK0EDeuXY7337sdn37yifYMS0Riun2ifaujC+URPwuaNcSHyFcihczZvLvXkIwUsevY+FC8fPYyfvDujejt6hZA5ftGRc3y7//8r2YEpg98eDSDitTed4ezOssYMNmQUkEQaMvUBNSGL8SjZRYkQSKDt24ViH72s/8m1tfW4tGjR3H69CltnNLeHxhU4MnPZPQ7NGTEDJqVmByWWZ0K6FC/Lf3jANeGQJZGMNVVncc0R+XQ0AFLgbKzU/rGVdxnsyTAO3v+fMzPL0juyQmiUbWgJRTsJZ3Xsjid0qPlvWRKnSZObNfyDQC1ILSPAzvQYyQprl368GhLN1wwKDPhlLvxpu7ClYrNaS6kf3d1qQBI4G8UtwtKoNh4ez77zZslNS4IFGGhKIHWgcbYmFnBuC0tLWrDowGAljSU0wqmiUZJWpFiqIZENbFcVIJ1Yw1Sbd5idfSbipoJCAeODs80hTZCMZHKR4cyP1XxEuo0plpcH/JgOX4MFAcFSaf1pZMiLRNgo0c2N9dNmabwinTY0IgRn+kLQCCIESO0f4I+I5zLs8BUUHe9LX9Rx3k1oTBg5T0IBF34R27Cz7kSAX7RR1c+y9TnfBuNkA2XnLOm4+eUyLX1zY2E5ymkCFTvfDGfy9hbCsy/L8+QKjypq2/jXcZdYylkqdGPBF+gKoWcIsDKgo7uXfRza4CCPC8KfzXdqsnwXRueAuLUh+f1hdapYmmFrk2aO+ybRIzo/doq5SUHxfwztZxG3FD85MMPhZ4kAQahR9LmoNrybhQh1BxjXaYnC2+tZ5nBEk+BZ0mSVGbmDtCcxIgZBsKw13JvFCLQEofSznhBCa0E9a//+hexlYg6GyDam0KNwWyQVV2hGk1v3WgOpLeFKgy/Le3zFnT3WwP/+xoV2RhjLhRyvGRIhJo3SrqKBG/ZbydyUbtdGtBpX5M5sxMpEgohoLu7pRWsAm3ST9lPQInzGSCqV9dXYy+TeMkgdDhZ5D8aEhjz9nScxHs3L8fVC2eiE+SjjPYGoq9/OH79yWextrkTo+PTQtfiEfLLv/2lEHXQejGH5XldunIlvvr6azdUhR7rVRLMs7eXUcg0nT2QgtfC8hvLFqaeKEVi7R0kFImOKbaTKNwUMpt79bdXQesZtlgoZii6WGSWgINtj7vfozxYvH9UgcMIp1rjPlPduLWXhM3qhChuXzxtl1XP1smTi55KUpMhp7PDKVGzCVko8moYqNklk1Oju+p9qgnxu4KfKqRWM+KbzZ36PY8ZYGMnb3WG27fJTQuhiHLv5VbZk9VQpmKYzAgVwjjlOjtt7Lm9LSS1EPMZjzQlENPU0B44LbickujcI/k2DRoSM7FLExlvtp9l7tCN5tyy9IZZnRQBKcALVbm03PT+4FmC+mQczJjgfLU8ldBk6PAO2S+KgruLEzbVZm0Rj4AKN0qOWqFR+0cHezE5Nh7v3LytwveLF6/i/pMn0UXTmNemzGFrbmY807YntAoV7JsU3CwvIMaEWJJmkvjZmBFHYZCiDk1ctMOLYalGhrSyLQ8l3V0Vs/g9M5loAEObJ0YBefry1QuNu1GvB0I5P3/uRgUFXxmMIufFPMzCkouzFC0PVfShkESMWWdPNVVKjrBYLqwFCkjcA/Ge2E1ZXKgiihLwNtZLLa8aw9ba8PzROkuWifeJTLjTj0txYcoUEX8aCEIM6f2b+JdiOV+c5QV+oTBdjBeteUmeGYHZWn+5grPBx3tI81umwb3SQ2d/ZB4gNYVcEawHUNwjYyS+jgd5ThSUC6BU61Uyn+lZwrydnpiQFwiyfsxDTGOZl2pQDAyo+Q9inYBoYfFNrL1Zj6nxsZidnojhQYqqJwIPLL5Zic3tvRibnI7Xr5fEXCQH2MXQG1bj4GA8efkiVja2g8cxMzMX+LHsIgdzeBhTs9NuOGcjjlhS87J5ztvnhSIucaXlKlw0ofCws7cfL1+9DOQTmJ8U4AAfcC4gb8S8X1lejjNnMbnc1n2dP3sqTo73o6+H3OYwDvcAP8GQynO4g+Y3+zEeFT7jxNQD2Z0Niu29vZiYnJJ5+MvXryUBJUQ7+3CiV/2XtxsVFaNot060a5MpkBKPKtTvYSxrQIGkQhKFKoarDGvd4ONnljzBUNieZxTDL5w7K3mLU6dmpbX9+PGjODzpiOk5jLZPy8x8eXEpGo3d+OG778TE5GTcfXBfzQzMg/d2XWQvAI0BbS54Mv7slVVE5xqY+zBn+HxeQwPPrLdjfR7vgwm41oZYKT6D2DsoYlO4Jud0rNyd+UOf0OuvX78SC05jm2AcGrsUuMvrYHJiTPHkMAVqpFUPDuLxsxfR09Pvhq3OAzcfuD4hVwXC204fmmPlqKxLMcQpRCGbd3gk3wh7LezpOiyxWzmxJeAoNvfTNBwe1nUwVylqw4JQEwIfJDGcbGZNo7vmguMWSxLKr4UYK2NmzgI11BUjmFnI+UiTkX2SphyxkM8/g4NoanFNNHIH8Q48OdY904hWDn6cUs3pq4Sf2/TMrAr1xOkw1FberDZ9EYh1uH+umffFvwG26+LCvK6HmJ7COp/Hnie2aVeXGmKAhWhUHJF/HZ7Es+cvY2GBc9M5GOM/MzMVQwO9MTzUL2WG6enJuHTtmhoDf/u3fxfLq7ClYa/AcoIlnR5XnGmZB8sXLE2E1TQQK8mxh5H2lgSlMMr5zX1y3nH2ffXVl9rXz587H4uL83oOACUYJ/w0YRhSX6DpTlMMw9yvv/oyRkfHYm52VlKN7K8jo2NqkK3ISNexJ/syc4295/KVKzHQ169zkmvh75a5NjtRa0rxPD5WgNSI8ywF0wJSeh6obiOEgiUDVT/ZQ1bMclOcXdwHz5tzwY0K5/j2lLIvpGtASI0lAEmyaJYPVr6Z6HhLH7n572tpRn7NZobPGl9fFa9rr3b87NyqKSlevkzZ+CwEPutf8W0ChJDlUbwArirzdbbWYp+RC/NzzggBK1NOS81S7alWLWjfi+v63UjzmSLwSxbtS06rwkrHDC2Qb32/Hfxh0GEV+Vv7vnLblG7j9wTIpLGc3pECLWSNwDLLyQRPf0nGgQHXuDX72wYAVV7Rfp3KP0oGWudMsUxboMs6fwqsWXFCk+nXlluoZpO+mS762xOuYn7VCHOeFGCsamPONQ30c2NiOI7xvckzvuYptTDNt5wfJetOPsF8aOw0or+nRwCDg601NSrOTQ/Hwc5WTE/PxMdf3FWjontwIhr7J7Gyse5GxZrZcfv73tdhaOhcOjY4l5yIfQ+WB7FDAZbYx5F9c93LMRv7G3VNgSR7umJsdDhwQ9pceRNXLpyLf/LHfxRDg/3x+NHjePj4cbxaWI6+wf7o6x8IyJ/7B5zXSAvuqrbT2DLY0g1ozvuQlCAgkOHB/hjp71eMd/nihe8bFb8rQf3++3+4IzC5b71M0WSbxY1C+yZ6R4GTkS5OcI2AYfG6s1tdZMuG2JBpN/7iL/8i7t+7G4sLC0YtoSUOpXNkVJQqvnYa2wpeCLJcoO+UZAhde1P0MWAb0eGsbnzq+hI08PlCFuyDIrOcEV86dNMYqpCVVSzl8z/86U9iAfTQk6eWt0jUGz8joWZzkdZxmkNK85rmRPouZJynzb8623UaE3yTAAqlWkWRLPaoIZLFat7DSLk0sm4aJPrQL21FF8YtwUMSWvRD7qt/cEAUfYw6q1HDZ9CFJchgvNn4SWTYzCmwEmRcunhBQRUFBzZ9GXIlgriZEB0faxyMBmh10SWLIk3I8hkIBdg2bSZIaqGQm5r0aeBMgsfni6K7C/3WXhkbm+tCDCk50DM1rZmCUJlOMQY1Z0AGyaBTz8eFDQVh0GV1yHcpWW8WeJJ14/nipJ/fN1vERRjQKhz8FE4ohnEtIB6ZHCTEPNM6mFsFOYVzPuhljNjOqPAsaQ8OSrde9M52qEbb9qHxT0QIa64SJUB81qM1JbYSQw7HYtmUWbebL3ahLb8JadYmRbHQMwpqcn6Jnp5JruYCTZy8/lpX39zlFGpmIcDBiY0aSTgKXWFkRRZ8M3CqZk8FqxrFRN4IySMjsYN4/713FdxzXRjVbTe2hTBygmO0AwlAoYdYM9IvRkokG528txN0M3Js3uZnJXSGDn6Kct5LeA3BPImyi9cgNL0fIF1HQbGQqFyH5cQKbesxUNMlabIOJJ00tn85eHOTtRUU+zV+6VtthPYZ8t2HjWk++s9UdoonNAMtb1FycpJp4xrb0ZzZpPBzcHLhYL8jGxVGHZFIsU7ZF5CdYV8BHc09iJVCQKmiyJGCKPZuozfxfoEZBejuOPpA6+/vxZ98+IOYmRiKo91GTIwOqzg5PjUb9x4+jS/vPIih0UlJhYyOT8bNGyBQPo6RoYHoEfsM5lhfXLx0OebxLpKhLs8X417TpXnu7IUwZLjGtc1NoeyePn/enJ9FUa5GZxnD+zlk8zPziO8qvDfPwKbRdY5hszGUFPX0PvLyduHJyY4Dd3+1yfGIcm/0WTW+lFwJ8Wmt5e/6amdU1D4BitYyMUamiyGXa64a6YWAr+Ye64ICqs+FNiO/37FvebxaBtzV3PjmNVbhl3EeGrYBtRM2I3/9bxenmWcq4jZ9JWggu0npYuFJTExMxpK8ePZVKJTkjhJunzUeD58PKvbnmdvefKk9SnKBIBALIZ+0/jJjp2mOFBNrCTRlFci5F6EyOzA4beizzAg9jInxSSXkoFIdR7jpzefo+icnxYbUHtPTI0YC98a+QhG1WCb7Mn/mJjjPd+PWtWtx/sxZxV6ra+vx9x9/Gh3EKN0U8y0R0jp/jOyrfUrnSxodeq83g6Tmi3afZBvZ38fFjNrvKOTS0EFiDUQ7xQEV+pOdw3Ow1IvnDY1K1uKli5f1WXzvzt27TcYFBciLFy7Gg4cPkg1DcdLsJ+7ZMl2eSYqFjk+EbiWxpTFFU6VQxIxX6RQzvjYjt2m2CooZgxiUkCbDnKf8j0JE7t/eiNtZb17XhdbU/Mm4mXGp5jmXqQZFNtPl05XSZdKdJ85NU1nOCseavsaSvSjDbjUZM/G3SarZXgVO0R6fJsowGoT+y4acEajExYMqeA6KXdgbc3Mzar7T5KewC1hnbu6UGAEUbgzIMGqWe8FrgDMYXzeul/UGg42iL4kxRSyZ9B4eyL+Jc/ezj7+Kwf6+uHThTAwOdEVjeyP6acLt7sfm1m6sbWxrHz7cPxTSGGPnrZ2t6B0cjPVGIza3t1U4wODy6OBYOYIQ+UjHYIoLg4D9IgvZjKEZ1Adaf/hZKR4tk3CZmncKuYiXFffGvT9+jP+GC6ac6/weSG7G7sL58/Hs2bOYmhiN0ZFBZlXAXEBLmrNM8rZipMAkBjTVEz0pG0aTAsS0JN8AOR3AzNqX4fjrhcVYWFzWXqRV2jz/Kw5I+EtOeJ85Zr1pLmUcIeAQDO6jI+1HJZ1aQDHJFmrf89lNkYkcAKka7QMCY1GAOYmf/OhH8fDB/bh27Ypkw+7evRMr6+sCGmAUigH14vxiLL95E1MTE3Ht+o14Of8q1tnTxEiCtWRwGXMddhRzRMCqzBNoiMBMpbl4+uwZFZZ5PfI3iktTVglpC54F/zXXIH4F7Ee9fWJNINMFs471Kj1+QCodnZLzQpaJ+N+NV84Ux8GWHTrRnJ2entK9c180qLa39+Lew8dqZimnS8Nz3qeJApc8rfNMZKg2G1vR3QfYa00yRzCBKRKfPXtGCF/mCbkNDWzObT6Ha+6SFJiL4pw3/A75S/n/+QwVLlvPj33fz4+CWeryA6JLFkrJqXLW8bmW8DHzlUaG8s3OTjXAX756JQaEG7nJqkvpFsaPcYHBB1qcwhvXh8zi65evXLDGR6LjWA0WzqbzSA8eGJhC3Mzz5izDtBpAEJ4O7Ak0lV20tr8Q18AYMneRNJTvBOfgFmoJsAnJW7rj3v1Hsbd3GJvsFxne8gw6OvAc6YmR4YEYnxiNU2dOxTvvvy8Jqn/7b/73aGzvxYCY/kfRjxfEvrQYxa6wbC6xlc879gj79nWLbcQ6palVzdurV6/GV199oTmNRBVNWvYYQJfMcb5oBtNsohlErYK96NWLecXep8+cjjtffi32CGcWCGoBHoZHJTODDwyNCkludrowDUuT+OXDDz7Q/opxPXtP5XdqiG0j7+s8VvWOXrwqaUC7qUU9RWs/5WFgmdFcRbWC39cempKkmoPpDcBZxBmlXCClmCXvnedYSUQxT+V3l7KBnIuWSS6PplRXSNZBKXSwrWlNycja3g4CgaXfE/kD76HPTCBXswaSxWmuu2o/7N0luag6jtjBalP63KdmlH6YJZ2tmkY2PNhdS4aVvcSgnRZ40WGUgw9iD3JR+S/A2k9AyzfBQeVdUXmfGLKAv/KeLIfka2zdY+UF7RGzmczEX2YM2KSc3YM1IxnPBEioVgUrK3N3se3qrbJJ4Tyz8gYD0iputz9dC1j71t9LWioBFeXroeZJmwRuYnKb4+K54DNS8b2ASZ7jznt9NboOKTG4dqA50IFU0kAc7LmWQExfcpv8HmNYuXc1a5A4U/ODOJ55tr8d/R1H8bOfvB9Tg92x29iMsbHx+OL+k9jcB808EjuHoUYFi481Q+PPzRszb9wM5Frtw4WsG/EIMlDlNzo5NSWAA2NI3AvI0TWLNc/FroixkaHo7YxYW5yPm1cuxdjwYKyvvIl/9ud/HvtHh3Hn3oP4zcefBKuGuGB3nybEcBwe0oDslSTozOxsLC4uag8GNHh0fKD9j3h/iMZwV1dMj49936hoX0Lf//2/jhEY32kh6URTSwmXKmKySbApcEBZ+w89SwelVVgg+NCmfXggSRAO8lu3bmlffPL4kSjaGGaTVLLhkByUbiqJlDbuphwP7AVrfCIzwMIvwzQlbtkxRoqlOudKFBP9zoYu2Zg97ssoHGhT6CVzcNy4cSOWV1YlGcJmQzFfMgxZqKwkUUidfZArUHOhkrrxUJrUOuwSpa9xSKkPEl1QK5ljtxCyKSPk4r0RjqVDVwUqHSNtxkJskIUyqOJWu/QTYyr68OGhJE50nYlEZ3xcjLFWPveuxgMou7ExBRVr62sxODTcRPfKfCypl8xugpsKIEhyHJw4iCljb5KMkv+pRFmBtk/7ppyCNKdTgsqUUuvDE9h1iDrv4ruSHbwKKDapqGCZKCHdj4/VgOC6CCrQYsV/gmDNzBYzNUxz77HOK8Z8agyAqhpSc4YEUpRFpIAwa0+zZArUOhAxXuugIGJkDUEsz833blaRA5jWHmB5ldY36yDmEK5mj2V5KNy7+fRdXwqcElGgQC4bABSWofdWIlKmZIUs4T1d2DTrSOsptXFLesoyaS7gFetJzxJUTPpi1N8VqqXJ9u9qqjDJC4HRXsCxCaSZWuUxImRsGzXdBtTIqiSSJdeQGlnj47r+f/yP/ySGBtD/JRl2ca3Glb1EJoVqBJg9wtgpWMtCMAE4Y0bSJjkwip8yyXICr/Wt1/s5q+C+Z5m4kmnxc/Kz1frS56Edm6yvNFqUBFeiHB3otBCw7Q2Zun7LA7gYTrPLAZ+rqWauEcg78JZkURaNC61TzJ324nlNwQoYa//gs8S+yeBdf8+CuQJFNfccLGqPpbibWvKsb8aJ9Ugzjv2H5oRYOanlnK6htoOmACM0tAC2ui8jmyMmx8eFniUU/NM//jAmRwej8/gg+ntNA+8ZGIzB0Yn4d//+P0RP/0jsHp7ESVdfdPcOxKWLl+KTjz9Sk+Jwbyf6sgCNljAeJl98/rnlqtBe7++XvBfJsiUUzFB79ORJXLp6Le49uK8CHHuQjQetS19Bt5oJmeALyd8m7dLOFtJqzz26/l7FTTcLjY4u+Zq3n1WZWpsYXftfa88HGGCmTsnNuGFAckc424amyjUv5F028Nnrq8HA3mjqv2ey0HXZIPdaKSPPVjFfXh7Z3HgrdfodjYpv3lt7I6AaX5IZSpNT0LvDIxg/WtebJB90txqKkmE0QtGNazcnlORIhsOSA5wVPH+KB3rfQ+uuVyGX+dp+nhajRcxFIe6qAW+/KSW/uc7cPDHToHI7rgmvA66Zv9tjySxSihMyx9vZSWTjvjV2xTClEOoCEctMIAMZXPr9kEwTKrqrW4VEkhxeMzI0rHvkdVsNmubeH9DeRVf+9vUbwVTAt+VXv/5N7MNoSuQk5xixi+arZEfMzqkmNc9Ucy4TcJscvP0lNlAa+hVbgfv+0z/7p3F4ciT5l0cPH+h+0VpXIVnFoL5oUIii8N/Dz3hWvZJrEvOtszPu3r3r4nOi4dH/xriZfwt9DXo0dbrZCwEQCHmL9B+GgSUb0LZ2Wmfw74vNW/eZOXaec/YF0f6u5D/PYSEajfCrNVpxKPOF80UylinlYuSim4EqhGVzUPuAGl9mmPAazmWvU6MgkepEirPJzqMpmcygkvYBEV+/a131/CwKJ6DYZUI9pPOCghOm2hRSjw6QUhiJwaF+yePw3BXXMJ9SkoWpo7kH2vjQRUoabPhbUEAgZgJktLKyrDhpcGggthtbKuztNrZUODw9OxtfffYgVta34p///CfRaKyryTEwMhTLa5uxc3AcG1s7sbqyjZKU2Bo0LDmH8fPYgekgWVkze7oCSc8d5wNTE5J7JL6DwTE6PBwvX84Hi2BqalrPjaa81mjGqcSkNFcoOiNTRGwBa6BkUznbKCAiGyeE+8BAvJqfj9s3bsbayrKMxs+cnY2OExfzBI45yD09C+V9/bC/VIFzkSMLcfaCo3ixLzlbirpIFN69/0Bn5R5IZhjDxIQnoChBcVM4t+ecchKxw1JuVVKlPsd1ZmUDzKxYxxMUx3l2JVmID4PmLiArClzkRvgy4amwvydk/+2b1+PRw/tqFtKsWF5eiqfPX8SrhUV5cCAzB/Dr5bMXMTQwFFeuXo2nL57Fy9cLcQAIQcwh5PXMhKO4ixG5ZfjMVFeceXys3A+EPQz7YmTV2cneQDEYyYxi1VbDlFyNZ8YzogCkvSMlXewD1C/AFONIE4GmBteCXyCIc8aKvZp4cnRkSGtoloaFfKMO4/HTF9HbN6h1qH0T1mWyUdkDiSmYC/zJ/F/bWIsfffCjOHfuvL5XXkk0YiQjOjgUu/imdXaJ2c0aOzy0jFIpEyjH2m4IHMf5w5ek1vJ83t93s5e1yrnA3K74T3EjHgaYycpTokPNblD6jLcAJJ2dOh+RVxaS3sFJ3L1zL54/eyZ5rcnJKcUonGE0qa7fuK5cCmlNYqSf/vSn8eD+/ZiemVbTZXFxQfk9xTkkd1l3oIBp7nz99deS/JS0cGeH2Aic6bC7mAvkpGIlHSKzsiEGoRqdWSzm34DQdnYa0dc3KFPs3Z3DePVqUabuBmkRpB7G3h7NgpmYmBiN6ekJ5XaXb9xQ0+d/+Z//15hfohnYGSMj47GzD0AAySTLV9P8IeTRmZ956ckxr/E+X8wkcqtLFy/G4yeP9EyQiuN7xP7UNBgLYpWZ6SkB3ZhHNCcAM7x88UrxJ4yKe3fvqolEcwMpOxvg4i+xH0+ePlUOznsSa1bugbk9ufGtmzcVa6BJT75eRXHYXrCZdncorlL8NcCJecfaL0AexzrNCsbZbAqfz8wlYpaK05z/WO601ir/bi9EK49QPuu8pfI3sRkSxV/SQAV+5PMKLOJ6UYG6LFnF3lYggSb0JmWI/HnJI7kicwAAIABJREFUOgCdnxKP1fTgvbkG1nkpWhAllv9VKW+k9IH2P11LNiqKMaz9OhvABfCoeMd1HF+Z8s02sF87CLE9zvJ+5rGseJfvmYFhloEbd1Z0qBi8GhxNlkqha/I5mEkopcHmV7PgX2CqyiK/C8eUAJVihhicZ9aWt5yWRJRjHTf0eA7VJKvalZpkxHbZNBWjs5RI5O/IszVQsgA9jJ8lsDRCTUko58IGvpY3Jr/P/KS+I8+i9DeTYkdbPMZeJRCm5PA4h5DZI9/piLHBvjjaXo8//ycfRuxuRvfJUQyPjsZndx7HSuMo+sdm4rirN14tLIh51QsDS3mf5bLdmOVcdq7P3/GuWl9dE4hVDaSDgzh95owYVAXM4ZxC6YEzi+e7s78TE+MjGFzF9tpKXLtwLkYG+uLj33wWw0O98ZOffhiXb16PpeWV+Pruvbj/8HEcdxzFyPBYNBp7arjGSVdMz8zF/MKSroP8vbsLwNmJ9lEYkSeH+3H29Oz3jYrfF/5//7M/zBEY2waR4mTbRSrrI2uT6SrkImh2OojedNwZdRFddKT0LZDr/PZOvPfeezpUXr96pYOb/0C6cKAQvCD3RLBD4EJiRPBMYETBWWg06asa/UnQLg243AStZ+hkkOSeAMDBGegiJ3kcQLw3Oy2baXendTXpdJIozi8sSj9dHgaSeIICjS6cUWVF22c8ylgVanoln3Uw+0C3V0IdGHyPAosOoTD6S/THNN/24dhuxpyyKllwFZuiEE9N9FQiQZJSyabtwogReTw7Nk5YK1wzer1CKzUI+Kxp6kaFCyKnT58RyljB6cREk/ZJUl1JA8UAni+JuJ56BinMiyrqMh2E0JYHg09GF/HTiLfoj1m0LXqBKab9ovgqqT6mGeD3sKSC/xQFME2emGccAAR9MkuSJA9JGUZ3A0oSFcikdBaHDGgvG1CWxuGwGxjJmJFWKcmBdGHL/HtPyZnBblWoquKtEcOWw/JhW1+t+l3+pPkNj0t1/as49O2ykN+p0CtC5aa0l+S7hBBMjcgcJ17fZFhk80jz0NVImVo6OEqNxWwEGWliVlQT1aECTTVPKjBzgFJB3Ld2uKYWaEsKzHOg2DasP1ONmTMEE2ZktRpe0j2VdEaaBdNsODiQFiT7AhF4JbSMDc9UwYmSeAqGLvxwxVWAVFMiizymEUvjyvVGodWOHbu2BXeSZemzBAFj5nG1JJbo0RRtSVJAeIg1RuPu2CgiIfrKk6Cl8899uhGR49lW5G02KrK4IXpvs3HhC22uh/J2KNmwtsnjZddCyVTwXMUw32ZLaq4CUgU7+UCrsObr9b5fBXcV21L/k6IJ+449eNyslLyFCtoOxDVHk0ViBo/1W0lWocxOjAzHT3/4fvTEcfQLKXkQQ0P90dPXE92Dw/Hx51/F/OKKmhY7+8dxgt5wV4+o8J99+plorl1qPnSqKMq8uXTpohK0Bw/uawyZN+zJQtn3IcNBMj8Q9+8/jB9+8KP4zccfaQ8or6NmUzHNw+Vt1Ecj/FB0do1w7U05t6pJ/+014e/4PVvPpb0x6WfTJvEkLxnOqJb8VdGcYXNVsb2uQ0H9SY1zi2LP71hvmQKIUcgu4GMA62uqRFMF70RhcU65YYVcms/Xkr9rb0C07utbd93c/+s1lQC3F3jrt/geyL7zF865WYhu//CQUJ8Vi9DUBH0oXynQTSmbI3+TfCPO+qmpGSF95ROjxiyazi4Y1hqosS/PAO97NnqvBmv22CyHkDKEzN1iR3IRkmxAQoeCS/oeEQtpz8v3lKSTzkDLUTJPQDwj+cB1qfF3gCSIARIUfDhjiY/kW5JNdmIqiiHsM3vyWtmUaS+Fnp6uzpibno53bt4U8Qok8C9+9XexurGRjfkjFe5K97zYENZL9lxr7gPVqP6OA8nmk27icO/+Ookf/PjH0T80ICbH00ePYggz5TQyVlFqbSO28dpIHXoX9rvi/PkLirWYm5ZsquS4xZhg3vBcYYtSSHWhw1KGjDlrREXMOlMTnddq2H97br79ndaNFpuJ4oZMr/dAVLo4UuyjunYjw52AV+OyGoFqJmUTvhqBLj6YTSEGahZsGHczM8wapWBXRUp+Buq3EKMC4mRDhnXrRpOlPCwJ5QY+z1pCQsnKLQk7y7DAPEBaZiAWF9/En/3Tn8fDh/cNphH7+EBeFsRFnH/VXKVgXqhBGIdaS8ehwgExt4Aiw2bpTk+Oxwm6942N+OG770VjfTM+//TLeOfda7q/ienxmJyZiU+/+Do2dw8iOjHg3ZTc67u3b6poLZNuGl09PfKoODg8jnNnz8ZOYzeWl5YVC82dmotldPZpRoyPap0in7W3uy8ZmC4xHfYS4exCC4VPGob9A4Px/MVLFdEp8i0uLcW5s+dUjKUAy7pAvx9ZqJ3d7djd3o3pyclYW1+Ns2emY3+P5oHX9gmU75RqotAmfzIYfsQP6fNHTMprzVTq0suJjXslV3UQa5tb8XLxjeQkuP7+fkvAAThSkazJrhNGtAn88c7iOVxFRLNaAZN1xzu3b6tJsPRmKQ3Y2ctpsNjw2/nXurygKG7AZnnn5o14/vxpzExPx3vvvqO9f2l5OZ69fCENcIrv0xNTsbe9owLONaR2Hj6MhTdvxCMuryM393ri6lXLuAEKcvGrBeJBgo1mEY0h1pgR7p3K2bhGCtuS+k0fMv0+0kiDQ1ozzGNiM8WTGZcVa0oyNx2dlnwU+xhT5r0Ywcuhg/17LybHJ2KcuUM+MTiU2vkRz1/OSz5HLFByx/QBMRvqSA2d3b0d5ZXIGMEAYj7+6Ic/VL6FTCh3SRzHFzEHsa3WqbyO9tSQY+0b6GeJU5r1m+sbKiSbiUFzy/lvT0+nmtBcK2PzxZdfSFpqfGxcTULiFxqHw8iWyROlI56/eKFx4hwkNiU+gynBMyKuGRkbU7MEyRHAHIwhcdLc3KzONnxZ+BPZo719exP09/anzw5NVViDxE69kiMhvuIz2GNgVvDZ5P0ra6tiXZyam40xPGLSE4m9S2bu2RzhXin4szYkC9rfJ9YhMR9HanfPgAr6NPnu3Pk61tdWFfudnByKxXTx4rmYmhrTdSJHd+b8BYEg/+YXv4onT59HD425w4j+QaTdenWWek82Kls5vtZHW02DIjO+Dl3dMvm+c/eOWPbIS25sbsT5c+e0tyD9xDOEcYbkGGe6GmZqdtpzkz1kfv61PD9AY3NtSJ/x+4zjZgPVAmGVFHsRMzCG3EvNCWQRmQPlwcX1sy6R1+JMB8zJG1DDKDCG2F4HmKODxLdqg84XWLxiNWaunf4JFSNV0boVa7oe4eYaMrdmQui92sBZ7UCbyi95kQ297RtRca9Ygm1+B2qgpXeWqwfw0IRyTKCjQSr2zbO8H9dfzATl8UhYw6Zvk8wudrulE30eK87Ork6TySzGZeXpriNVQ/Ct2KHpTWX2pcC86XfXZEVmjvY2aM3v3WJa2GuyvX7gWKjZE8nYqPXpSHTrNbZEqlCsLYc14Ek/qtTjO5oVAv7I/9JAWTeSDdhpB1Q1AYjVPHDHxkCZ8h7JekSTHZNgjpZSgBvqjs3Ss7NZO/nWLVRbRmMvCd+eXp2n7IXMYxhzrAmuv5oXla9b/qsjOrpOYge/2p7uGOztjL6Tw/izP/lRbK8sxOToUAwMjsSvf3sn1vc7o3toIg46OmVgjReO4y/qIp6DXAd1QrHxiLm6u7X30ohmRio3zDnhOphlyLx3J/td4BNkUEOgvP3GZty+fkV+FXe++DKQjxkeGYoff/gjsSmmZmZibWMlPv38M7H1iIMGBvDv6Yr+gSEZbnd190pmWflRX5887JgezMGzc9PfNyr+oRTg+5//4Y3AaMOF9EJ+u5DoImklQ0UHZzXUpsSBXJRrFa2yoHPz+g0dbA8fPhSyicRBHgS9PXHhwnmZZqN7S0AKYh50jILVtkMEdBUICFFPB4fl+cDmpA2sp1uoIw6hRmPTSWxHh/WdG9vWyY+W7wKFDg513p/Dn4IGxc6dvd3mhmI0E0mq0Xw0TAgQQeFwbZLa6DLapU4BroVrkjzPzq5eR5ABDZRghBQfjTmhkdPQWHqlWQyuYrcLREbfQXNjUxfKME8t3l9HVJlxEwQTpKcmP+Oh5H3bElqMNwV9Amo+G9aFm1AUWfeU2J06faqJSlJhR9qXls2QqbRkjzb0vtaCtR6gDoMOAgWzOLhO3zt0YzZyKMqJJG87eat4WYlVoVVNxw6h/Dh4CO59znZJ85VEAwowgR/PgDl3/8H9phk2TS5QQMyjaqBYzzEkadA01D42bZrCPc0qyf5s76gbLiRISgER6Oi50PRKmTHuUwWnDjejXLhrr+q0FyQrSmhJRmhdZRFQCMhEfBQC5Js7RqFCq7hUdFHCwzIlLwSGG2mWanCR25GJEBlHlr2oAErohzQz82tan9x835RxKhk4U2hb9/LNa3WC6LnBV117oUXkW5KIEQoiJGVmc6C/6+aUklIKyaAm0IUdHlYCVe/nILyYOVmlzHtV8JMNFqH4C72X5u2F1CAo9v5BcRLWje9ExpeSMfM4VpCvxlCa2hu9w77XMggrNIjZPvjk2OS7CsN67yxOtVN8a/ycuLdMbqFkF+rQ6PkKIlsof363aYTe9iDqOZYMSatAbqSt5mw2PUp2zt/LoDYD+CZaOJE/ZmCknE9KnFAVLdQ4E8jX7TnAPOV5FtuOud5Dc6jDTQUo/FcvzMW1i+djbKA/OiS9gOHisYLBofGxePTiVTx69kpNhbXNbZmQHmFg3D8Y165el9Yv6EX2ZYq1NONoMvL55y9cUPDNukcCiiQeFDYMLBJt9kzOmstXLsdHH/+muXezt3APFA6EvhTKC63phuRHtF6z0Vr3+s3ie3uTurphDlQ95yrodzGz1TAodBmJVxPtf4Su/JiKphQKReXXfK/AnoTCng21H1UxiHEoE9liVKhYqqad/TKqCaWCaRr80Xat9VNzg8JONa7eur/fE+LU/tP++vb3qO/XHKU4gokmY838o6jEOLCWYFouLb+Jgb4BIT9BaVJALNo55wN+UrwHxVCKLzJ4VCPgQPPCiWRrX/T5YzYjD0bnUMr5eM2afl6SX2aCMHaWxpR8Sv+ACkoAK9RYSgkuAQe6usTQK9R8MTDYZ5bevHGchV8JQIr0ZgCpCgsC6rjQnvIhkiGF4hzeF1k1YiBvXcfBCQc76QfvvCt2wfjEZHz828/jBcwSFbGzKCGqvlF77aaXLemBkhs6FjLrW19pzFp7OPsbYzYxPS00OEVD+YQga3Bw4HP46EhAlINdF/0ZO66hWGIlQVWSRrUeqoggScihQbOgsnlr4Ii9lHg/Cs3VmGhJD7ph/Q9/tV7Ec65EupgExH58mcmYflZ5H7UCi3UhdHo2E+pz25tfxVxzwyLPkfSD43vVGG826QF+SJrSRTRiWRUS93azUZoyZm2SjNyNPXncJBZjUuCYZCClvjNjx3xiP6RZxPNgbnG/xIiF4qRACXKXgrMaagPso73x7NmLmJ2cjM21DXmcUcC3VNVBjAz1xwmF5cODuHbpotCCjx7cU1F8cXE1egf74tL1m/H3n3wWByecCd3x5s2KWEFgQphDW7s7ccJ50d0tNDRr5tTcqWhs7ShfoFCMTBpo+b0Da+hzDxTdd3cPYmZ6Qp4ArEHiYDUJZAS8qfu8fPlqPHr8RA1o9l2APQb8IOXTiKmpKcXOSNFcunwpFl/Pqzg4Mz0ZnV0gzvez+UsxENkhI2YpLh6mLFtzP6V5xPres08LE5PCAjmVGk0JxppfXo3VDUyGkffrFLodg3HyGM1BnTs+QyiUMmfY28SeyGJeE6ARnWrqvnP7lkzBka7kDCHnIJ4iH6gGnK4JM1oMmft7Y2piPF6/eimWyvvvvaf1xzjjp/Hy9avA2RymPPr7xwdHMk7HJ+LRsxeSgGNX6umhaOqcQM2Q9bVkkwF0aEl9FPPM7Hw35QxKsoSpQF0+NHWfMGDZd/Hy4VlKVnhvL9ZWQZf7vc1071CBHeYBklQ63/AcRGavsyOGhwZlpu2C8aQM50HdKu/YP4wnz17FyMiY2fWYoMsTqoWA5rUUzZg/CwvzAleJrTM+HrffeUd/qvHS3aP1wjxk35KkcRYCbUR9qNyGJgKNnOXlN8qJ2cc4V2iecU3kx3UecTbTCHny7ImaGpyFZ5Plgh+h5FZpsqZ0Ls9DZ2p6ARKfw7bA/4v8ZvnNcryen9c4bmxsqQnOM+/q6I6Z2alAfgvfBXLakgqiQOgY1YwDNxZgrzQ0ZhTwyLdoui8tLcWv/u7vJHeFRBt59/Xr15trdmZmRmuPnBV2v1kVJ03vDfZ9Coe7yKt19URvD14NryW1BGPjRMBC5zZdHSdx653rMrRmfjN/Tp89q7z0F3/9t3HvwaPo7O6Lrq6+6KF5Ty7MekxpMNaFC8itIrwYTOyrff1x+tSpePDwodYu7IjHT56ooUdzk30GeTie/QryopKk7FVTCDAkUnKsqWdPnypPZf0szC8kyAnwhZUDuFfWUXev/SlKPaA3gWpc2+VLlwTeoiHy/PkLmzn3GNyEeTznRF9vf6LYvb4ZV3th+eyhW0pcbpUGF1IVDwGsaCvCV/zSikkdt5ZEUuVElX86dvJaMYCnYi5L/rLfVh7Eawpt38qT8mRNoJRACQk28TN13UGxpK7XQJPm++ra098tGe4Gm1ieyr9DzEcNx/J0ym3ye46vW/n1IYy5fD9/jmP2AoW56ZbXlABJgwsyv0zm7zfj5hojg7ey7iD2ZfpKtMtBGSlpGWiFg5mLE8O3gdNaeUFbk8JBbwsn1Uw8fR/l7VkG0ZUnVw5YTIhSf3BTJnNJMaIT1FzemymzW7UxP2uzcX3mWMLSl5UabnVNeQMajwSjME6cZQLJaQ9oyXsBUsD3hmZ0gcdUI0v1kJ7eTsXmw0MD0XGwG5ODPfFPPnw3NhZfxPTEWHR09sRHn9+P/e6hiL7RAMJFzLW49EbxA3MBDykaxuxDADpcayMPHdBnk0dxLrG+aKDXPREzcq7BqGIvBIwjFmZPVwz290ZvV0dsrCzG+7dvRX9PZ3z12dcxMNAdY6MTcePW9fjFLz6KC5dPxY9+/G709nfJo+fOnfuxtbUTc6fPxjDssJ39ODyi2X0YW40d1TY5q3oBqGFOD1us+9QffUc0/w+Hxt+/4vsR+P/rCCD9xIKX5l0aoskgLAtjPtgwObXUEhs9nXw0bgk6q8vORvreu+8JBfjJJ5/E1NSkAnkCnYMjTPtGFMSA5CB4puhc0gLyndjbV4AruRbpxBt9zaFCYk8AMDDgAsH16zfi/v17KmqiG8/rYGHUgUvyT3OFYI3f44CngEWCxe9hmMNCZjOpgrEQ1IUAVJKTRmap+djT6wIGgacQK7199tPI4q/Q4mkkjiQCxYJumerZBFybL2wPKOmp/U7XWNrqyFtxoB+7o1vUfwcURpzrwEq9fd6DpBR/CX7kBsSW5CSIHmFMUKyT5E02GgisoCDzehBSmCNKZukIzdGhFtUevchDG1LZE6JD2qFch6RUjo0qN1LCiYAbDj5YQSMUOkOF67z20hcs9DnXjJHi/sFeTE1bToMvgvWtzYaerQ21jJwQFW93R3OIM3yWYglNoE6CO7N9mG88U2jPoOMI3EFqk7TxXrwPiQ73z3jVfVIU28O/oMcUfOtjG4WmeQKyulmMN+LYAYz/fBt1/PbPjPJqUUY9ZzJw/I5NocooVVQmEZNRHw1EyekYiSGJo5TW0Oe74pP0SzeXqnBXqFStEwX5brg1g78MDLW+MUJM2mcz0GjvarRds4J9NQ97m0ho08hdtNaYpTkrB3glaDVmGGzKQA9vCRDGe/tKNCuQlClfb78OYo1H22eXBrrYPH4K6QsD84SxabE8cmhcpJXXoL0HykOGgMToM7MnhIqQ7raLVUp4c90WkpexU9KZEnT63Zx/CuzSmNZzpSXz1QpeW3JMDgxLCsrIowzdmwGfkM1p1vXtCJTCmoupLcS85wPSUULkF6IpnzuFySbdOaVK+MxqoKrpksF8Fa+5rip2sBuJcZCNVf6EOiu9XBXpD2S2enSIbNRJ7O+exH/7F38SHQf7MTs2Gt3hwi8I2mG0+Pv74v/5m7+LrR3Q9SNCwlHApWFMs5JC0pdffmWEPYinvDaZUg4NxdT0jBA39+/fT7NsB8as6TeLbyQjw1q8cvWSZGdM23VzSmdcBtu8//r6phJ5EkUS265u728870Lje+/0OitKtxMYI/NUYM65XEXYkuNo3zv4O59Rr+Ez+N2jo2RCqOBRiCQ/S/YnZCTav2ot87u8RiZu2VjW88/krtmQIjnN/UJSbU10uxt3ZfBdSLR6/98Xx3yzUcG/m/Mli1JVYKbQMDY2rKXB82MvV7FbrCZL/YCA5vmytiSH0mufqDpfMNy8euWyPJqWlpYDmRONJ9KBJaFRzdvU0/VW2VqP9ewYA5IRn7KpFZ1sIj0f7/ja6yiI4ZlDjEBRygCFUX0mMpM0yRgv9kc0cVmvFECLXaX9EdmxwwOhi7k/GhUgeWEnCdWuhmWiGaUljXTenhKwxkYjpiZH48fvvadGxfDIWDx68jQePXsae8xpSSGW75SRoW6S+5jgmZTXgYoRetrfTm1k3K6CPWen4z/uYXxqKrqRskF7OGXl0O1VU+3Ycw82Z9moMBbVmJA0zZFlI0rDuOQbqnjJ2S86f8pCcdEVp3F2WuJkx3tdFg3aZQF/3xxtBxkICDOEVIYTbzf4XdBgOARSacpN2G+HmErAmiyocu28vMxDa75zz0q0U9eZa3JTxEUfNfiPDqXNTqPNGuGsQwNBys+C8SJW8nmeaNDmDZ4o/uEZEcMRI9E8qbXL/sNYbtPE6+mWPj/XS5GWfYLrkw70wWFMz0ypkCWZzX384EAm7sTjJw9jam4qnj9/FqcmZ+MwNaOR4CFg3dvbjv2dRsyOjcQEDaaT47h17UJsb61pPnf39MfhSVc0DiK+vP8kVja3Y32rESB//ugnP4zXL56o0AZzbv/wKPZPTuL14opQ1adPnYm1lTWBSigKSvZnY13FURoTsMpoVFBvGx0dEDCKQsLS4pLkXYnvmMOTkxNqVMCeoIiAdA/7PYCiudkZje/q+kZcunBefkfIxBIDLM3Px8zMZPQPdEdfX3eCofDOO4ljtKO7WJeWvKWQTVxBPCBvHGJHnesu4DGuFLaZJ+wV63gp4Ofx1QMZh8ucWywNv15rTzEohTozyiigw6qCgcEc6uulgMOcwDuK5wby3BIuNPS5B9Y3ckpc4+jIWHPN2AQa/4+tmJuZiY31tXjx/JmkZqamp1SsWd1Y03jwDDjLKTifPXU2NrY2hSxf20L+gkbIbrOhyxlcDU3FBJiSYmaea6kQzfybu2Wus+7VhAE9SwF7B+aGvTTMroCZZhlfciYK7XW2VEOP84JCMGeGYphmYc376djoiFgvk2PjAauDdQXggfy0sb0Tr14vqRAkeVzFSJ2OGcjLBGrxXkgePP/qVWzvNgRS4Xv4Uvz0Jz8Voltm5RkHED9ULk2OBIuducv3nz19pntnLpIL00i8du2qPCK4J9YzrBful2tamJ/XfdGkZaxu3b7t2KOzU3G14mQAWfKwsswpkmI0vWhUcSbCLCIn/vrOnXjw8LnOX88Znw2YP5ND/vznP4vzZ89pDAW0S2ll9hX8xTj3WrEfHoMb8kocn5xQ7o+fw/MXz+R1wn7JWqDg/7Of/TybP95biLXYaMnpmResmwcPH6k5efb8OZ1j5LiwDpkP6+R1m5vx8uWreAyTD78FgB3DfWJWXLh4XlJ05A0YbJMr/V//51/FvQePY2cXUEGX2H/4/VGcFKMiZWO1VgS0s38Hz5xzHLbE4vIbNX+RucJ/g3snHmU9+Fw6iQf37yl3kFfO8aFMsokT+P07X38ds9Mz+vvS4hs9Nxp7KEG4nmCgJHUSmtOOHyw9yHqXHPMxef3puHrlSvzyP/7SDO9stPM65iuND95PnjWHeHwZeAOTyM0PN1A54Jj/jCnfo+nB70t2LCWElbelNCM5GecYZyW/W0xRxUnpnSIMep5RlrRunfkqQuOnkHmc10T5mbXYlI5PUrUgz12fowbS1s9dw3ehv9QdyucGmcnabxhD/VznsJlRJatcMV675K2kieRZaTWPt6W5nS/bt7AkiEvWOSWlUupIzYCM36rhIsZCngVu9Nh02nF/Av4EYjUQUjlgetW0KxoovzCCrDUeTigUtzQZFQpxK6armoQDhwJButFTpuDNEkKznmGGhZsMlsey5KHrWa5p8V61z1e9TnNX8459vVP1IceOmdsqR2oB5bj2yi8MbAE4hp9Ph+Jbfo8zk3OB+Ub9jv2t5EyV0yRDpLOLhueumPe7m2tx9dxM/KP3b8byqycxMzkexx1d8elXj2Kno19m2lu7B8rOF5eWtVd6WDuCBrDAiz2WgDf79iRosiI9zuerRsjZPjQYG0hRJyCIBiW/S/1sLz28JifGo7vjOJYW5uPDD96LzjiOB3fu6L7Pnr4QP3j/3fg3/9v/Ef0DSPQdxF/+iz+PU6dPSxLz448/jt/+9kEMjw3GtRs34vHjZzE6OoVIf2xsNOwPSV2OZnJ3x/eNit+fAHz/0z/EEZjcs56hO8je0ChIawNKuRMXTW3MKn3m1GplUyGwQbLh/fffV1Dy4P4DHeIVoNFNJElicxNKdW9PSTQIjiZ6/PAoLly8qMDszZtlvGGENiEAo6Dswg3Ur3EZdEHblhbowUG8nn+dBxFSCcgIuQiBZjIasSQ5fJ05cyaWV1bUjd7d3zXKvSuplpKMMCqfe5L5bF+/kj4VPSgWhXXvdFDUoSANvyPJmhAgsJkRfLKZD4+MxOv5RX02zRtpXUcIWaEkVYfsgZJLNRQY40RuVpFFmzvNCvT3kqZaBRDeg+QsrknYAAAgAElEQVSHZ8FBwEZpZgOJ2aTGuQzVOGRAni4tLQpNxH0xvhzaNtsi4Abp40YEaBQ2/6JYtyfWHE7MA5mdJ62zHWHxTesFIaVSEkYbf+pim8o3Gvv7uzE2bkNDTgmemZofiQCrGrkQ93moYvLH/VMMUTFDCR6GfrsKyjlYVISLExc0EjGjogyyIwMDQgAxPminyiw7G1WgrziQSBKNvnfBgedDMdvBkgOl/5xGRQU7RQl0UbANIv27Ng3paHbK0JBmW9NEMX0BZDRPA5GflVFu+ny4AG+0mtApIBoyGCqUa/Njs0jdXohkDbRQFaYJVwGv/XJLCs5FFxfGmsWllHByUE4T1OuyCtt8nyCE65QWJaboUOzTAJ45u7uzFx2wL7QPtYI4f44LuGoEyagri7h+QjnGDuAUFBVaR8wUmgTlo2Gpo5KQchHPBehC1RTduNB+BIoKoFOKrVC9CvJTBo9GhYpPJYSeQaPnjP8r34gqnlVzynOkVUytYpl0UL+xwKowzji0ywk5EWgxOxR+5Vz2HM5GRY5PzdMqTlqz33O1gnteo8/hvXRf9muRxMxxi0pvuYOD6JSeaMSRjI5P4l/9xc9ie3UlTo1NRB/Ff5pMoN2GhuK3X92Npy8Xoq9vyHrOx6AR92JgEO3pQaHTvvzya6GCSfK4NzWX0QDdJkDrjqvXriqg/vruXUkisI/MnTolhDdIYtbA9PRkPHr0UNIJzAwVBZvG6yf6PZrwz5+/FAOI/VmyCemTwBzgc+ur5nfNbckndXUKaQMrrRiK1TTwc1AqkrJDJHAuHnt/QnqCZpl9GGpOFRNCzLAuiuBG3tceVOvXiahRyvVVKDczAzLhS+uV0uXXPptzwc2qtwvX/zmNippX7ftie6OivYhLo+L0qRk1tpkrnEFcH3sCSE/2BO3LQupjbr9heRjJr/hMZIzsIYUcx2LTYFuJotCCnqfqlbdR9fl+rakac76nMcZjL5taDIF1kXP/EHLX4AviEpL3QqVxJup65GnhMWavRXKG88jsMhJYJze8D8+Wuc1eQcHVhXdznWgwimWKbxJMhUDekYJQv+Rwzp+ZjZtXrirb6+rpjeXV1fj8669dhAFFTMMVz4s9ZDGL0eB9uvY44wjyPPoOj4pqfhuAwVjvqdAxc+pUbOsMtmcI0kHaNyj+dHUJ7czZrDmdxXliJyXSeR5ZyqjVnK0ml1gl7Bdpes18Re/XoAj7hbCvAljQe1CgybX5XWfUt4/XVrvbDRQjuEmqJT2aMZ4YYmritM4OgUL29yWLUmeeCxpZdMjkW02LZKZJuz/PJstQFhrUBZ+JiXHFjpLTSyNMNcClYQ6jiqJTmdr7cwqBqSJHjguN15LnAmlb57EMnbPJbz8xinMuevlzMDm/GM+eP9fnE6MXi5SxYV5NnZpQ8XV7YysmR8c15iTnewe7sbqyFKND/XG8sx3nZqai+/Awzs6NxchgjwrYgyPjcdTRF1/eexr3ny3EYWd3HGTecOvG5VhefKWzd/+4M5ZW1mLm1FysbGxKk35majr2d8yKYN7hNYGkzNZuI0ZHBhSHLi9junwSExNjijPJPTD/ZX+gMAgzYHtrO8ZGxyW5QmwPQ8PP3dJXNDJevZ6XTA1jCBLy4vnz0djcpO0pDXwkJfAcgCV9fMw6zeKKzuMym/U6Yc6TQ5UPFiAHeQ2lvrbM6ym+9/fGm9W1WFwEbGW0rxsV5ctjvS2KIhQgeA/JEvb2NfXBuQdiY9Ya+Q+fz1hR/OVM5HkSZ29uNszowNh7zwUf7UNxEhfPgeLvjefPnqq4evHihehCVvX4SICmVy9fxf7OXmxvNeInH3wo8NDjp48DdXk8VUDqM7btsUnFD8WYZVzZP3St3V0aY/Z6z1mfNexTPAv2ytVVZIRc2FKD8OAopiZ5hgMxP7/YZACJVZFMIoBoyOMQFCCZ4TjR7DQYOICiZibxTSCGAI2PhwESZ/vx6tVSs0EBo5PrtoSowTs0KqyP3hGvXr5M9kgyLg4PZRj9wx+8r7OqPNW2dxoqZksSDM+xDory2/aRattXkEriPPnggw/eiivEiADJ3uXxIoaBCQQ47+q1a8qB3dyxXjyNChhQzKNib25tuUkhP78EZtCs++yzz8WSwiCWJhZgNIBj3POf/vznaqYwj3heMB/kqXR4EEeYeyd7/vPPv5AMCU+P5jFNBeYR+eX4hJkSNO4BycEcIYbjM9ibPKY2oOYZ8sxpxqxtbMb6ekM5PnHX1RtXtEdSH2BNkRMwN+58fVfm2ccy6qWJdxzvvnM7rl27LLATCAjAK53dvfHxR7+Nz7/4OtbWt2JwaCS6+waiu8dNJcU9Oc/YGwFLlQcW846aw+r6qvIvrv/163nNPZ73ixfPJU9Hc/Tx48c6E8RAOTkWMIFYgHrFk4cPNc8wgl+cX9J5MzQ0IlYZEm1c09Y2LCCvA54HZx51BT6L/WJ0yMxT9PBpbgE6dFPBhXh+VaTylMm0XCNodMejnJGc4+whTZZ6p8F7blS52O4YpcX8ZT+pfMiSXWaqJf6wueZZG9WsVywl0Bcm2QXKK7moFji06krtcWzlLQINtPl6NhsVzQaH319gAOS8UvZNoIE8Y6khSD45mxra81IJo6R6xWquIkMVzFO6s+6xrs/xq8/vyuNb+Z337IrvLW3V8uSo5oSBQslIasphOY8qRloxNxxPN3GRzfhcfJm2ZkXzQ6vX7UBLe4dLei3viWqiVIzOnq21+A0VAkt4m3XiGNfv0YyFm7Uq5yn8jPcqvz/Wks2p3fAz2KItH643y92/nreBgW5UqG6UNReBfHUO2nPN8Sg1N3uecT/s6fidwnCkEdBYXYsfv3Mx3r9+Id68eBxn5mbE5vzoiwexftAVPcOT0dM/JCbF64UFqWYQj+/t8xw7tN9Sg4TNLCm4bhqup2N1ZUX7Heuv2G+cO+zzyEidO3tG5xrNTYAv+CkO9AGM241GYyN+/MH7sb+zHQ/u3VOMOTM1G9evXIu//n9/GSMwB7c24l/+q79Qnjo1OxXXb12NFy9fxMPHSDE2lJeurDail1y5s0ds7arLarp8z6j4dtj//Xf+sEdgXGZM7gBzuFXRuqiRBLYcTi6AONGVsWvS00Gug5RACxaUCIV4dUO7utSBX1haUIBWskFK/Dkw+5B7gu486UB0/yAePngkmtSm6NCmfvEaklU6qmdOn9GCBVHExkXSwWZAcduajNbBZw8kWCtEmVARiwS3TsT6+3v1exRPFdRl48UI2Jbea23mkmbqTjkgXVNXFkiN2rW2d5co5CQFBGqvX72O7V2zBqpIwcaGTiVfBDEEhyQCKrzgxyCTT58GRdst9H0V2cvAW2ia7i4lJxRMVpZXpHXH4U6wJMOszU3dI+OCjioGl9YAtbwJ90rDqEyrVCxOlE51wFX0l5YxXiY+QIr6S+JB0C2tU5lwGeVgarmLPDzDarx8U0aKjZ9nQQKBNqqeN8l00nFl4iTUWk82ZSzDsX90oCBYRW0huntcHNnZsWE7jZSkvaKv3NS2PDDyjEQCum6ZuHIYNpHGzM1+gm8XqEzdM6KaomUhQ9B1rwCmAkzvBIVeyD+z+FQan63A5rv3jRpb3luBc+qcE2wxxhTxGF8FmArSU6okjd5dCHKhpD6rkBxCuYuBIMyYA5FsmphN6shGa64ZlHyDqtl+2cnycXDmwrvGOpEaDoJaHhUEPzJlJmnLIhcoHhW7Kfo1dZk93/waB7hcrgs0WexK5KsDzRY9V3IJeY2FnG4iWUT1bS9UtSOMc8xg8SQzqgqehRAyo+FISLwK3lxUQ07CzBs+v1gZRkG6kFWsimpUVOGXe1PRJI0zHeQ7mK37bTaevoGodePBCH5JW5WUT6GDyyg5R6QCOs3XYgNlUtG0OGsL5E0Gsc9IJScUAarpVUGrpeUsm6NGGL4/ILiRguhipRxHT+dx/Hf/4k9ja3kpzs7MRccJchgRY3NnpdX9tx/9VujMk2O8Qnqjp9em8xQQQRcii/Hw0WP70pArlBQe0iGNba0Hzq5333tXzAvWBpq9zAWK3jQfxidG4/joIBaXFpqeO4VqglUFAob9GYkBCgLyTtrGLHdQ41sGn0IGZUIkllsaVVYRmOfGeYmkgpIbD1SzkdRO9ZbhvGj1JHUE4G5Ks5bYb7Rv1JrK96FYwt5bc6W563RYi54v9r8msy2lQpqMj+YayD0q9+1ax94f6svXXY0+z992pFZ7JvX2ntZqDr7t0aP3ODmJuZlJFVjUlNy1bnclxchbiLVyeKxxJ4HY3t2ODhVbKQY56YE9xxcNZ1CdxARKVPMSy0/KaK66q2T9pcSlG7NG4pHYMudYc0Ldpo6/5glmtDQO+lxENhK/pEc6lahULMW5Veufzy7UaiHYeF8VNSlGdXao2eZ4J4uUKS0gzxEhtWCK0VTrir2dvbh47lTcvn499vesjcvV/erXv5bEmRWeOSNAXxdTNM+zNgQdb+yGJfSz1hPXPEg0Xxl8V5NUsdjEBBPWYwU1n+vOOcS7IE8idFf6I/EwZAOce3fNdctAmXXp5g0GwSnhBOIwzzHODJqJbrx7jvk5W6aTWE7v+U2UxHcesa37rDN0YnyiTTPdxWbiRD6rEniKHJ4bZv3wp/yVknVTa1H7QiKqq8hTzw9EfDXAqxDA2AOaQJaO1/kWDEKBWazCp3xmbPCtPaLpG2XvD17Deq9mBQk7wyT0OmajAAWSHSgE8MlxzM7MaNx5P5oWX3zxhVioNTpcH0XjvoG+6B3qVbHyaHdfDebR4VHtlaD/8D3risPoPTmOMYyUz5+Jw+3lmJ0eic6uvujqHYrljZ346Lf3Y3PvWD5Eb1ZX4vY7t+L4eD+WFl8p2T6M7lh4sxqXr16J7b39ePniZUxOTsfO1raeNQ3qyanJeDX/2qCliRGdd6x7o8UHxS6BVVH7Hs9Hc4K4o8tGsrwXTS6ANrC8AVkRAyvWEBhqzMa/3d3yNkBedlIa+JZgQm4Ohl9np9lbAFzk6wMgI4spYkQn01rsVdh6fWapiy3OM2W+93ZRhY6nT17IoFusyA5yMK95AzdKmsbFGfYX4nTQ73pNMhplMN9hyZ/Srq+zQya9yFW1gRWQMaJ5SExz5eIFIdSJeQFVXbl8OTD/rrgXuRp8gDZWNwLTe5gtz168iANJVHa7mZ8Sidwj85l8i1hV/lXpL8gYw9ZgL0e338wqYgQz+pivsN85e3kGzYZqImaRbbXXyqLlntJjsNjS5Fqr62sGjSWwy2vAHiYgYWenpmJqciIbSgbfccYvL2/Ia8EqOI5Tfd2w32BWHCimETNicTHIK3g2MNd51kLxX7wQt2/dEpuFRhH7BKh2JC5hZ5AHCyQDIpnm6D6o3P2m5C9NIsncilVv4Bz7G0h7xv/+/QdCC7969VqfR67JXGLMbt66GVuNzeY89N7bpfnt2KwzxsdhrtvrjsYFUmiMu0FY+/KK4PmfP3de+ZiKunleSM8eVPzRnvYSYgLYD0gf4fsyPTsbn3/2udYQ1zI9M6M9VdLCabzLHifD+80tmXP760TPhfOPvejLr+7ExNSMgH6fffFF9PV3xwcffqBr5z7F5j80Q/HTj38ribGOjkN5yMD2uH7tkphRPFfGcWRsIgaGRuKTTz+Pv/mb/xg9vf2x2diN8YmpZKQYXIDnodh1jL3kmHb0LGgGLa28UaOCuf9IMWhvXLxwXj4sPGPAf7B5Xs+/UmNqdX1dzC/iRuohTx4/kk8HfhcwKjjnyF2X3qzE2pr9LBu7lrcuJi6KFKXQwDgST5L/uTjbEcsrbzKvTU8xnonFPZvgDBV2MbjvN7CQn/I8iB05T2pPcljpInNJ1lZuS07DF7m689zyXjLQstah0eRuorcajAZWVbGc9zGIwobd1ZRo5jGVkzgZbfqWGHHv3yhgiM7RUiqQB6K7NK3c1Xkjv0djtHwy+GaBjoo93p77Ki9rSxOrh2H2Z0lYOW80+p/IxzGM4/+2fCyvu0ANVWfhPioWb4GIMm9/K752Xl17a+V3GopiBifASIMj5En++R2NCl0ZYLNkcpSHh2NWx9MFyqznLEBd5qOO5wukWQAONzPYI6vBUnNCNcTyN1G+zi8bpFVfkjDUnPH5VzLwVfcpOSWdo9ozkd+zRDfND2JuAyELTAkYlv7+QRxsb8Yf//h2XJqbiI2l1zE7NRmN3YP47O6TOOgejpOeoTjq6FYDd2u7of2Se2CP0Wel9wljAXCORilNV8y03Rg4FLCN+qU88iQrexQTk1Pa0xgTDhQAe+TB5AqHh7tx7drF2NtpxIN796O3qztmaVRcvRF/9e//2jKax0fxr//1v4pf/M3fxPLqWly4NBPXblyNmbmZeD3/Ju4/eBivXq9qvxocHBFLlAYJDReYYt83Kr4z8P/+m3/IIzBzcGwJnSwYcDiLdgtyNA3NiiZuE1U2FOsOslD/0U//kYLjJ0+fip4tE76dXSUM9+7dixMJ6p0oqHIC0WEUOPIOff1KDEBrfPrpb4WGovOvpCgPbQoDFDBOnzkVT588VfA7PT0TiwsLopxyeEP7baK283Qq6vytWzfj6dNn3sNlVocJVX8TbcCm5OTtxIWozg4X/79xoCqpBcXOZso1JZKd4I3gxuaVh9IOffrkieSGCMp1XcdsqqZZUhyHscA9EbiR8JnSb6RlIYSqEKbGEc2dYwILIxpkYptG1ehmohfLmFXhg+dF0AtahXui0Ccj4sNDoVPKaNV0bEsalFEwY6OiGsWuXWsjqzmVaATkXfgcEmDej//4N3+KOkqClkVTAhJLQ0H/tmQH925ZGQc8PHvYC8y7QoZVQUn68RTfZCrar3tRp1168tsxMDgQSE6IEnh0pPslyeF6tneNUFRil0ZHvhcaKTbeguLP+0Ilp/hKwdOeJMxNmgRG+tazK8RN3bOpmRS4yyzMAVUFuyWDU4UY/5kNgjLpzaLQW3tIRkduNLgwKM3clPCoBoQRDE7yVDjJeaziEhqmMnnPwOUbm1QxK5So6Hm58SLmBwi1/n7NmaJzKkhUsNYKZpu02/zcQo9L77Wp8e0CVTUDXaSyvBvPl/Gm2ChEhBpoDmaMCEv/i7bmQjPAKSPvkuQSPdXPo5BorQCrVfz/9l7dxoxpjrZKeEaqlflaziXuzXOauZ6SPVlQVVEI5k9KifD5or/muFUs2UKntILpVhHVtTgH++0hXYX2DhBZoyqENeWGXOiTPBFrMtFRzZAwuz2OZTEdIxAzwqik5kpGxXulg9dKPsz+cMLEs+P9haRBiidN1YqNwJ7OGUG5DFr+bmMtbl+/EHNTY3Gyvx9n507Hzi5o9IEYmpiK//DLX8beEfKDA9HbbRkx1rQKyBhoQv+fnIxf/+YjSeVkNK5rEOqYogqF4b0DNSrYB5D1ELKuw4UT3m9yaiJW1lbi5YsXOqtI4jmLJPOQyYwYgsg/qLjkYgFJ8cUrV+SP02CvIXmTrJmeaK6LzjjheWfjiiAS5GPtyRW0f1esIMaT9PfNDjLDyHR9ChZZYdIzt7k3jT2SUEzcKZKVRwwyEDR7jmNb/j5e05WY/JfEKU2EVCKylBgmBdztzVbRX43CLMBYdgkptcOU2MBIeuUthoMMHTs7YnZmqkkbNyLOKCm+zKKyJCVjzDNcXlvVXNBZTLGuv1/7PT+3rMuQxqw98apmpZNEJ30av9xf1LjVPCtzSZ+T3BNzgTFm7lSiS4GnGDVIiRADqcna4QZbU/c3jBL1+X/cvK9qTCpZzeSQ4kLtDUbgW8ucguAJLBIQwmLQOZlkbM/MTsYHP3hfDXtiEcxHf/3xpzLpZQ6VXID25GTUuTheTSYn254b3m8MNnAxrdkgZx1gHn7iexgaGIzO3u4YHMHvoKGiFfs476PmMn/Kawvkt1G4anI0GXGtJmM1j9zk7owOxR1mWjCmyjjTG2hgcMgM3ATVAPKoM4X7kLE0vJMyrc6m9NsNNu+dVYRRoaG7K6DlMz9YczJ2HxxSXCaWZZ6hTY+iHEL2dNZ2MXOq+JA1luyAp/SZ9t5CUdqeSGzWzi7tNcSEmo8pZcGeTsGL5NPymDTtjy1/lp9p8IXlOuqzGQ95PG3BOBjWGlFzRchG/GnMbmUFUKRCxmBxcSlOnzmt9/ns8881JwEHwC5gXg0MggY/iD3iKc6L4+MYHh5VzD9MMbOrI7Y31mMQIM92I/7oh+9GY+11DPUjszKu/168Woo7959FV/9wnLlwKT794vO4cu1KrLIXv5qPsxfOxUlXf9y9/ySuX7sc65uNePHiZVy+dFlgG9hGFPzGJ8eFQGZNse+PjI1qj0dOpxDBZ86cMhgJabXUt2aiF9MMZtbONszbhhoCOkP2duXJMTTYL6TypcuX48WzZzE00B9zs9OxubmuPl4xqcS0zeKUij2wDIX+JBb2WkYSjuInL8MvR0zLNKRFgoc9ZWxyInZ292RKPzo6Hm+WV+U3I0bLwVHuHxRoQub0iqlgOqKRvb1tBjlSGAP9yuFU1BZ4xeAg2LjyL8D4fHDIzENiylwDGI4y586dORNPnz5x4f/4IC5eOBcXLl3SzziPGZOF1/NiuyPLyB789MXLWF7dxOa7WcBjewEFjtkwps72Z+iUpBfMH+5jdnZOYz4/b2Q6MYgbSkbZg1onL2IOM/+4Vs4TZHLGx0aU13CeWGPf+yHr0KhgF9rwCRIghr2rH+nA0JnNXjoxOhaz05MaK+TFMIJgTmxs0Sjuiq30crD5cMnQWIKLvYyxhgFB0UmMGXmuWT4P/4szZ8/Ehx/8WFJpyDjxLGHCTUyOiywDQ5T4BIYP48sc5bkQM7E183obMuOncCLpD2KHxTdL8eTRY4HZMKFnLMhhaJIhk3nj1o1EGSOxwjiwZ3do7tFQ4Xobm1uxsIR/yZaMW9nTMV7H72iCPLy/TzKZM1Mz8fT5M40hbKfefppieOCQ/x7E+bNnJX1IXPTy5YvY2WmoWAZIDC+Ky1euqKjHHF9YXNDzowlC3EUjhL0VmWjYBjIc7+6ORw8fGaTQEZJhe+fdd+Prr7/Ss0QN4ebtmzrf8dHgdXt7B3Hnzh01bzCTxVfizNxsrC7Nx8WzZ+Ld27eEsObMGxmdiPHZU/Hpp5/Gr/7u17GxuR0DQ/g5HgTniiRwTgos4XmkZjGMkt5eSXYdd0bMzHhuCmQxO6eYA0Q0eT7NjcFB4tDOePHyZTR2dnV+qyEhtmev6hswTFibzG2aFJyh+NewHxM/ih0AkG7CcsiK5bNByfPmi2Yr65yzSiwrvaY783qD+vjijCRH5my1VFRJzLbOQH6XM6zO8AJsVN5HrFZMi4odiPsFnGj+DDa1gaMGmDofFatC3oiOa93EL5BcMhBSHdr5pQF4ha7XTWRDoD5bjQTj+5txd8V0UusAfDkIGNF1LQHbWJv9Zp0pRjlO1qxikrcBGo7oW42R9pi5gFlvx9HeIyqnq3yg1Dma3ZJmGt6Km8v7geuq5kk1V8SsTYZHxSsGFTo3qzoQa6v8Aa0ukMxsmpNteXPtZQZMWubSDSOPo6Tc0jtD+1mGiRXjVEOF8W0CIZNtU8+uYlg+q+YGZw9fBU5BXpX/FQil6aOYShEGYdgjQudUMkaJSyQPnTKBjAHPW55HCQYgN+pkT97djLHh3vjv/+WfR+dBQxJQR7u7MdA/FEfRFb/57Vdx3D0QHb0D0dU/FAvLq7G51VDDHXl5wMOc0QIaJXCR8394bKRZD2JdUFdT3S2VNyQlnB6pAAPwGBSoUWA2ZMP2YnNtJX7+8z+OlcWleHT/YXR3dsfFC5fF/vzVf/xVgnqP4n/8n/6H+Ku/+r/V8N7dO4grV8/F7du3dL+jU1PxyW8+iq++vBNbm/tx7eaVGBybEBPk8PDk+0bFf0mi+/1r/zBGYHwbxLkNPNksCfKNzHIhQOgOEGSSZrHmK2ZWFJUxMAXhAtJVyKxTp2TOZbPJhjYV6OFQUsvkEyiRCtpQKedOKdj+4ssvhJgFvaGF3w2izR4KaLAiK/X02VMZa7NhPnnyRBTaQk0QaFCAJ4ggQCo0OMUtaXUXgoUmyI61MSsAtFZrOOFPiSXLwhQa3AUMgjQVWISCLMkCAnNrzxIoEFAhqUTwNzw6pG6r9VVtdEdSYuMwIwugbPGZUMsITFs0O9N9eQYKyIVMNs1Y1DcC3L39GJ8Yd2f38LBZFGHTZvwYBw4BBTWJ7GbMB4eHsqlgup8Pik4nsHkwKljpImhvRCdBVRYaeDZGilkWB61ejHB1mCFXUUlQHnKW1LF0lgrRJJhouJZONgHSENq6lpRgTvEaAmZn3xGjY8NKAEoOhASikJMEa2urqwpcCPYpWglRlojHQrEWosjNHaMTJXXV26s5jDxYSR4YpWU6urwhDo8s9yCjcky1fZAS5BZzSKwjac1bA9PPywWEklpxve/bjYpv7hIqo6XqT8sM2RqmBH3WtjTdt0IeEgqCVsV1J/aT4VpsFvZ2sbtZpkoJDlC3vjQHs3V/BAl6zoUYyQsteY1CszDGLmpZVkLojwyYuC6aP06u85GqiG/EmEwC87qZQy6IQbE3WkJJd8pvfHOcXLRq1d2qCKBnncFYBT2m4bJ+WkW6t9/v28Gqf+65ItppGh57NBOdnAZ8lqMxI0WMp/w8N0rels0qdFGhi5vkBgpJao94hBX8fsezk1ZmNkKE5mVtNxshbQOS72H0uhsv/krJqjQJz4fvglciZlQwy8YXCVU1P2C7KaDWHtitvWNnf09ozZIiQ2dZBQSM5aRcsReHe5tx+9rFGOztjDF0fbthUUWMT83FZ1/fj7//+LdCafO5NH7HJyZcVEPbus8MsP7Bwbh/736MTYxrfEWzzjkAk0008AzM//Iv/zJ+85vfqIhFsUSI4+1tscpeL8zHyuqyGxQnIRmXQ0wNU54O1C7rnaegRPHoWGjlS1evxvIg9kAAABsASURBVL3792OjsSkvIX5XxUvCUPYMGpblqZNsQs4jo8VaerTfGRVkw8P7r/Vd+bOMyctLxQmKqdhqlrYh2VUey6YTfzZ2to3GStp7e9LyD0cmFKfN5jLDrpqrTvq+tWdpirlwCwNCiNTuLhVCmVM0jZQMUThN01+kJWamp7SXwoTg+RBDaC/LZgWNCu6V580ZiUQC12NJA2vGgyQmIeCssl8MiKtWQlPr2GNrplgxRMxucHGe5UaRgWRH953IShJwzf9ccyQw3AOsT5iArIlK8ApNx2cV2q4YqqB227/qJFCs0Satxzi6+GBgwt5eQ2b0IEy1t+C9tdWI2emJeP/2TRVDZTzd0xeffXEn5peWzJjMhFbHqOQK2hpLuQ/UHsT18nmlRcw5Uwi7moOOU3bcBKLADxo8WRRuhtCw9/8onjGeXFczsVS6lnMniw0lGamiQzYqqgmrs1VmomgOW35NMQfN8zwj3KT3eWMkoUe4kmLfe/rGNNGarSKNnl021JHT4dykMOazLw3XM5jUOuYeSgYsWYlNHWvXKpoISM8pQCxuBivRF7tSp0eTeVNFIjW8MlaSnnaCPVgbhdr2vPceXCxVyX6U51XJEdJI78MrIWUjU2qFNUIDBBBGgQCIkZ89ex7//M//WTx8+CjlG1w4ccEc77jxWJyfj7GhwVh5s2wWNOsC9Pz4eGyurcq48rCxEe/duBznT03E3a8/j6npuZiYmo2nz17H8xcLcdzZE+cuXoqJmelYWFqKlwuvhXYlle/sodjuotz62mauH4pvO5JNwdSSPYxCr+P0XknFoiXNz2hWUCzltVpPKRcp7Xm70KeR7Ens7dv3oNHYUdFd+/3xSZw+PSezW5o89kLZjLOnKax3yiuH84S9UB4U3WZ/VVMQfXg08ylmM2XE5h4ZdMMqdd8poKkYzXnT3SMU5/QsxtNbQk4iB4exbifN02LzCuxjLzB5fB0dqgnDuhJbINnA8kdArgjwSndXk8UNMw1wFuNIU1GeDKDsj0/ivXdux8bmupqPAL/IQTBJn5odj3du3lYg2hX/X3tn+hvXeV7xhzPkLNxXiZRMiaRkx7Hd2HWBIm6aFg2CFi2KtI0RoH9nky7px6JFtMSpHcdybYuUKIqSSIoUxXW4qvid87wzY9ku0I8tTMAW15l73/suz3KWqu6dPXwVeYv+wag1GrH80DIUyHhZohDwDzlFNWavzCoHUuwnMIXb2qwDirUwIygwO4dwkVT68WIJjGY+c5jSZDTebRJf0Ljetw0ucyHLUrFaX13MOc6F0zQk13UcH8fk6Fg0FEeHEPqc2wdHR/Ho8Vr09w9q/yCvYT8qsoIChSTohIMfGSPYFaBktd9k85Bnzt49NTUpOSD+k28JjeTeHuWE7DMuqBoERBPjtOXmEmcLjRgaQ8gCkftSuCdnswRnRTJ7vXgatA6V81Z6K7F7sBvP9/bi2rXrMT42HkQl52eYv3r+HcMuZ+LRVDw8jN99/Lu4t/LQ0paHBzExNqY4CK+Ss+MTKQMwvjdu3Y6Nzc0YGRuTOoCauUdHMTw0kCCjXjE8eI3dvVb86M9+GG+++Zb20Fp6UMI8weeG+UPDROMyMaWcQDGYZM6I8ytiGzx4uBxrG0+1jp9tb0vu7fq166pJ0NxhzGBAERswJ27/+tdxf2VFzIox5JUuTsXm2pOoV6vx7u+/bS+y03PJFdaa/fFfn30eN27diu0dpJZ6oonx7el5VDGDT08Z2EYGLDal5PBwdSX6GnUBL2DmwsrHUHvp7qKYFJOTE2r0jY8Nx8LCguSokdwCqc18X/zirvbM6YvTarKV2F55fIIVjsnpJLcaykfZ35jn+veMpiVnr+sIAO/kG4GXgorc7DnOCxXPZO5ATEXjutQOiG0KIKo02LsL0WaxF8BGMlATuc86Jb/jbOK9rcpg9mE5cy2lBditR+BDAy+deaiAnhLK8uNJNqdjpw6AoLAtyn6hODulkjLEbYdRRW1D9YSUJ6Kx49wgFQUyRyhNXuXnmT90gIAvZ4POo0qx3u/7co745TjYsXkyOFJO08DcPAJK9pUv083U+FL8lWbg2oeMvGs3JspYF+aGmfyWxGQvNXDQUl+lmVByvnI/BTSoOhaynCgEpBesGO1pYu7GhudX5zVejvydqxd51bZcVAIVBbLyCOR+50a7vpNy8p4jKS+dTA9GVnkZ/rTJYKXu5XzuSGuJD2o2YkFT82J/Vk7UE81aT5we7sb0RD3mLk/GEM3qM2pJeC/1xAe/vRM9fXXFHCd0j/tqce/+gzg5tpQ06woGF3GCvBxTVrl/sClJNpRJlB/UkIZ3HUl1Rf1rcBJjR7zVV8Hz9SRGh1E7OYqNJ5vxF3/+/djaeBr3F+9FNXpj7sq8mp03b95IwPh5vP+z9+OXv/xX1QtbreO4fn1OdVXOzffe+8OYmZ2Ng+fP47PPPo3PFx9GbXAgpi9djnhR+bZR8fI0/fbr//sjMHKADnhTCWDRfCtddTYrUIUEYByOHJJnuSnOz82pqADLAbQOi4iECsM2NhAYBRQhj0+Po95AyiJlfKq9Ms3md2BGUKzf30NP2+gRb6QuwpDkg9AgyIHuC+qEpATpJ36f4JtiBR9Fh5l/KWqA1nAw3yfmBa9XimxCRGZSqe4vki0YEubmqJhO3f2SsKObZ2SqkTbefNlgSXL6mwMKSHgdjMowE0MrlGYLwQ+NIAo4NGsIqgmqlKjs7elgkYxRs64ihGrpiS6nOFqK/O1ie9LHQVxQUHBjp1fSW+pCRwiNUeiMFMsKIoMDX0jrPHjFWmkyfpZ3EfJC+pSgSZpqDpyjAQ+6mcBaCAqjWY0issSIyhOiv1tBohg8tg/3DETkqXFio+5S8PD9hgIqDkWeAUgW5lKj1ohqX0WNCv6WnzM3MTflmkhEKBYyl0QFbLW6tMCNBi8IDMalIK44JJXs9/VqfGEBcT+8DgeVpBKE9rL+eWEcuJCbCArpG6epYaLoxSqR5idIMjeCsn6RZ30p5WSx4iU0R7uU1A5QSpAAchfUnhEnKu7LbM3NLL7XbsJkwYjnWIKMwr7pbjIIqQKqQqgpozkLepS/K+byFJu4L9NbXZz1egO1W7S47UHDz4pEEOtQQTc+A2p4WsaHe+R9lDimz0aZJyWI5PVVJFYB6mW1/Ax9viTl4gCxMEyMqLaUHe+nsVPx8JsaFV//fSe9DgRpnklHVIV6PykVP4W+8fuVgrQRzGYXqZCV899/o/+3m6ku3vlrXuubGhWdNkM2MdS0tD5okdwqiUMpZun6vxJm+r0YE1FT03y4JI08IyGbkKKT5EjR+nfwrsZR6pNapszzht8Dmcu+gdwB99Ko9cbZ8WEcHW7HT/7qx7H7bDOGB0ChHMXo+MV4vP4sbnzwUdT6m3HCmPHaBInjNC1cUCII7R8clFzE0tKSm+a5f2j+YQIoPVT8KowMYv/lfMKEzIyQHqFk5ufn4u7SYhY/WyoYkXzJdB7k/MFBjE+C8qcZ4NciaSfhvPbaq7G4tGQTVJKxNNarvACpXAklmkWTNv2Dun0iCgrq6yIGS6WZMSXmQhaliu+RmCv5h5IMkQa3m6buaqVMGEheFUV6pa/q/kca/n0l0fqfYxc3+7xuNC+7Gm4uJrdBxZl0mtFT9sic5e39si4ZOxdkxNiq9arRbnO8Zjvh4dlKSkMNghPFHcwpSx+Z5dJBulrXd2vrWXs9kiAguVAS+9wtuhBvblQw3qWZUM5zGSQXecti6qeiISxBF64BAHBWEY+0C+S5rkui6kTFib6bNtz7keUJuvoF2guVpXeSYF1LFvBAspJ/9zco2hfN3x7FYBRkFq7OyqzextP1WLq/EkuwR1PCxOddYUZl0pnPsZthYgRcFr9Tk7iAJIhBtJZhoapxZQYpCZxYVtkbbTfV03zRkhFG6xVGRXuXTf8o+6O4aMF60nxmOqvwaT8V4hPOFIEAkHlKZqrYRGqMARJwc8R63WlinQxQox07H+W5OC5gngHEcHOMvy8SA74qNwbtG9PbMbHM5oXlBvJoL1KL+b3c5pP91PE8cnPH54LXJ8UnM06RJOJz5i5jxtlJY4Fr5gwuhajSRC6AjbZMYJ6bYvcSF6TmOnsC5zxrk3scGhnSz+23MahzuTQKVcCSmfuZCnDsQdMzU7Gz/SyGQOpyLccnMTYxEYdHJ0JHjw0Pxunhfpwe7Mb4UH9cm52KrY21GB4di6mpmVhaXo3FeyvRGByK5uBQXJqdjUdrT8R65R7Y+w+Pacwxx040JqC1YeQQkxGDUURnvQkwlAU5muiAgYhxKeoYYNOreKPso5qjySTiebEHPd/d1R7PfsJzZcwpPlj65SxaBwdx9epsrK2t694w0qYhQNFNDSfmNRrZR8ihGjyiomPKUhDLs96tOQ77GIPbghCF1WLJtHp/Q6wHZJ9gK9AEUHEDJlJKoOlZSnbO8RP5BOck18jUpqAjlPrBgeRm2KPIiWAJsE+RCwAEoghMoZv5hGcTcwIUJ2cH8S4G5GoI7dsU9Nq1hZgaH1dhnTsm3saoegzfkNOzuLt0P7YACeW5QsFca7JSlbk0PiCWhDLauuResAH66jUVbIssaAFIcf5ZUz/HSFJLyGjZg4Ez3LEu8lfO2fhcDTnYBZVKPNv2WcB6kR+M9oMeMfpPj1oxM3Uh+hsNSc7yLGkCbGxtyheBU9YxxLkaBgKc5HkFQ1QF354XYgcwbjSQS1NbsUsyk3n/K7OvSEbSYK0TFdevLlxp92oZK+WHZ2eaWyBrQeDTpGAfxIh6bx8T4zMxBsjDYauMDA7FALLHO89jZmZaBfTmoH2OWAfNRn+MTF6Mk+NzeW/QWNjf2Yn93R3FMrAA1zY3Y219U1LBFy5MxfzVKzEyNBT9jaYYG+TVvM5+6zBu3v6N9NvHxsdjZ3fXiHmBzlg3vTExMRbDg/26T+SiFuYXtHMaxMXaYI1VBCjgeRMbMraSelKR1N4fnC80CUfGRuLjTz6J+8v325JhNAvefuedmBibaJs6I3lIo4XYDJYra2zxi881LmiDwkC6NH0hpqcvqoFJHCFm7uRULK+uxs1bt+PBysNoDAyKjRgVAAuWG6TBxnvyTGmcrTy8rxiFJhAMNOIR2DLIpbEvXbo0E08erQrMxrigY0/TEENtCu3IwPAxhRLE+rrWJWc262N7d8fAMuSLmAsoFSQzW14g2QRjfAqLQfJZe3gJpQ9CxmfFB1Ey2xWkQ1t+rzxXlU8lgKnEUGpY5zriZ2W+83mRGFTsk/6RnP/cD+utsADK+i1Hrc9c78eckAXoovi2DcRz3mQGmOXH2ns2vgNd3onOVd3w9fXr/21gJd/muTH2qsmkN4Jfn6YF98g8NKOQz4vXxJcQDiVMSDaDw+fiS9qROvq6ULqTX5q14kZMd6Oik+eViMGgGQNoij8FZ4r8EBTDOb8pc8Cxi+NXPkojpPP8OBvs21HGvjtAKTm8Abf2z3D+VkzBHU9ZajZz0QSVGvDh3L3k6wJMZmPE1+N4jmvXuLfHz8Bc1cxKoyLvLbnEfrb5XtwnZ3GJ0ct9SiWF+mPOBDXVxNTzfqOGSDIqxodq8eb1y1GvnEbvi7MYbA5Eta8ZPdV6fPzp3Tg4Pos6sc8LGGn9ce/+sszo7QlmwBRfI7vn+6hEb62qM3Nrc9Pm7CldSv2PWh45P+c+dU1iARhTYsg16jHQDzDuOJ6ub8Zf/+WfxOryo1h9sKzGwvwcPjxjcfPmzajVfR8/ff/v4p//8V8U7yLp9MZ3X9Ne89uPPom+vkqMT03He9//AzlabR0exJ1PP4319adSJfhW+ulLIf+3X/x/GIHpcLBV2ALauKqVDBB9GMASAJkDlZADcGFuTl3Nu3fvKsAg0Gdxiwp12IqnGzZ34QMEFAG2KfbjOuSgTQ40B2JxaTGGRkaUPPAebJBsOPwN13Hl6hU1QljwsBUoRqEf7mKw2Qa8d0FLyfjrsBVv/d5b8eSxTbYJ+ihos3myscngJk1FeR2o93wQkNuszsGx8m/px3c2/XbxBgRYUuhJ6kBKkPQ9QP5qYDAGh4d0nTt7uwpoCOCEinvRo6bE9vNtmWk5OXRjgITGLXlr/nHgSIOZsc0gWY0jivgyC3OxuJgMUZjqblQURKTMovGR2EerNOUCspDCvYJIExJc0iNmUqhRkUbdILiErDs+VnBJE8KIX6N1Sa5FPYXiiawSXgqim3OIdfT3ua/SMBELRE0ZDmG/DoE49809EMjyfgTmKjwgq0HCIqP3uqjLHCAEv4whh4SeXUpwFCmoQpO32VinyeAignXSSVjRIaWJxGsQSJJYoF8spgDNgETYiCUhrwh0Tb1mFOhp/DqyGTIVTQ+Jgmbh70qg4LmVgUu7eN0BnLoQ2NG0V4ACbRXDTz27Ykrdkf7pZkCUwrVus6sZUvwoJDWTdHVLzhhpI738NNcSSqN4JySboB0AZRGu3fhJgzVJXlEUaRsOO8grzRseIIVh7kVMJ6SmhJQgifGcYh/RtUAxTf30b2gjtNkfpaHQQcE4+C6UZQVyyfZ5ec8u8+Lr9nI9sTbDxsuThJeGmBEsvlY3tJDoSUmZTNQKMlxI5XyDrzYqCjEgUetdjIp2o689X7LwLINfNw1Yw0brlmK3A0k3qnJPyXnQHWBLWipZOX4t8MJGnCsNyKaOCnrZmNCeUu1xEay3V8mKC8IuBl26PCOml2ShKM6gE3x6FHHWir//2U9iHckEzHcbQzEyNhkffvxZrG5sylR777AlKYPj1pHWP2PN3sIaHhpGIzykCQzqRz42uR8wtpZGAXFoJCnB/tW5qyrg4BXEc+D7GCB+8NF/es8hGG4OaK0XlDRz7sLFC0ruV1YfqgGvNR4Rs3NXY3llRck6jQqkLOS5QwIk8+9zYk43BkQ/71dxp8yvDjLpqzPNa7TQzS2NyHsWpJQTACOn5fujJkr6n7hf0JYmqiONh5wa3kfqbnve/u8YFQXhVq7Vsl+yMlCBleJC+Zn3MRlQp1RYScTEqkl5MiD+pUjMBYHsbTbrNhat9OiZSfIomW7Wa3eRh9cQiKKPZqHp+mIRVGmooq29nue0C88qZOUcFQMwM+iSfBVmRTnfu5M+Faa7EPUYrirpTISdDV/HY2PDpphmWlliqzwn7o39rMN0BH3tM7Rd2lbe7SKNrieLDRQ+283ZnohGDc16I8hLkRIjPoxlX7++IONAn+u98XR7J+58+rkKbmpuFX3gLAapmSxGpJubxXtHjUsllj4DnPR57y57WEmq3aB+oQaFEzrLB2g9FDk0xTCcJZ53AkhkXFEAIpyZmg/abCwHoYZh8UOR3i9NLMAdLt6wnxXD6LLnlzkljzIlzt7AStPW52zno3ztAkHeg7yy6lr3kh9JlDTN2hIIWp6tMHKyYC1dbsscyucj0aduWHl8PX/MrJQJMmsbg8m+mlnGan65sL54dzFGJ8ZUsCPGYv8g7lazHTZwSomJeVZkESkEp1dG8QCTFDTylvLJ2VfhntfQ12kQybWoSA9afn3dEowgqSX/Yx8MGFGWsewNcCgHe7sxNDCoOcx86x8eVjH/O69ei/3trdh++iRGBxrxysXxGB8aVENgcmomHjx8HJ99QZO5GZMz0zHzyqwY0uiyEzf3AAyRUCBFvUNJclKIbhdBpEVeMds7vVFAfAuYcmSDZu6XmFLPr2iVMzY57zhbnm6RyDMGBxrL8QmAUhtmPqefAtrwFCKYD5IgOzmKSzPTkvrDp0D7OYAFzW/iKLOXaHax7gFF8Tcu6Ha8/Th/aDpQwCFHEMsA1twp52U9nm5uSl5n/+BQZwmeGjQbWD/EHPy3ubmVcmBIKwLWOYiRoREVbGEWs+dTYKE4+XRzSzH17CuXNI8eP14TM8JSmztR663Gd157TYCy6QsXdC/I+Eim5+m65KAmJyZiYW7eBdKTM2nvc6CAsl/f3JRkFQV4Jpf97c5VYGJukVeV2BK5qBKnCARRsw8TMrBat6BSM89hEthfyWhanymW3JX0T7USW1vbLqRlZ5gxlVfA+ISAb3yfQpJQ1iqCnot9cH5yHBcnJsVKGEL6cX8/xibH49nuTmwjY5UoX/YtMX6zUeHmBbE366VP43Ry3JKPCfsa98Q5wD3Kn4xmS6UnXnv1VRWtHj1aleTk1QUMt7/nfKni2E0Mc0AZraOYnp5WTs28vnPnjuYpYwfYj+b7yPBgtGjcVSoxiuwaMQy+hNWI7775phouN351I55tt6KShTbF39WqDF0JgWn0HwPuOmSOVqLZgDV+KumnN15/PTXfa5LRpCEFe+bf/v0/1EDDZHx/vyVPSE5ETKf7++uSiQN48OTRI3nfwFRhzPABZJ3QEBHLgjPxhFyfhoeLejSiASAWhDWd+ef7u/FPv/iF5jBsH0lOnVfij3/wXswvzOv5Yqotj8aBARWEYZAufXFX48f+xz1h/k4M+r233wqM1okl5Hd2+VKsPliJX924GY/W1qNSrUUPTRX+rVRlPO+9uRITk5Px5PGq9kBQ1jTgmvWmgIliiYjpMSzPFZ45jRFYSsOjo6oLsKcTE/N8AU8iF6Wmw7kR17BGkC6lLiFmFzlSveYGPSAvZE1V5zCDQevh9EwNORes3TQyM9D+Wm4QOUZE8aIw9GgbCOiWjFE+5+/Ym0otoYDU+Jo4tBSYeb1SgDeKvE85HN830r+cu5zr5Ft5roshzLN2HOc4yb/LOlGzqi2xliC4lIkj76fe0A3ukA9AOzfpgLvKdRQmWonXAIkK+6E16UZUiS07Bf4O8MzBQ3rJdEmF+hozsm3jSjoAkxJzFK8P5UQvxR4lhiqxfpHiVGyv2pd9VUp5opxlYq9IktGNU35PwN4E4hqk5yaBSwf2aXSc3ol/PPbnLvbn8xRYg3pOelEItJismpL7eUjcvLDfYsdku9xiqR0YQFLiTOfHfu7kwB3AlWPWBFplDUSxH3kP4F8x3S0vzudFJtVxoOtBmtcpl1mArNSr6vWeODl4FvOXR2P24kScHx3G9YVrcfvWhzH/6uvx4SdfCDRxhmdYD15r9Vi6tyy2BPuU4tZk3vB6xZ+EsXrl0uXY2FgXm5M8l7OXuhDr2HHaueQLFaOlj6EBk9TGTuL51nr8+Ed/GvcXl2Nt9aHyqIWF6wJ4w6gA5MD7/e1P/yZ+/g8/l8wrOc47b78h/xnk7ohN8P9699239PUf/fAH0RhoSj7v1u3fxH8DABsndDLwolsAAAAASUVORK5CYII="/>
</defs>
</svg>
